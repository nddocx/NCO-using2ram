module counter (clk,
    csb00,
    csb01,
    rst,
    addr00,
    addr01,
    din00,
    din01,
    sine_out);
 input clk;
 input csb00;
 input csb01;
 input rst;
 input [7:0] addr00;
 input [7:0] addr01;
 input [15:0] din00;
 input [15:0] din01;
 output [15:0] sine_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire net115;
 wire clknet_0_clk;
 wire \sine_out_temp0[0] ;
 wire \sine_out_temp0[10] ;
 wire \sine_out_temp0[11] ;
 wire \sine_out_temp0[12] ;
 wire \sine_out_temp0[13] ;
 wire \sine_out_temp0[14] ;
 wire \sine_out_temp0[15] ;
 wire \sine_out_temp0[1] ;
 wire \sine_out_temp0[2] ;
 wire \sine_out_temp0[3] ;
 wire \sine_out_temp0[4] ;
 wire \sine_out_temp0[5] ;
 wire \sine_out_temp0[6] ;
 wire \sine_out_temp0[7] ;
 wire \sine_out_temp0[8] ;
 wire \sine_out_temp0[9] ;
 wire \sine_out_temp1[0] ;
 wire \sine_out_temp1[10] ;
 wire \sine_out_temp1[11] ;
 wire \sine_out_temp1[12] ;
 wire \sine_out_temp1[13] ;
 wire \sine_out_temp1[14] ;
 wire \sine_out_temp1[15] ;
 wire \sine_out_temp1[1] ;
 wire \sine_out_temp1[2] ;
 wire \sine_out_temp1[3] ;
 wire \sine_out_temp1[4] ;
 wire \sine_out_temp1[5] ;
 wire \sine_out_temp1[6] ;
 wire \sine_out_temp1[7] ;
 wire \sine_out_temp1[8] ;
 wire \sine_out_temp1[9] ;
 wire \tcout[0] ;
 wire \tcout[1] ;
 wire \tcout[2] ;
 wire \tcout[3] ;
 wire \tcout[4] ;
 wire \tcout[5] ;
 wire \tcout[6] ;
 wire \tcout[7] ;
 wire \tcout[8] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__inv_2 _061_ (.A(\tcout[0] ),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _062_ (.A(net112),
    .Y(_025_));
 sky130_fd_sc_hd__mux2_1 _063_ (.A0(\sine_out_temp0[0] ),
    .A1(\sine_out_temp1[0] ),
    .S(net84),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _064_ (.A0(\sine_out_temp0[1] ),
    .A1(net76),
    .S(net84),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _065_ (.A0(\sine_out_temp0[2] ),
    .A1(net75),
    .S(net84),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _066_ (.A0(\sine_out_temp0[3] ),
    .A1(net74),
    .S(net84),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _067_ (.A0(\sine_out_temp0[4] ),
    .A1(net73),
    .S(net84),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _068_ (.A0(\sine_out_temp0[5] ),
    .A1(net72),
    .S(net84),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _069_ (.A0(\sine_out_temp0[6] ),
    .A1(net71),
    .S(net83),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _070_ (.A0(\sine_out_temp0[7] ),
    .A1(net70),
    .S(net83),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _071_ (.A0(\sine_out_temp0[8] ),
    .A1(net69),
    .S(net83),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _072_ (.A0(\sine_out_temp0[9] ),
    .A1(net68),
    .S(net83),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _073_ (.A0(\sine_out_temp0[10] ),
    .A1(net82),
    .S(net83),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _074_ (.A0(\sine_out_temp0[11] ),
    .A1(net81),
    .S(net83),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _075_ (.A0(\sine_out_temp0[12] ),
    .A1(net80),
    .S(net83),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _076_ (.A0(\sine_out_temp0[13] ),
    .A1(net79),
    .S(net83),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _077_ (.A0(\sine_out_temp0[14] ),
    .A1(net78),
    .S(net83),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _078_ (.A0(\sine_out_temp0[15] ),
    .A1(net77),
    .S(net83),
    .X(_006_));
 sky130_fd_sc_hd__xor2_1 _079_ (.A(net107),
    .B(\tcout[1] ),
    .X(_017_));
 sky130_fd_sc_hd__and3_1 _080_ (.A(net109),
    .B(net105),
    .C(net102),
    .X(_050_));
 sky130_fd_sc_hd__a21oi_1 _081_ (.A1(net110),
    .A2(net105),
    .B1(net102),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_1 _082_ (.A(_050_),
    .B(_051_),
    .Y(_018_));
 sky130_fd_sc_hd__and4_2 _083_ (.A(net109),
    .B(net105),
    .C(\tcout[2] ),
    .D(\tcout[3] ),
    .X(_052_));
 sky130_fd_sc_hd__nor2_1 _084_ (.A(\tcout[3] ),
    .B(_050_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_1 _085_ (.A(_052_),
    .B(_053_),
    .Y(_019_));
 sky130_fd_sc_hd__xor2_1 _086_ (.A(\tcout[4] ),
    .B(_052_),
    .X(_020_));
 sky130_fd_sc_hd__and3_1 _087_ (.A(net96),
    .B(net93),
    .C(_052_),
    .X(_054_));
 sky130_fd_sc_hd__a21oi_1 _088_ (.A1(net96),
    .A2(_052_),
    .B1(net93),
    .Y(_055_));
 sky130_fd_sc_hd__nor2_1 _089_ (.A(_054_),
    .B(_055_),
    .Y(_021_));
 sky130_fd_sc_hd__xor2_1 _090_ (.A(\tcout[6] ),
    .B(_054_),
    .X(_022_));
 sky130_fd_sc_hd__and2_1 _091_ (.A(net88),
    .B(\tcout[7] ),
    .X(_056_));
 sky130_fd_sc_hd__and4_1 _092_ (.A(net95),
    .B(\tcout[5] ),
    .C(_052_),
    .D(_056_),
    .X(_057_));
 sky130_fd_sc_hd__a41o_1 _093_ (.A1(net95),
    .A2(net92),
    .A3(net88),
    .A4(_052_),
    .B1(\tcout[7] ),
    .X(_058_));
 sky130_fd_sc_hd__and2b_1 _094_ (.A_N(_057_),
    .B(_058_),
    .X(_023_));
 sky130_fd_sc_hd__xor2_1 _095_ (.A(net84),
    .B(_057_),
    .X(_024_));
 sky130_fd_sc_hd__inv_2 _096_ (.A(net111),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _097_ (.A(net111),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _098_ (.A(net111),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _099_ (.A(net111),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _100_ (.A(net112),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _101_ (.A(net112),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _102_ (.A(net112),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _103_ (.A(net112),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _104_ (.A(net112),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _105_ (.A(net111),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _106_ (.A(net111),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _107_ (.A(net111),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _108_ (.A(net111),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _109_ (.A(net111),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _110_ (.A(net111),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _111_ (.A(net113),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _112_ (.A(net113),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _113_ (.A(net113),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _114_ (.A(net113),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _115_ (.A(net113),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _116_ (.A(net113),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _117_ (.A(net113),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _118_ (.A(net112),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _119_ (.A(net112),
    .Y(_049_));
 sky130_fd_sc_hd__dfrtp_1 _120_ (.CLK(clknet_2_1__leaf_clk),
    .D(_014_),
    .RESET_B(_025_),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_1 _121_ (.CLK(clknet_2_0__leaf_clk),
    .D(_015_),
    .RESET_B(_026_),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _122_ (.CLK(clknet_2_1__leaf_clk),
    .D(_001_),
    .RESET_B(_027_),
    .Q(net53));
 sky130_fd_sc_hd__dfrtp_1 _123_ (.CLK(clknet_2_0__leaf_clk),
    .D(_002_),
    .RESET_B(_028_),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_1 _124_ (.CLK(clknet_2_0__leaf_clk),
    .D(_003_),
    .RESET_B(_029_),
    .Q(net55));
 sky130_fd_sc_hd__dfrtp_1 _125_ (.CLK(clknet_2_0__leaf_clk),
    .D(_004_),
    .RESET_B(_030_),
    .Q(net56));
 sky130_fd_sc_hd__dfrtp_1 _126_ (.CLK(clknet_2_0__leaf_clk),
    .D(_005_),
    .RESET_B(_031_),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _127_ (.CLK(clknet_2_1__leaf_clk),
    .D(_006_),
    .RESET_B(_032_),
    .Q(net58));
 sky130_fd_sc_hd__dfrtp_1 _128_ (.CLK(clknet_2_0__leaf_clk),
    .D(_016_),
    .RESET_B(_033_),
    .Q(\tcout[0] ));
 sky130_fd_sc_hd__dfrtp_1 _129_ (.CLK(clknet_2_0__leaf_clk),
    .D(_017_),
    .RESET_B(_034_),
    .Q(\tcout[1] ));
 sky130_fd_sc_hd__dfrtp_1 _130_ (.CLK(clknet_2_1__leaf_clk),
    .D(_018_),
    .RESET_B(_035_),
    .Q(\tcout[2] ));
 sky130_fd_sc_hd__dfrtp_1 _131_ (.CLK(clknet_2_1__leaf_clk),
    .D(_019_),
    .RESET_B(_036_),
    .Q(\tcout[3] ));
 sky130_fd_sc_hd__dfrtp_1 _132_ (.CLK(clknet_2_1__leaf_clk),
    .D(_020_),
    .RESET_B(_037_),
    .Q(\tcout[4] ));
 sky130_fd_sc_hd__dfrtp_1 _133_ (.CLK(clknet_2_1__leaf_clk),
    .D(_021_),
    .RESET_B(_038_),
    .Q(\tcout[5] ));
 sky130_fd_sc_hd__dfrtp_1 _134_ (.CLK(clknet_2_1__leaf_clk),
    .D(_022_),
    .RESET_B(_039_),
    .Q(\tcout[6] ));
 sky130_fd_sc_hd__dfrtp_1 _135_ (.CLK(clknet_2_3__leaf_clk),
    .D(_023_),
    .RESET_B(_040_),
    .Q(\tcout[7] ));
 sky130_fd_sc_hd__dfrtp_1 _136_ (.CLK(clknet_2_3__leaf_clk),
    .D(_024_),
    .RESET_B(_041_),
    .Q(\tcout[8] ));
 sky130_fd_sc_hd__dfrtp_1 _137_ (.CLK(clknet_2_2__leaf_clk),
    .D(_000_),
    .RESET_B(_042_),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_1 _138_ (.CLK(clknet_2_2__leaf_clk),
    .D(_007_),
    .RESET_B(_043_),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_1 _139_ (.CLK(clknet_2_2__leaf_clk),
    .D(_008_),
    .RESET_B(_044_),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _140_ (.CLK(clknet_2_3__leaf_clk),
    .D(_009_),
    .RESET_B(_045_),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_1 _141_ (.CLK(clknet_2_3__leaf_clk),
    .D(_010_),
    .RESET_B(_046_),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_1 _142_ (.CLK(clknet_2_3__leaf_clk),
    .D(_011_),
    .RESET_B(_047_),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_1 _143_ (.CLK(clknet_2_3__leaf_clk),
    .D(_012_),
    .RESET_B(_048_),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _144_ (.CLK(clknet_2_0__leaf_clk),
    .D(_013_),
    .RESET_B(_049_),
    .Q(net65));
 sky130_fd_sc_hd__conb_1 mem_i1_115 (.LO(net115));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 ram_256x16 mem_i0 (.csb0(net17),
    .csb1(net114),
    .clk0(clknet_2_2__leaf_clk),
    .clk1(clknet_2_1__leaf_clk),
    .addr0({net8,
    net7,
    net6,
    net5,
    net4,
    net3,
    net2,
    net1}),
    .addr1({net85,
    net87,
    net91,
    net94,
    net99,
    net101,
    net103,
    net108}),
    .din0({net25,
    net24,
    net23,
    net22,
    net21,
    net20,
    net34,
    net33,
    net32,
    net31,
    net30,
    net29,
    net28,
    net27,
    net26,
    net19}),
    .dout1({\sine_out_temp0[15] ,
    \sine_out_temp0[14] ,
    \sine_out_temp0[13] ,
    \sine_out_temp0[12] ,
    \sine_out_temp0[11] ,
    \sine_out_temp0[10] ,
    \sine_out_temp0[9] ,
    \sine_out_temp0[8] ,
    \sine_out_temp0[7] ,
    \sine_out_temp0[6] ,
    \sine_out_temp0[5] ,
    \sine_out_temp0[4] ,
    \sine_out_temp0[3] ,
    \sine_out_temp0[2] ,
    \sine_out_temp0[1] ,
    \sine_out_temp0[0] }));
 ram_256x16 mem_i1 (.csb0(net18),
    .csb1(net115),
    .clk0(clknet_2_2__leaf_clk),
    .clk1(clknet_2_0__leaf_clk),
    .addr0({net16,
    net15,
    net14,
    net13,
    net12,
    net11,
    net10,
    net9}),
    .addr1({net86,
    net89,
    net90,
    net97,
    net98,
    net100,
    net104,
    net106}),
    .din0({net41,
    net40,
    net39,
    net38,
    net37,
    net36,
    net50,
    net49,
    net48,
    net47,
    net46,
    net45,
    net44,
    net43,
    net42,
    net35}),
    .dout1({\sine_out_temp1[15] ,
    \sine_out_temp1[14] ,
    \sine_out_temp1[13] ,
    \sine_out_temp1[12] ,
    \sine_out_temp1[11] ,
    \sine_out_temp1[10] ,
    \sine_out_temp1[9] ,
    \sine_out_temp1[8] ,
    \sine_out_temp1[7] ,
    \sine_out_temp1[6] ,
    \sine_out_temp1[5] ,
    \sine_out_temp1[4] ,
    \sine_out_temp1[3] ,
    \sine_out_temp1[2] ,
    \sine_out_temp1[1] ,
    \sine_out_temp1[0] }));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_246_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_247_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_248_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_249_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_250_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_251_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_252_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_253_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_254_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_255_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_256_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_257_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_258_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_259_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_260_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_261_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_262_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_263_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_264_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_265_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_266_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_2_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_2_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_2_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_2_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_2_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_2_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_2_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_2_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_2_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_2_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_2_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_2_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_2_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_2_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_2_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_2_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_2_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_2_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_2_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_2_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_2_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_2_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_2_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_2_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_2_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_2_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_2_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_2_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_2_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_2_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_2_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_2_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_2_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_2_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_2_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_2_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_2_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_2_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_2_Right_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_2_Right_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_2_Right_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_2_Right_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_2_Right_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_2_Right_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_2_Right_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_2_Right_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_2_Right_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_2_Right_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_2_Right_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_2_Right_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_2_Right_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_2_Right_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_2_Right_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_2_Right_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_2_Right_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_2_Right_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_2_Right_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_2_Right_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_2_Right_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_2_Right_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_2_Right_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_2_Right_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_2_Right_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_2_Right_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_2_Right_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_2_Right_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_2_Right_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_2_Right_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_2_Right_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_2_Right_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_2_Right_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_2_Right_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_2_Right_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_2_Right_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_2_Right_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_2_Right_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_2_Right_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_2_Right_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_2_Right_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_2_Right_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_2_Right_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_2_Right_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_2_Right_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_2_Right_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_2_Right_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_2_Right_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_2_Right_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_2_Right_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_2_Right_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_2_Right_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_2_Right_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_2_Right_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_2_Right_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_2_Right_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_2_Right_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_2_Right_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_2_Right_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_2_Right_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_2_Right_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_2_Right_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_2_Right_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_2_Right_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_2_Right_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_2_Right_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_2_Right_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_2_Right_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_2_Right_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_1_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_1_Left_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_1_Left_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_1_Left_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_1_Left_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_1_Left_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_1_Left_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_1_Left_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_1_Left_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_1_Left_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_1_Left_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_1_Left_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_1_Left_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_1_Left_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_1_Left_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_1_Left_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_1_Left_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_1_Left_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_1_Left_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_1_Left_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_1_Left_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_1_Left_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_1_Left_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_1_Left_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_1_Left_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_1_Left_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_1_Left_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_1_Left_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_1_Left_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_1_Left_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_1_Left_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_1_Left_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_1_Left_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_1_Left_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_1_Left_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_1_Left_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_1_Left_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_1_Left_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_1_Left_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_1_Left_444 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_1_Left_445 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_1_Left_446 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_1_Left_447 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_1_Left_448 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_1_Left_449 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_1_Left_450 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_1_Left_451 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_1_Left_452 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_1_Left_453 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_1_Left_454 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_1_Left_455 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_1_Left_456 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_1_Left_457 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_1_Left_458 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_1_Left_459 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_1_Left_460 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_1_Left_461 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_1_Left_462 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_1_Left_463 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_1_Left_464 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_1_Left_465 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_1_Left_466 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_1_Left_467 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_1_Left_468 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_1_Left_469 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_1_Left_470 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_1_Left_471 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_1_Left_472 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_1_Left_473 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_1_Left_474 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_1_Left_475 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_1_Left_476 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_1_Left_477 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_1_Left_478 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_1_Left_479 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_1_Left_480 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_1_Left_481 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_1_Left_482 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_1_Left_483 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_1_Left_484 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_1_Left_485 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_1_Left_486 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_1_Left_487 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_1_Left_488 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_1_Left_489 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_1_Left_490 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_1_Left_491 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_1_Left_492 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_1_Left_493 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_1_Left_494 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_1_Left_495 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_1_Left_496 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_1_Left_497 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_1_Left_498 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_1_Left_499 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_1_Left_500 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_1_Left_501 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_1_Left_502 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_1_Left_503 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_1_Left_504 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_1_Left_505 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_1_Left_506 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_1_Left_507 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_1_Left_508 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_1_Left_509 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_1_Left_510 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_1_Left_511 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_246_Left_512 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_247_Left_513 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_248_Left_514 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_249_Left_515 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_250_Left_516 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_251_Left_517 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_252_Left_518 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_253_Left_519 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_254_Left_520 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_255_Left_521 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_256_Left_522 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_257_Left_523 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_258_Left_524 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_259_Left_525 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_260_Left_526 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_261_Left_527 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_262_Left_528 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_263_Left_529 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_264_Left_530 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_265_Left_531 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_266_Left_532 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Left_533 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_534 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_535 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_536 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_537 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_538 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_539 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_540 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_541 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_542 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_543 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_544 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_545 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_546 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_547 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_548 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_549 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_550 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_551 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_552 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_553 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_554 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_555 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_556 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_557 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_558 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_559 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_560 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_561 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_562 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_563 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_564 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_565 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_566 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_567 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_568 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_569 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_570 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_571 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_572 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_573 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_574 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_575 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_576 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_577 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_578 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_579 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_580 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_581 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_582 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_583 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_584 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_585 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_586 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_587 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_588 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_589 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_590 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Left_591 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Left_592 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Left_593 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Left_594 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Left_595 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Left_596 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Left_597 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Left_598 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Left_599 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Left_600 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Left_601 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Left_602 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Left_603 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Left_604 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Left_605 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Left_606 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Left_607 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Left_608 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Left_609 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Left_610 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Left_611 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Left_612 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Left_613 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Left_614 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Left_615 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Left_616 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Left_617 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Left_618 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Left_619 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Left_620 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Left_621 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Left_622 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Left_623 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Left_624 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Left_625 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Left_626 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Left_627 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Left_628 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Left_629 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Left_630 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Left_631 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Left_632 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Left_633 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Left_634 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Left_635 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Left_636 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Left_637 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Left_638 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Left_639 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Left_640 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Right_641 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Right_642 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Right_643 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Right_644 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Right_645 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Right_646 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Right_647 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Right_648 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Right_649 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Right_650 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Right_651 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Right_652 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Right_653 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Right_654 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Right_655 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Right_656 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Right_657 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Right_658 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Right_659 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Right_660 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Right_661 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Right_662 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Right_663 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Right_664 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Right_665 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Right_666 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Right_667 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Right_668 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Right_669 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Right_670 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Right_671 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Right_672 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Right_673 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Right_674 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Right_675 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Right_676 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Right_677 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Right_678 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Right_679 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Right_680 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Right_681 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Right_682 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Right_683 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Right_684 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Right_685 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Right_686 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Right_687 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Right_688 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Right_689 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Right_690 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Right_691 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Right_692 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Right_693 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Right_694 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Right_695 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Right_696 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Right_697 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Right_698 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Right_699 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Right_700 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Right_701 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Right_702 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Right_703 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Right_704 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Right_705 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Right_706 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Right_707 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Right_708 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Right_709 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Right_710 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Right_711 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Right_712 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Right_713 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Right_714 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Right_715 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Right_716 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Right_717 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Right_718 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Right_719 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Right_720 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Right_721 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Right_722 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Right_723 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Right_724 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Right_725 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Right_726 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Right_727 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Right_728 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Right_729 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Right_730 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Right_731 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Right_732 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Right_733 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Right_734 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Right_735 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Right_736 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Right_737 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Right_738 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Right_739 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Right_740 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Right_741 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Right_742 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Right_743 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Right_744 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Right_745 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Right_746 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Right_747 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_2_Left_748 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_2_Left_749 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_2_Left_750 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_2_Left_751 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_2_Left_752 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_2_Left_753 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_2_Left_754 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_2_Left_755 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_2_Left_756 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_2_Left_757 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_2_Left_758 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_2_Left_759 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_2_Left_760 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_2_Left_761 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_2_Left_762 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_2_Left_763 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_2_Left_764 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_2_Left_765 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_2_Left_766 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_2_Left_767 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_2_Left_768 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_2_Left_769 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_2_Left_770 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_2_Left_771 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_2_Left_772 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_2_Left_773 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_2_Left_774 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_2_Left_775 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_2_Left_776 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_2_Left_777 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_2_Left_778 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_2_Left_779 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_2_Left_780 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_2_Left_781 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_2_Left_782 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_2_Left_783 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_2_Left_784 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_2_Left_785 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_2_Left_786 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_2_Left_787 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_2_Left_788 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_2_Left_789 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_2_Left_790 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_2_Left_791 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_2_Left_792 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_2_Left_793 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_2_Left_794 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_2_Left_795 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_2_Left_796 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_2_Left_797 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_2_Left_798 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_2_Left_799 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_2_Left_800 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_2_Left_801 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_2_Left_802 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_2_Left_803 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_2_Left_804 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_2_Left_805 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_2_Left_806 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_2_Left_807 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_2_Left_808 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_2_Left_809 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_2_Left_810 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_2_Left_811 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_2_Left_812 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_2_Left_813 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_2_Left_814 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_2_Left_815 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_2_Left_816 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_2_Left_817 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_2_Left_818 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_2_Left_819 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_2_Left_820 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_2_Left_821 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_2_Left_822 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_2_Left_823 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_2_Left_824 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_2_Left_825 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_2_Left_826 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_2_Left_827 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_2_Left_828 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_2_Left_829 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_2_Left_830 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_2_Left_831 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_2_Left_832 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_2_Left_833 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_2_Left_834 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_2_Left_835 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_2_Left_836 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_2_Left_837 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_2_Left_838 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_2_Left_839 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_2_Left_840 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_2_Left_841 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_2_Left_842 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_2_Left_843 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_2_Left_844 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_2_Left_845 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_2_Left_846 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_2_Left_847 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_2_Left_848 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_2_Left_849 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_2_Left_850 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_2_Left_851 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_2_Left_852 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_2_Left_853 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_2_Left_854 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_1_Right_855 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_1_Right_856 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_1_Right_857 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_1_Right_858 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_1_Right_859 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_1_Right_860 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_1_Right_861 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_1_Right_862 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_1_Right_863 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_1_Right_864 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_1_Right_865 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_1_Right_866 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_1_Right_867 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_1_Right_868 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_1_Right_869 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_1_Right_870 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_1_Right_871 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_1_Right_872 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_1_Right_873 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_1_Right_874 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_1_Right_875 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_1_Right_876 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_1_Right_877 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_1_Right_878 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_1_Right_879 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_1_Right_880 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_1_Right_881 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_1_Right_882 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_1_Right_883 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_1_Right_884 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_1_Right_885 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_1_Right_886 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_1_Right_887 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_1_Right_888 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_1_Right_889 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_1_Right_890 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_1_Right_891 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_1_Right_892 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_1_Right_893 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_1_Right_894 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_1_Right_895 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_1_Right_896 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_1_Right_897 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_1_Right_898 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_1_Right_899 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_1_Right_900 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_1_Right_901 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_1_Right_902 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_1_Right_903 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_1_Right_904 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_1_Right_905 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_1_Right_906 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_1_Right_907 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_1_Right_908 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_1_Right_909 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_1_Right_910 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_1_Right_911 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_1_Right_912 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_1_Right_913 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_1_Right_914 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_1_Right_915 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_1_Right_916 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_1_Right_917 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_1_Right_918 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_1_Right_919 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_1_Right_920 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_1_Right_921 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_1_Right_922 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_1_Right_923 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_1_Right_924 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_1_Right_925 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_1_Right_926 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_1_Right_927 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_1_Right_928 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_1_Right_929 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_1_Right_930 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_1_Right_931 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_1_Right_932 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_1_Right_933 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_1_Right_934 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_1_Right_935 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_1_Right_936 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_1_Right_937 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_1_Right_938 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_1_Right_939 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_1_Right_940 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_1_Right_941 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_1_Right_942 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_1_Right_943 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_1_Right_944 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_1_Right_945 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_1_Right_946 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_1_Right_947 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_1_Right_948 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_1_Right_949 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_1_Right_950 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_1_Right_951 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_1_Right_952 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_1_Right_953 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_1_Right_954 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_1_Right_955 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_1_Right_956 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_1_Right_957 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_1_Right_958 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_1_Right_959 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_1_Right_960 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_1_Right_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_1_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_1_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_1_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_1_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_1_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_1_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_1_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_1_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_1_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_1_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_1_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_1_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_1_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_1_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_1_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_1_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_1_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_1_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_1_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_1_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_1_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_1_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_1_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_2_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_2_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_2_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_2_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_2_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_2_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_2_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_2_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_2_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_2_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_2_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_2_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_2_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_2_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_2_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_2_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_2_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_2_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_2_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_2_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_2_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_2_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_2_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_2_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_2_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_2_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_2_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_2_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_2_2491 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(addr00[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(addr00[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(addr00[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(addr00[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(addr00[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(addr00[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(addr00[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(addr00[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(addr01[0]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(addr01[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(addr01[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(addr01[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(addr01[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(addr01[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(addr01[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(addr01[7]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(csb00),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(csb01),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(din00[0]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(din00[10]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(din00[11]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(din00[12]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(din00[13]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(din00[14]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(din00[15]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(din00[1]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(din00[2]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(din00[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(din00[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(din00[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(din00[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(din00[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(din00[8]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(din00[9]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(din01[0]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(din01[10]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(din01[11]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(din01[12]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(din01[13]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(din01[14]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(din01[15]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(din01[1]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(din01[2]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(din01[3]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(din01[4]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(din01[5]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(din01[6]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(din01[7]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(din01[8]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(din01[9]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(rst),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net52),
    .X(sine_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .X(sine_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net54),
    .X(sine_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(sine_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(sine_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(sine_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(sine_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(sine_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(sine_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(sine_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(sine_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net63),
    .X(sine_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net64),
    .X(sine_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net65),
    .X(sine_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(sine_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(sine_out[9]));
 sky130_fd_sc_hd__clkbuf_2 wire68 (.A(\sine_out_temp1[9] ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 wire69 (.A(\sine_out_temp1[8] ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 wire70 (.A(\sine_out_temp1[7] ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 wire71 (.A(\sine_out_temp1[6] ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 wire72 (.A(\sine_out_temp1[5] ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 wire73 (.A(\sine_out_temp1[4] ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 wire74 (.A(\sine_out_temp1[3] ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 wire75 (.A(\sine_out_temp1[2] ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 wire76 (.A(\sine_out_temp1[1] ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 wire77 (.A(\sine_out_temp1[15] ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 wire78 (.A(\sine_out_temp1[14] ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 wire79 (.A(\sine_out_temp1[13] ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 wire80 (.A(\sine_out_temp1[12] ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 wire81 (.A(\sine_out_temp1[11] ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 wire82 (.A(\sine_out_temp1[10] ),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__buf_4 fanout84 (.A(\tcout[8] ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 load_slew85 (.A(\tcout[7] ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 load_slew86 (.A(\tcout[7] ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 load_slew87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 load_slew88 (.A(\tcout[6] ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 load_slew89 (.A(\tcout[6] ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 load_slew90 (.A(net93),
    .X(net90));
 sky130_fd_sc_hd__buf_2 load_slew91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 load_slew92 (.A(\tcout[5] ),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 load_slew93 (.A(\tcout[5] ),
    .X(net93));
 sky130_fd_sc_hd__buf_2 load_slew94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 load_slew95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 load_slew96 (.A(\tcout[4] ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 load_slew97 (.A(\tcout[4] ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 load_slew98 (.A(\tcout[3] ),
    .X(net98));
 sky130_fd_sc_hd__buf_2 load_slew99 (.A(\tcout[3] ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 load_slew100 (.A(net102),
    .X(net100));
 sky130_fd_sc_hd__buf_2 load_slew101 (.A(\tcout[2] ),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 load_slew102 (.A(\tcout[2] ),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 load_slew103 (.A(net105),
    .X(net103));
 sky130_fd_sc_hd__buf_2 load_slew104 (.A(\tcout[1] ),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 load_slew105 (.A(\tcout[1] ),
    .X(net105));
 sky130_fd_sc_hd__buf_2 load_slew106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 load_slew107 (.A(\tcout[0] ),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 load_slew108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 load_slew109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 load_slew110 (.A(\tcout[0] ),
    .X(net110));
 sky130_fd_sc_hd__buf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_4 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net51),
    .X(net113));
 sky130_fd_sc_hd__conb_1 mem_i0_114 (.LO(net114));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload0 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload1 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__D (.DIODE(_001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__X (.DIODE(_001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__D (.DIODE(_012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__X (.DIODE(_012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__D (.DIODE(_013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__X (.DIODE(_013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__D (.DIODE(_014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__X (.DIODE(_014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__D (.DIODE(_015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__072__X (.DIODE(_015_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(addr00[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(addr00[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(addr00[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(addr00[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(addr00[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(addr00[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(addr00[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(addr00[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(addr01[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(addr01[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(addr01[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(addr01[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(addr01[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(addr01[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(addr01[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(addr01[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(csb00));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(csb01));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(din00[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(din00[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(din00[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(din00[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(din00[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(din00[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(din00[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(din00[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(din00[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(din00[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(din00[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(din00[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(din00[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(din00[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(din00[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(din00[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(din01[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(din01[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(din01[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(din01[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(din01[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(din01[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(din01[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(din01[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(din01[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(din01[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(din01[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(din01[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(din01[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(din01[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(din01[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(din01[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[0]  (.DIODE(\sine_out_temp0[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__063__A0 (.DIODE(\sine_out_temp0[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[10]  (.DIODE(\sine_out_temp0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__A0 (.DIODE(\sine_out_temp0[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[11]  (.DIODE(\sine_out_temp0[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__074__A0 (.DIODE(\sine_out_temp0[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[12]  (.DIODE(\sine_out_temp0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__A0 (.DIODE(\sine_out_temp0[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[13]  (.DIODE(\sine_out_temp0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__076__A0 (.DIODE(\sine_out_temp0[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[14]  (.DIODE(\sine_out_temp0[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__077__A0 (.DIODE(\sine_out_temp0[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[15]  (.DIODE(\sine_out_temp0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__078__A0 (.DIODE(\sine_out_temp0[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[1]  (.DIODE(\sine_out_temp0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__064__A0 (.DIODE(\sine_out_temp0[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[2]  (.DIODE(\sine_out_temp0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__065__A0 (.DIODE(\sine_out_temp0[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[3]  (.DIODE(\sine_out_temp0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__066__A0 (.DIODE(\sine_out_temp0[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[4]  (.DIODE(\sine_out_temp0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__A0 (.DIODE(\sine_out_temp0[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[5]  (.DIODE(\sine_out_temp0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__A0 (.DIODE(\sine_out_temp0[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[6]  (.DIODE(\sine_out_temp0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__A0 (.DIODE(\sine_out_temp0[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[7]  (.DIODE(\sine_out_temp0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__A0 (.DIODE(\sine_out_temp0[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[8]  (.DIODE(\sine_out_temp0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__A0 (.DIODE(\sine_out_temp0[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[9]  (.DIODE(\sine_out_temp0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__072__A0 (.DIODE(\sine_out_temp0[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[0]  (.DIODE(\sine_out_temp1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__063__A1 (.DIODE(\sine_out_temp1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[0]  (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[1]  (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[2]  (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[3]  (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[4]  (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[5]  (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[6]  (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[7]  (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr0[0]  (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr0[1]  (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i0_csb0 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[0]  (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[1]  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[2]  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[3]  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[4]  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[0]  (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[10]  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[11]  (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[12]  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[13]  (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[14]  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[15]  (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[1]  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[2]  (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[3]  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[4]  (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[5]  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[6]  (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[7]  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[8]  (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[9]  (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__Q (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__Q (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__Q (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__Q (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__Q (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output59_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__Q (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__Q (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_output61_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__Q (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__Q (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__Q (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__Q (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__Q (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__Q (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__Q (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire68_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__072__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire69_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire70_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire71_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire72_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire73_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire74_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__066__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire75_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__065__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire76_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__064__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire77_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__078__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire78_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__077__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire79_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__076__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire80_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire81_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__074__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire82_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_X (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__078__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__077__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__076__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__074__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__072__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__095__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__066__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__065__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__064__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__063__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew85_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[7]  (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew87_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[6]  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew91_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[5]  (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew94_X (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[4]  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew97_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[4]  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew98_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[3]  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew99_X (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[3]  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew100_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[2]  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew101_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[2]  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew104_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[1]  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew106_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[0]  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__100__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__101__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__102__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__119__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__118__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__104__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__103__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__062__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__111__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__117__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__116__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__115__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__114__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__113__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__112__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__128__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__129__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i1_clk1 (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__131__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__132__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__133__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__134__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i0_clk1 (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload0_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i0_clk0 (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i1_clk0 (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload1_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_009_));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1148 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1167 ();
endmodule
