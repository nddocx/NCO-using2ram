VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter
  CLASS BLOCK ;
  FOREIGN counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 650.000 ;
  PIN addr00[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END addr00[0]
  PIN addr00[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END addr00[1]
  PIN addr00[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END addr00[2]
  PIN addr00[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END addr00[3]
  PIN addr00[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END addr00[4]
  PIN addr00[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END addr00[5]
  PIN addr00[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END addr00[6]
  PIN addr00[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END addr00[7]
  PIN addr01[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END addr01[0]
  PIN addr01[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END addr01[1]
  PIN addr01[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END addr01[2]
  PIN addr01[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END addr01[3]
  PIN addr01[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END addr01[4]
  PIN addr01[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END addr01[5]
  PIN addr01[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END addr01[6]
  PIN addr01[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END addr01[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 492.750 646.000 493.030 650.000 ;
    END
  END clk
  PIN csb00
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END csb00
  PIN csb01
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END csb01
  PIN din00[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END din00[0]
  PIN din00[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END din00[10]
  PIN din00[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END din00[11]
  PIN din00[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END din00[12]
  PIN din00[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END din00[13]
  PIN din00[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END din00[14]
  PIN din00[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END din00[15]
  PIN din00[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END din00[1]
  PIN din00[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END din00[2]
  PIN din00[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END din00[3]
  PIN din00[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END din00[4]
  PIN din00[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END din00[5]
  PIN din00[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END din00[6]
  PIN din00[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END din00[7]
  PIN din00[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END din00[8]
  PIN din00[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END din00[9]
  PIN din01[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END din01[0]
  PIN din01[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END din01[10]
  PIN din01[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END din01[11]
  PIN din01[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END din01[12]
  PIN din01[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END din01[13]
  PIN din01[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END din01[14]
  PIN din01[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END din01[15]
  PIN din01[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END din01[1]
  PIN din01[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END din01[2]
  PIN din01[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END din01[3]
  PIN din01[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END din01[4]
  PIN din01[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END din01[5]
  PIN din01[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END din01[6]
  PIN din01[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END din01[7]
  PIN din01[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END din01[8]
  PIN din01[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END din01[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 255.040 550.000 255.640 ;
    END
  END rst
  PIN sine_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END sine_out[0]
  PIN sine_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 319.640 550.000 320.240 ;
    END
  END sine_out[10]
  PIN sine_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 346.840 550.000 347.440 ;
    END
  END sine_out[11]
  PIN sine_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 329.840 550.000 330.440 ;
    END
  END sine_out[12]
  PIN sine_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 326.440 550.000 327.040 ;
    END
  END sine_out[13]
  PIN sine_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 340.040 550.000 340.640 ;
    END
  END sine_out[14]
  PIN sine_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 336.640 550.000 337.240 ;
    END
  END sine_out[15]
  PIN sine_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END sine_out[1]
  PIN sine_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END sine_out[2]
  PIN sine_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END sine_out[3]
  PIN sine_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END sine_out[4]
  PIN sine_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END sine_out[5]
  PIN sine_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END sine_out[6]
  PIN sine_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 323.040 550.000 323.640 ;
    END
  END sine_out[7]
  PIN sine_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 333.240 550.000 333.840 ;
    END
  END sine_out[8]
  PIN sine_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 343.440 550.000 344.040 ;
    END
  END sine_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 39.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 328.250 176.240 339.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 628.250 176.240 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 328.880 329.840 340.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 629.170 329.840 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 328.250 483.440 340.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 628.250 483.440 636.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 544.420 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 544.420 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 544.420 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 544.420 487.870 ;
    END
    PORT
      LAYER met4 ;
        RECT 529.580 35.120 531.180 332.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 529.580 337.040 531.180 634.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 21.040 629.900 544.420 631.500 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 328.250 179.540 340.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 628.250 179.540 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 328.250 333.140 340.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 628.250 333.140 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 328.250 486.740 340.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 628.250 486.740 636.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 544.420 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 544.420 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 544.420 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 544.420 491.170 ;
    END
    PORT
      LAYER met4 ;
        RECT 533.260 35.120 534.860 332.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 533.260 337.040 534.860 634.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 21.040 633.300 544.420 634.900 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 544.370 636.565 ;
      LAYER li1 ;
        RECT 5.520 10.795 544.180 636.565 ;
      LAYER met1 ;
        RECT 4.210 10.640 544.180 641.880 ;
      LAYER met2 ;
        RECT 4.230 645.720 492.470 646.000 ;
        RECT 493.310 645.720 542.710 646.000 ;
        RECT 4.230 4.280 542.710 645.720 ;
        RECT 4.230 4.000 115.730 4.280 ;
        RECT 116.570 4.000 122.170 4.280 ;
        RECT 123.010 4.000 128.610 4.280 ;
        RECT 129.450 4.000 135.050 4.280 ;
        RECT 135.890 4.000 141.490 4.280 ;
        RECT 142.330 4.000 144.710 4.280 ;
        RECT 145.550 4.000 151.150 4.280 ;
        RECT 151.990 4.000 157.590 4.280 ;
        RECT 158.430 4.000 164.030 4.280 ;
        RECT 164.870 4.000 170.470 4.280 ;
        RECT 171.310 4.000 176.910 4.280 ;
        RECT 177.750 4.000 180.130 4.280 ;
        RECT 180.970 4.000 186.570 4.280 ;
        RECT 187.410 4.000 193.010 4.280 ;
        RECT 193.850 4.000 199.450 4.280 ;
        RECT 200.290 4.000 205.890 4.280 ;
        RECT 206.730 4.000 209.110 4.280 ;
        RECT 209.950 4.000 215.550 4.280 ;
        RECT 216.390 4.000 542.710 4.280 ;
      LAYER met3 ;
        RECT 3.990 507.640 546.000 636.645 ;
        RECT 4.400 506.240 546.000 507.640 ;
        RECT 3.990 497.440 546.000 506.240 ;
        RECT 4.400 496.040 546.000 497.440 ;
        RECT 3.990 494.040 546.000 496.040 ;
        RECT 4.400 492.640 546.000 494.040 ;
        RECT 3.990 483.840 546.000 492.640 ;
        RECT 4.400 482.440 546.000 483.840 ;
        RECT 3.990 480.440 546.000 482.440 ;
        RECT 4.400 479.040 546.000 480.440 ;
        RECT 3.990 470.240 546.000 479.040 ;
        RECT 4.400 468.840 546.000 470.240 ;
        RECT 3.990 392.040 546.000 468.840 ;
        RECT 4.400 390.640 546.000 392.040 ;
        RECT 3.990 388.640 546.000 390.640 ;
        RECT 4.400 387.240 546.000 388.640 ;
        RECT 3.990 385.240 546.000 387.240 ;
        RECT 4.400 383.840 546.000 385.240 ;
        RECT 3.990 381.840 546.000 383.840 ;
        RECT 4.400 380.440 546.000 381.840 ;
        RECT 3.990 378.440 546.000 380.440 ;
        RECT 4.400 377.040 546.000 378.440 ;
        RECT 3.990 375.040 546.000 377.040 ;
        RECT 4.400 373.640 546.000 375.040 ;
        RECT 3.990 371.640 546.000 373.640 ;
        RECT 4.400 370.240 546.000 371.640 ;
        RECT 3.990 368.240 546.000 370.240 ;
        RECT 4.400 366.840 546.000 368.240 ;
        RECT 3.990 364.840 546.000 366.840 ;
        RECT 4.400 363.440 546.000 364.840 ;
        RECT 3.990 361.440 546.000 363.440 ;
        RECT 4.400 360.040 546.000 361.440 ;
        RECT 3.990 358.040 546.000 360.040 ;
        RECT 4.400 356.640 546.000 358.040 ;
        RECT 3.990 354.640 546.000 356.640 ;
        RECT 4.400 353.240 546.000 354.640 ;
        RECT 3.990 351.240 546.000 353.240 ;
        RECT 4.400 349.840 546.000 351.240 ;
        RECT 3.990 347.840 546.000 349.840 ;
        RECT 4.400 346.440 545.600 347.840 ;
        RECT 3.990 344.440 546.000 346.440 ;
        RECT 4.400 343.040 545.600 344.440 ;
        RECT 3.990 341.040 546.000 343.040 ;
        RECT 4.400 339.640 545.600 341.040 ;
        RECT 3.990 337.640 546.000 339.640 ;
        RECT 4.400 336.240 545.600 337.640 ;
        RECT 3.990 334.240 546.000 336.240 ;
        RECT 4.400 332.840 545.600 334.240 ;
        RECT 3.990 330.840 546.000 332.840 ;
        RECT 4.400 329.440 545.600 330.840 ;
        RECT 3.990 327.440 546.000 329.440 ;
        RECT 4.400 326.040 545.600 327.440 ;
        RECT 3.990 324.040 546.000 326.040 ;
        RECT 4.400 322.640 545.600 324.040 ;
        RECT 3.990 320.640 546.000 322.640 ;
        RECT 4.400 319.240 545.600 320.640 ;
        RECT 3.990 317.240 546.000 319.240 ;
        RECT 4.400 315.840 546.000 317.240 ;
        RECT 3.990 313.840 546.000 315.840 ;
        RECT 4.400 312.440 546.000 313.840 ;
        RECT 3.990 310.440 546.000 312.440 ;
        RECT 4.400 309.040 546.000 310.440 ;
        RECT 3.990 307.040 546.000 309.040 ;
        RECT 4.400 305.640 546.000 307.040 ;
        RECT 3.990 256.040 546.000 305.640 ;
        RECT 3.990 254.640 545.600 256.040 ;
        RECT 3.990 208.440 546.000 254.640 ;
        RECT 4.400 207.040 546.000 208.440 ;
        RECT 3.990 198.240 546.000 207.040 ;
        RECT 4.400 196.840 546.000 198.240 ;
        RECT 3.990 191.440 546.000 196.840 ;
        RECT 4.400 190.040 546.000 191.440 ;
        RECT 3.990 184.640 546.000 190.040 ;
        RECT 4.400 183.240 546.000 184.640 ;
        RECT 3.990 177.840 546.000 183.240 ;
        RECT 4.400 176.440 546.000 177.840 ;
        RECT 3.990 171.040 546.000 176.440 ;
        RECT 4.400 169.640 546.000 171.040 ;
        RECT 3.990 79.240 546.000 169.640 ;
        RECT 4.400 77.840 546.000 79.240 ;
        RECT 3.990 10.715 546.000 77.840 ;
      LAYER met4 ;
        RECT 50.000 627.850 174.240 632.225 ;
        RECT 176.640 627.850 177.540 632.225 ;
        RECT 179.940 628.770 327.840 632.225 ;
        RECT 330.240 628.770 331.140 632.225 ;
        RECT 179.940 627.850 331.140 628.770 ;
        RECT 333.540 627.850 481.440 632.225 ;
        RECT 483.840 627.850 484.740 632.225 ;
        RECT 487.140 627.850 509.900 632.225 ;
        RECT 50.000 340.720 509.900 627.850 ;
        RECT 50.000 339.800 177.540 340.720 ;
        RECT 50.000 327.850 174.240 339.800 ;
        RECT 176.640 327.850 177.540 339.800 ;
        RECT 179.940 328.480 327.840 340.720 ;
        RECT 330.240 328.480 331.140 340.720 ;
        RECT 179.940 327.850 331.140 328.480 ;
        RECT 333.540 327.850 481.440 340.720 ;
        RECT 483.840 327.850 484.740 340.720 ;
        RECT 487.140 327.850 509.900 340.720 ;
        RECT 50.000 40.720 509.900 327.850 ;
        RECT 50.000 39.800 177.540 40.720 ;
        RECT 50.000 22.615 174.240 39.800 ;
        RECT 176.640 22.615 177.540 39.800 ;
        RECT 179.940 22.615 327.840 40.720 ;
        RECT 330.240 22.615 331.140 40.720 ;
        RECT 333.540 22.615 481.440 40.720 ;
        RECT 483.840 22.615 484.740 40.720 ;
        RECT 487.140 22.615 509.900 40.720 ;
  END
END counter
END LIBRARY

