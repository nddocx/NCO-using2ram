VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter
  CLASS BLOCK ;
  FOREIGN counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 750.000 ;
  PIN addr00[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END addr00[0]
  PIN addr00[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END addr00[1]
  PIN addr00[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END addr00[2]
  PIN addr00[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END addr00[3]
  PIN addr00[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END addr00[4]
  PIN addr00[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END addr00[5]
  PIN addr00[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END addr00[6]
  PIN addr00[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END addr00[7]
  PIN addr01[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END addr01[0]
  PIN addr01[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END addr01[1]
  PIN addr01[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END addr01[2]
  PIN addr01[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END addr01[3]
  PIN addr01[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END addr01[4]
  PIN addr01[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END addr01[5]
  PIN addr01[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END addr01[6]
  PIN addr01[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END addr01[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END clk
  PIN csb00
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END csb00
  PIN csb01
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END csb01
  PIN din00[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END din00[0]
  PIN din00[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END din00[10]
  PIN din00[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END din00[11]
  PIN din00[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END din00[12]
  PIN din00[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END din00[13]
  PIN din00[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END din00[14]
  PIN din00[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END din00[15]
  PIN din00[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END din00[1]
  PIN din00[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END din00[2]
  PIN din00[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END din00[3]
  PIN din00[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END din00[4]
  PIN din00[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END din00[5]
  PIN din00[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END din00[6]
  PIN din00[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END din00[7]
  PIN din00[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END din00[8]
  PIN din00[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END din00[9]
  PIN din01[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END din01[0]
  PIN din01[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END din01[10]
  PIN din01[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END din01[11]
  PIN din01[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END din01[12]
  PIN din01[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END din01[13]
  PIN din01[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END din01[14]
  PIN din01[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END din01[15]
  PIN din01[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END din01[1]
  PIN din01[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END din01[2]
  PIN din01[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END din01[3]
  PIN din01[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END din01[4]
  PIN din01[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END din01[5]
  PIN din01[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END din01[6]
  PIN din01[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END din01[7]
  PIN din01[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END din01[8]
  PIN din01[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END din01[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 336.640 550.000 337.240 ;
    END
  END rst
  PIN sine_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END sine_out[0]
  PIN sine_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 363.840 550.000 364.440 ;
    END
  END sine_out[10]
  PIN sine_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 394.440 550.000 395.040 ;
    END
  END sine_out[11]
  PIN sine_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 391.040 550.000 391.640 ;
    END
  END sine_out[12]
  PIN sine_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 387.640 550.000 388.240 ;
    END
  END sine_out[13]
  PIN sine_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 380.840 550.000 381.440 ;
    END
  END sine_out[14]
  PIN sine_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 384.240 550.000 384.840 ;
    END
  END sine_out[15]
  PIN sine_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END sine_out[1]
  PIN sine_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END sine_out[2]
  PIN sine_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END sine_out[3]
  PIN sine_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END sine_out[4]
  PIN sine_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END sine_out[5]
  PIN sine_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 367.240 550.000 367.840 ;
    END
  END sine_out[6]
  PIN sine_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 370.640 550.000 371.240 ;
    END
  END sine_out[7]
  PIN sine_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 374.040 550.000 374.640 ;
    END
  END sine_out[8]
  PIN sine_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 546.000 377.440 550.000 378.040 ;
    END
  END sine_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 39.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 328.250 176.240 389.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 678.250 176.240 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 328.880 329.840 390.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 679.170 329.840 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 328.250 483.440 390.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 678.250 483.440 737.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 544.420 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 544.420 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 544.420 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 544.420 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 544.420 641.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 529.580 35.120 531.180 332.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 529.580 386.000 531.180 682.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 21.040 704.700 544.420 706.300 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 328.250 179.540 390.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 678.250 179.540 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 328.250 333.140 390.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 678.250 333.140 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 328.250 486.740 390.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 678.250 486.740 737.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 544.420 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 544.420 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 544.420 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 544.420 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 642.750 544.420 644.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 533.260 35.120 534.860 332.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 533.260 386.000 534.860 682.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 21.040 708.100 544.420 709.700 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 544.370 737.310 ;
      LAYER li1 ;
        RECT 5.520 10.795 544.180 737.205 ;
      LAYER met1 ;
        RECT 4.210 10.640 544.180 737.360 ;
      LAYER met2 ;
        RECT 4.230 4.280 542.710 737.305 ;
        RECT 4.230 4.000 80.310 4.280 ;
        RECT 81.150 4.000 157.590 4.280 ;
        RECT 158.430 4.000 164.030 4.280 ;
        RECT 164.870 4.000 170.470 4.280 ;
        RECT 171.310 4.000 176.910 4.280 ;
        RECT 177.750 4.000 180.130 4.280 ;
        RECT 180.970 4.000 186.570 4.280 ;
        RECT 187.410 4.000 193.010 4.280 ;
        RECT 193.850 4.000 199.450 4.280 ;
        RECT 200.290 4.000 205.890 4.280 ;
        RECT 206.730 4.000 209.110 4.280 ;
        RECT 209.950 4.000 215.550 4.280 ;
        RECT 216.390 4.000 542.710 4.280 ;
      LAYER met3 ;
        RECT 3.990 555.240 546.000 737.285 ;
        RECT 4.400 553.840 546.000 555.240 ;
        RECT 3.990 548.440 546.000 553.840 ;
        RECT 4.400 547.040 546.000 548.440 ;
        RECT 3.990 541.640 546.000 547.040 ;
        RECT 4.400 540.240 546.000 541.640 ;
        RECT 3.990 534.840 546.000 540.240 ;
        RECT 4.400 533.440 546.000 534.840 ;
        RECT 3.990 528.040 546.000 533.440 ;
        RECT 4.400 526.640 546.000 528.040 ;
        RECT 3.990 521.240 546.000 526.640 ;
        RECT 4.400 519.840 546.000 521.240 ;
        RECT 3.990 443.040 546.000 519.840 ;
        RECT 4.400 441.640 546.000 443.040 ;
        RECT 3.990 439.640 546.000 441.640 ;
        RECT 4.400 438.240 546.000 439.640 ;
        RECT 3.990 436.240 546.000 438.240 ;
        RECT 4.400 434.840 546.000 436.240 ;
        RECT 3.990 432.840 546.000 434.840 ;
        RECT 4.400 431.440 546.000 432.840 ;
        RECT 3.990 429.440 546.000 431.440 ;
        RECT 4.400 428.040 546.000 429.440 ;
        RECT 3.990 426.040 546.000 428.040 ;
        RECT 4.400 424.640 546.000 426.040 ;
        RECT 3.990 422.640 546.000 424.640 ;
        RECT 4.400 421.240 546.000 422.640 ;
        RECT 3.990 419.240 546.000 421.240 ;
        RECT 4.400 417.840 546.000 419.240 ;
        RECT 3.990 415.840 546.000 417.840 ;
        RECT 4.400 414.440 546.000 415.840 ;
        RECT 3.990 412.440 546.000 414.440 ;
        RECT 4.400 411.040 546.000 412.440 ;
        RECT 3.990 409.040 546.000 411.040 ;
        RECT 4.400 407.640 546.000 409.040 ;
        RECT 3.990 405.640 546.000 407.640 ;
        RECT 4.400 404.240 546.000 405.640 ;
        RECT 3.990 402.240 546.000 404.240 ;
        RECT 4.400 400.840 546.000 402.240 ;
        RECT 3.990 398.840 546.000 400.840 ;
        RECT 4.400 397.440 546.000 398.840 ;
        RECT 3.990 395.440 546.000 397.440 ;
        RECT 4.400 394.040 545.600 395.440 ;
        RECT 3.990 392.040 546.000 394.040 ;
        RECT 4.400 390.640 545.600 392.040 ;
        RECT 3.990 388.640 546.000 390.640 ;
        RECT 4.400 387.240 545.600 388.640 ;
        RECT 3.990 385.240 546.000 387.240 ;
        RECT 4.400 383.840 545.600 385.240 ;
        RECT 3.990 381.840 546.000 383.840 ;
        RECT 4.400 380.440 545.600 381.840 ;
        RECT 3.990 378.440 546.000 380.440 ;
        RECT 4.400 377.040 545.600 378.440 ;
        RECT 3.990 375.040 546.000 377.040 ;
        RECT 4.400 373.640 545.600 375.040 ;
        RECT 3.990 371.640 546.000 373.640 ;
        RECT 4.400 370.240 545.600 371.640 ;
        RECT 3.990 368.240 546.000 370.240 ;
        RECT 4.400 366.840 545.600 368.240 ;
        RECT 3.990 364.840 546.000 366.840 ;
        RECT 4.400 363.440 545.600 364.840 ;
        RECT 3.990 361.440 546.000 363.440 ;
        RECT 4.400 360.040 546.000 361.440 ;
        RECT 3.990 337.640 546.000 360.040 ;
        RECT 3.990 336.240 545.600 337.640 ;
        RECT 3.990 69.040 546.000 336.240 ;
        RECT 4.400 67.640 546.000 69.040 ;
        RECT 3.990 65.640 546.000 67.640 ;
        RECT 4.400 64.240 546.000 65.640 ;
        RECT 3.990 62.240 546.000 64.240 ;
        RECT 4.400 60.840 546.000 62.240 ;
        RECT 3.990 58.840 546.000 60.840 ;
        RECT 4.400 57.440 546.000 58.840 ;
        RECT 3.990 55.440 546.000 57.440 ;
        RECT 4.400 54.040 546.000 55.440 ;
        RECT 3.990 52.040 546.000 54.040 ;
        RECT 4.400 50.640 546.000 52.040 ;
        RECT 3.990 48.640 546.000 50.640 ;
        RECT 4.400 47.240 546.000 48.640 ;
        RECT 3.990 45.240 546.000 47.240 ;
        RECT 4.400 43.840 546.000 45.240 ;
        RECT 3.990 41.840 546.000 43.840 ;
        RECT 4.400 40.440 546.000 41.840 ;
        RECT 3.990 38.440 546.000 40.440 ;
        RECT 4.400 37.040 546.000 38.440 ;
        RECT 3.990 35.040 546.000 37.040 ;
        RECT 4.400 33.640 546.000 35.040 ;
        RECT 3.990 31.640 546.000 33.640 ;
        RECT 4.400 30.240 546.000 31.640 ;
        RECT 3.990 28.240 546.000 30.240 ;
        RECT 4.400 26.840 546.000 28.240 ;
        RECT 3.990 24.840 546.000 26.840 ;
        RECT 4.400 23.440 546.000 24.840 ;
        RECT 3.990 10.715 546.000 23.440 ;
      LAYER met4 ;
        RECT 50.000 390.720 509.900 676.425 ;
        RECT 50.000 389.800 177.540 390.720 ;
        RECT 50.000 327.850 174.240 389.800 ;
        RECT 176.640 327.850 177.540 389.800 ;
        RECT 179.940 328.480 327.840 390.720 ;
        RECT 330.240 328.480 331.140 390.720 ;
        RECT 179.940 327.850 331.140 328.480 ;
        RECT 333.540 327.850 481.440 390.720 ;
        RECT 483.840 327.850 484.740 390.720 ;
        RECT 487.140 327.850 509.900 390.720 ;
        RECT 50.000 40.720 509.900 327.850 ;
        RECT 50.000 39.800 177.540 40.720 ;
        RECT 50.000 22.615 174.240 39.800 ;
        RECT 176.640 22.615 177.540 39.800 ;
        RECT 179.940 22.615 327.840 40.720 ;
        RECT 330.240 22.615 331.140 40.720 ;
        RECT 333.540 22.615 481.440 40.720 ;
        RECT 483.840 22.615 484.740 40.720 ;
        RECT 487.140 22.615 509.900 40.720 ;
  END
END counter
END LIBRARY

