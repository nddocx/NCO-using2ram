module counter (clk,
    csb0,
    rst,
    addr0,
    din0,
    sine_out);
 input clk;
 input csb0;
 input rst;
 input [7:0] addr0;
 input [15:0] din0;
 output [15:0] sine_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire clknet_0_clk;
 wire \sine_out_temp[0] ;
 wire \sine_out_temp[10] ;
 wire \sine_out_temp[11] ;
 wire \sine_out_temp[12] ;
 wire \sine_out_temp[13] ;
 wire \sine_out_temp[14] ;
 wire \sine_out_temp[15] ;
 wire \sine_out_temp[1] ;
 wire \sine_out_temp[2] ;
 wire \sine_out_temp[3] ;
 wire \sine_out_temp[4] ;
 wire \sine_out_temp[5] ;
 wire \sine_out_temp[6] ;
 wire \sine_out_temp[7] ;
 wire \sine_out_temp[8] ;
 wire \sine_out_temp[9] ;
 wire \tcout[0] ;
 wire \tcout[1] ;
 wire \tcout[2] ;
 wire \tcout[3] ;
 wire \tcout[4] ;
 wire \tcout[5] ;
 wire \tcout[6] ;
 wire \tcout[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;

 sky130_fd_sc_hd__inv_2 _040_ (.A(net61),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _041_ (.A(net54),
    .Y(_008_));
 sky130_fd_sc_hd__xor2_1 _042_ (.A(\tcout[0] ),
    .B(net62),
    .X(_001_));
 sky130_fd_sc_hd__and3_2 _043_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .C(\tcout[2] ),
    .X(_032_));
 sky130_fd_sc_hd__a21oi_1 _044_ (.A1(\tcout[0] ),
    .A2(\tcout[1] ),
    .B1(net66),
    .Y(_033_));
 sky130_fd_sc_hd__nor2_1 _045_ (.A(_032_),
    .B(_033_),
    .Y(_002_));
 sky130_fd_sc_hd__nand2_1 _046_ (.A(net50),
    .B(_032_),
    .Y(_034_));
 sky130_fd_sc_hd__xor2_1 _047_ (.A(net59),
    .B(_032_),
    .X(_003_));
 sky130_fd_sc_hd__and3_1 _048_ (.A(net49),
    .B(net47),
    .C(_032_),
    .X(_035_));
 sky130_fd_sc_hd__xnor2_1 _049_ (.A(net60),
    .B(_034_),
    .Y(_004_));
 sky130_fd_sc_hd__and3_1 _050_ (.A(net49),
    .B(net47),
    .C(\tcout[5] ),
    .X(_036_));
 sky130_fd_sc_hd__o2bb2a_1 _051_ (.A1_N(_032_),
    .A2_N(_036_),
    .B1(_035_),
    .B2(net65),
    .X(_005_));
 sky130_fd_sc_hd__and3_1 _052_ (.A(\tcout[6] ),
    .B(_032_),
    .C(_036_),
    .X(_037_));
 sky130_fd_sc_hd__a21oi_1 _053_ (.A1(_032_),
    .A2(_036_),
    .B1(net64),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_1 _054_ (.A(_037_),
    .B(_038_),
    .Y(_006_));
 sky130_fd_sc_hd__xor2_1 _055_ (.A(net58),
    .B(_037_),
    .X(_007_));
 sky130_fd_sc_hd__inv_2 _056_ (.A(net54),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _057_ (.A(net54),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _058_ (.A(net54),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _059_ (.A(net54),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _060_ (.A(net54),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _061_ (.A(net54),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _062_ (.A(net55),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _063_ (.A(net55),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _064_ (.A(net55),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _065_ (.A(net55),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _066_ (.A(net55),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _067_ (.A(net55),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _068_ (.A(net56),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _069_ (.A(net56),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _070_ (.A(net56),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _071_ (.A(net56),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _072_ (.A(net56),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _073_ (.A(net56),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _074_ (.A(net56),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _075_ (.A(net56),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _076_ (.A(net54),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _077_ (.A(net54),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _078_ (.A(net54),
    .Y(_031_));
 sky130_fd_sc_hd__dfrtp_1 _079_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[3] ),
    .RESET_B(_008_),
    .Q(net36));
 sky130_fd_sc_hd__dfrtp_1 _080_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[4] ),
    .RESET_B(_009_),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_1 _081_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[5] ),
    .RESET_B(_010_),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_1 _082_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[6] ),
    .RESET_B(_011_),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_1 _083_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[7] ),
    .RESET_B(_012_),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_1 _084_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[8] ),
    .RESET_B(_013_),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _085_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[9] ),
    .RESET_B(_014_),
    .Q(net42));
 sky130_fd_sc_hd__dfrtp_1 _086_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[10] ),
    .RESET_B(_015_),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _087_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[11] ),
    .RESET_B(_016_),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _088_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[12] ),
    .RESET_B(_017_),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _089_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[13] ),
    .RESET_B(_018_),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _090_ (.CLK(clknet_1_1__leaf_clk),
    .D(\sine_out_temp[14] ),
    .RESET_B(_019_),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_1 _091_ (.CLK(clknet_1_1__leaf_clk),
    .D(\sine_out_temp[15] ),
    .RESET_B(_020_),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_4 _092_ (.CLK(clknet_1_1__leaf_clk),
    .D(_000_),
    .RESET_B(_021_),
    .Q(\tcout[0] ));
 sky130_fd_sc_hd__dfrtp_1 _093_ (.CLK(clknet_1_1__leaf_clk),
    .D(net63),
    .RESET_B(_022_),
    .Q(\tcout[1] ));
 sky130_fd_sc_hd__dfrtp_1 _094_ (.CLK(clknet_1_1__leaf_clk),
    .D(_002_),
    .RESET_B(_023_),
    .Q(\tcout[2] ));
 sky130_fd_sc_hd__dfrtp_1 _095_ (.CLK(clknet_1_1__leaf_clk),
    .D(_003_),
    .RESET_B(_024_),
    .Q(\tcout[3] ));
 sky130_fd_sc_hd__dfrtp_1 _096_ (.CLK(clknet_1_1__leaf_clk),
    .D(_004_),
    .RESET_B(_025_),
    .Q(\tcout[4] ));
 sky130_fd_sc_hd__dfrtp_1 _097_ (.CLK(clknet_1_1__leaf_clk),
    .D(_005_),
    .RESET_B(_026_),
    .Q(\tcout[5] ));
 sky130_fd_sc_hd__dfrtp_1 _098_ (.CLK(clknet_1_1__leaf_clk),
    .D(_006_),
    .RESET_B(_027_),
    .Q(\tcout[6] ));
 sky130_fd_sc_hd__dfrtp_1 _099_ (.CLK(clknet_1_1__leaf_clk),
    .D(_007_),
    .RESET_B(_028_),
    .Q(\tcout[7] ));
 sky130_fd_sc_hd__dfrtp_1 _100_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[0] ),
    .RESET_B(_029_),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_1 _101_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[1] ),
    .RESET_B(_030_),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_1 _102_ (.CLK(clknet_1_0__leaf_clk),
    .D(\sine_out_temp[2] ),
    .RESET_B(_031_),
    .Q(net35));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 ram_256x16 mem_i (.csb0(net9),
    .csb1(net57),
    .clk0(clknet_1_0__leaf_clk),
    .clk1(clknet_1_1__leaf_clk),
    .addr0({net8,
    net7,
    net6,
    net5,
    net4,
    net3,
    net2,
    net1}),
    .addr1({net43,
    net44,
    net45,
    net46,
    net48,
    net51,
    net52,
    net53}),
    .din0({net16,
    net15,
    net14,
    net13,
    net12,
    net11,
    net25,
    net24,
    net23,
    net22,
    net21,
    net20,
    net19,
    net18,
    net17,
    net10}),
    .dout1({\sine_out_temp[15] ,
    \sine_out_temp[14] ,
    \sine_out_temp[13] ,
    \sine_out_temp[12] ,
    \sine_out_temp[11] ,
    \sine_out_temp[10] ,
    \sine_out_temp[9] ,
    \sine_out_temp[8] ,
    \sine_out_temp[7] ,
    \sine_out_temp[6] ,
    \sine_out_temp[5] ,
    \sine_out_temp[4] ,
    \sine_out_temp[3] ,
    \sine_out_temp[2] ,
    \sine_out_temp[1] ,
    \sine_out_temp[0] }));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Right_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Right_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Right_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Right_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Right_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Right_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Right_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Right_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Right_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Right_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Right_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Right_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Right_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Right_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Right_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Right_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Right_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Right_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Right_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Right_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Right_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Right_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Right_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Right_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Right_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Right_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Right_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Right_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Right_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Right_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Right_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Right_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Right_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Right_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Right_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Right_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Right_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Right_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Right_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Right_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Right_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Right_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Right_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Right_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Right_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Right_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Right_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Right_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Right_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Right_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Right_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Right_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Right_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Right_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Right_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Right_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Right_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Right_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Right_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Right_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Right_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Right_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Right_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Right_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Right_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Right_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Right_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Right_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Right_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Right_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Right_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Right_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Right_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Right_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Right_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Right_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Right_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Right_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Right_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Right_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Right_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Right_444 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Right_445 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Right_446 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Right_447 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Right_448 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Right_449 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Right_450 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Right_451 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Right_452 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Right_453 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Right_454 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Right_455 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Right_456 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Right_457 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Right_458 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Right_459 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Right_460 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Right_461 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Right_462 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Right_463 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Right_464 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Right_465 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Right_466 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Right_467 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Right_468 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Right_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_2_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_2_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_2_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_2_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_2_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_2_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_2_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_2_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_2_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_2_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_2_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_2_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_2_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_2_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_2_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_2_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_2_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_2_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_2_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_2_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_2_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_1208 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(addr0[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(addr0[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(addr0[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(addr0[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(addr0[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(addr0[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(addr0[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(addr0[7]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(csb0),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(din0[0]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(din0[10]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(din0[11]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(din0[12]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(din0[13]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(din0[14]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(din0[15]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(din0[1]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(din0[2]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(din0[3]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(din0[4]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(din0[5]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(din0[6]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(din0[7]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(din0[8]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(din0[9]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(rst),
    .X(net26));
 sky130_fd_sc_hd__buf_1 output27 (.A(net27),
    .X(sine_out[0]));
 sky130_fd_sc_hd__buf_1 output28 (.A(net28),
    .X(sine_out[10]));
 sky130_fd_sc_hd__buf_1 output29 (.A(net29),
    .X(sine_out[11]));
 sky130_fd_sc_hd__buf_1 output30 (.A(net30),
    .X(sine_out[12]));
 sky130_fd_sc_hd__buf_1 output31 (.A(net31),
    .X(sine_out[13]));
 sky130_fd_sc_hd__buf_1 output32 (.A(net32),
    .X(sine_out[14]));
 sky130_fd_sc_hd__buf_1 output33 (.A(net33),
    .X(sine_out[15]));
 sky130_fd_sc_hd__buf_1 output34 (.A(net34),
    .X(sine_out[1]));
 sky130_fd_sc_hd__buf_1 output35 (.A(net35),
    .X(sine_out[2]));
 sky130_fd_sc_hd__buf_1 output36 (.A(net36),
    .X(sine_out[3]));
 sky130_fd_sc_hd__buf_1 output37 (.A(net37),
    .X(sine_out[4]));
 sky130_fd_sc_hd__buf_1 output38 (.A(net38),
    .X(sine_out[5]));
 sky130_fd_sc_hd__buf_1 output39 (.A(net39),
    .X(sine_out[6]));
 sky130_fd_sc_hd__buf_1 output40 (.A(net40),
    .X(sine_out[7]));
 sky130_fd_sc_hd__buf_1 output41 (.A(net41),
    .X(sine_out[8]));
 sky130_fd_sc_hd__buf_1 output42 (.A(net42),
    .X(sine_out[9]));
 sky130_fd_sc_hd__clkbuf_2 load_slew43 (.A(\tcout[7] ),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 load_slew44 (.A(\tcout[6] ),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 load_slew45 (.A(\tcout[5] ),
    .X(net45));
 sky130_fd_sc_hd__buf_1 load_slew46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__buf_1 load_slew47 (.A(\tcout[4] ),
    .X(net47));
 sky130_fd_sc_hd__buf_1 load_slew48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_1 load_slew49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 load_slew50 (.A(\tcout[3] ),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 load_slew51 (.A(\tcout[2] ),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 load_slew52 (.A(\tcout[1] ),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 load_slew53 (.A(\tcout[0] ),
    .X(net53));
 sky130_fd_sc_hd__buf_4 fanout54 (.A(net56),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_8 fanout56 (.A(net26),
    .X(net56));
 sky130_fd_sc_hd__conb_1 mem_i_57 (.LO(net57));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\tcout[7] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\tcout[3] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\tcout[4] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\tcout[0] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\tcout[1] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_001_),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\tcout[6] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\tcout[5] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\tcout[2] ),
    .X(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__092__RESET_B (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__Y (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__053__A1 (.DIODE(_032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__052__B (.DIODE(_032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__051__A1_N (.DIODE(_032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__048__C (.DIODE(_032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__047__B (.DIODE(_032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__046__B (.DIODE(_032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__045__A (.DIODE(_032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__043__X (.DIODE(_032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(addr0[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(addr0[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(addr0[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(addr0[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(addr0[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(addr0[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(addr0[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(addr0[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(csb0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(din0[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(din0[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(din0[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(din0[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(din0[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(din0[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(din0[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(din0[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(din0[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(din0[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(din0[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(din0[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(din0[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(din0[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(din0[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(din0[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew43_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i_addr1[7]  (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew44_X (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i_addr1[6]  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew45_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i_addr1[5]  (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew51_X (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i_addr1[2]  (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew52_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i_addr1[1]  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew53_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i_addr1[0]  (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_X (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__074__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__072__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__079__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__080__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__081__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__082__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__083__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__084__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__085__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__086__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__087__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__088__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__089__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__100__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__101__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__102__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i_clk0 (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_clk_X (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload0_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__090__CLK (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__091__CLK (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__092__CLK (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__CLK (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__094__CLK (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__095__CLK (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__096__CLK (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__097__CLK (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__098__CLK (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__099__CLK (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i_clk1 (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_clk_X (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\sine_out_temp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\sine_out_temp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\sine_out_temp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\sine_out_temp[3] ));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1122 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1189 ();
endmodule
