VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter
  CLASS BLOCK ;
  FOREIGN counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 800.000 ;
  PIN addr00[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END addr00[0]
  PIN addr00[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END addr00[1]
  PIN addr00[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END addr00[2]
  PIN addr00[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END addr00[3]
  PIN addr00[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END addr00[4]
  PIN addr00[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END addr00[5]
  PIN addr00[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END addr00[6]
  PIN addr00[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END addr00[7]
  PIN addr01[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END addr01[0]
  PIN addr01[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END addr01[1]
  PIN addr01[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END addr01[2]
  PIN addr01[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END addr01[3]
  PIN addr01[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END addr01[4]
  PIN addr01[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END addr01[5]
  PIN addr01[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END addr01[6]
  PIN addr01[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END addr01[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END clk
  PIN csb00
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END csb00
  PIN csb01
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END csb01
  PIN din00[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END din00[0]
  PIN din00[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END din00[10]
  PIN din00[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END din00[11]
  PIN din00[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END din00[12]
  PIN din00[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END din00[13]
  PIN din00[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END din00[14]
  PIN din00[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END din00[15]
  PIN din00[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END din00[1]
  PIN din00[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END din00[2]
  PIN din00[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END din00[3]
  PIN din00[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END din00[4]
  PIN din00[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END din00[5]
  PIN din00[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END din00[6]
  PIN din00[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END din00[7]
  PIN din00[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END din00[8]
  PIN din00[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END din00[9]
  PIN din01[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END din01[0]
  PIN din01[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END din01[10]
  PIN din01[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END din01[11]
  PIN din01[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END din01[12]
  PIN din01[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END din01[13]
  PIN din01[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END din01[14]
  PIN din01[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END din01[15]
  PIN din01[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END din01[1]
  PIN din01[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END din01[2]
  PIN din01[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END din01[3]
  PIN din01[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END din01[4]
  PIN din01[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END din01[5]
  PIN din01[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END din01[6]
  PIN din01[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END din01[7]
  PIN din01[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END din01[8]
  PIN din01[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END din01[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END rst
  PIN sine_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END sine_out[0]
  PIN sine_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END sine_out[10]
  PIN sine_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END sine_out[11]
  PIN sine_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END sine_out[12]
  PIN sine_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END sine_out[13]
  PIN sine_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END sine_out[14]
  PIN sine_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END sine_out[15]
  PIN sine_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END sine_out[1]
  PIN sine_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END sine_out[2]
  PIN sine_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END sine_out[3]
  PIN sine_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END sine_out[4]
  PIN sine_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END sine_out[5]
  PIN sine_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END sine_out[6]
  PIN sine_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END sine_out[7]
  PIN sine_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END sine_out[8]
  PIN sine_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END sine_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 39.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 328.250 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 328.880 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 328.250 483.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 328.250 790.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 328.880 944.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 328.250 1097.840 789.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 1194.400 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 1194.400 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 1194.400 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 1194.400 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 1194.400 641.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 1154.260 35.120 1155.860 332.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 328.250 179.540 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 328.250 333.140 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 328.250 486.740 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 39.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 329.170 793.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 10.640 947.540 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 328.250 947.540 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.540 10.640 1101.140 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.540 328.250 1101.140 789.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 1194.400 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 1194.400 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 1194.400 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 1194.400 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 642.750 1194.400 644.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 578.340 201.040 579.940 212.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1157.940 35.120 1159.540 332.080 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 1194.350 788.885 ;
      LAYER li1 ;
        RECT 5.520 10.795 1194.160 788.885 ;
      LAYER met1 ;
        RECT 5.520 0.380 1194.160 789.040 ;
      LAYER met2 ;
        RECT 6.070 4.280 1159.510 788.985 ;
        RECT 6.070 0.350 80.310 4.280 ;
        RECT 81.150 0.350 180.130 4.280 ;
        RECT 180.970 0.350 186.570 4.280 ;
        RECT 187.410 0.350 193.010 4.280 ;
        RECT 193.850 0.350 199.450 4.280 ;
        RECT 200.290 0.350 205.890 4.280 ;
        RECT 206.730 0.350 209.110 4.280 ;
        RECT 209.950 0.350 215.550 4.280 ;
        RECT 216.390 0.350 534.330 4.280 ;
        RECT 535.170 0.350 537.550 4.280 ;
        RECT 538.390 0.350 540.770 4.280 ;
        RECT 541.610 0.350 547.210 4.280 ;
        RECT 548.050 0.350 550.430 4.280 ;
        RECT 551.270 0.350 560.090 4.280 ;
        RECT 560.930 0.350 566.530 4.280 ;
        RECT 567.370 0.350 572.970 4.280 ;
        RECT 573.810 0.350 579.410 4.280 ;
        RECT 580.250 0.350 589.070 4.280 ;
        RECT 589.910 0.350 595.510 4.280 ;
        RECT 596.350 0.350 605.170 4.280 ;
        RECT 606.010 0.350 611.610 4.280 ;
        RECT 612.450 0.350 618.050 4.280 ;
        RECT 618.890 0.350 643.810 4.280 ;
        RECT 644.650 0.350 647.030 4.280 ;
        RECT 647.870 0.350 650.250 4.280 ;
        RECT 651.090 0.350 653.470 4.280 ;
        RECT 654.310 0.350 656.690 4.280 ;
        RECT 657.530 0.350 659.910 4.280 ;
        RECT 660.750 0.350 663.130 4.280 ;
        RECT 663.970 0.350 666.350 4.280 ;
        RECT 667.190 0.350 669.570 4.280 ;
        RECT 670.410 0.350 672.790 4.280 ;
        RECT 673.630 0.350 717.870 4.280 ;
        RECT 718.710 0.350 724.310 4.280 ;
        RECT 725.150 0.350 727.530 4.280 ;
        RECT 728.370 0.350 733.970 4.280 ;
        RECT 734.810 0.350 740.410 4.280 ;
        RECT 741.250 0.350 746.850 4.280 ;
        RECT 747.690 0.350 753.290 4.280 ;
        RECT 754.130 0.350 756.510 4.280 ;
        RECT 757.350 0.350 762.950 4.280 ;
        RECT 763.790 0.350 769.390 4.280 ;
        RECT 770.230 0.350 775.830 4.280 ;
        RECT 776.670 0.350 782.270 4.280 ;
        RECT 783.110 0.350 785.490 4.280 ;
        RECT 786.330 0.350 791.930 4.280 ;
        RECT 792.770 0.350 798.370 4.280 ;
        RECT 799.210 0.350 804.810 4.280 ;
        RECT 805.650 0.350 811.250 4.280 ;
        RECT 812.090 0.350 817.690 4.280 ;
        RECT 818.530 0.350 1159.510 4.280 ;
      LAYER met3 ;
        RECT 4.000 120.040 1159.530 788.965 ;
        RECT 4.400 118.640 1159.530 120.040 ;
        RECT 4.000 116.640 1159.530 118.640 ;
        RECT 4.400 115.240 1159.530 116.640 ;
        RECT 4.000 113.240 1159.530 115.240 ;
        RECT 4.400 111.840 1159.530 113.240 ;
        RECT 4.000 109.840 1159.530 111.840 ;
        RECT 4.400 108.440 1159.530 109.840 ;
        RECT 4.000 106.440 1159.530 108.440 ;
        RECT 4.400 105.040 1159.530 106.440 ;
        RECT 4.000 103.040 1159.530 105.040 ;
        RECT 4.400 101.640 1159.530 103.040 ;
        RECT 4.000 79.240 1159.530 101.640 ;
        RECT 4.400 77.840 1159.530 79.240 ;
        RECT 4.000 69.040 1159.530 77.840 ;
        RECT 4.400 67.640 1159.530 69.040 ;
        RECT 4.000 65.640 1159.530 67.640 ;
        RECT 4.400 64.240 1159.530 65.640 ;
        RECT 4.000 62.240 1159.530 64.240 ;
        RECT 4.400 60.840 1159.530 62.240 ;
        RECT 4.000 58.840 1159.530 60.840 ;
        RECT 4.400 57.440 1159.530 58.840 ;
        RECT 4.000 55.440 1159.530 57.440 ;
        RECT 4.400 54.040 1159.530 55.440 ;
        RECT 4.000 52.040 1159.530 54.040 ;
        RECT 4.400 50.640 1159.530 52.040 ;
        RECT 4.000 48.640 1159.530 50.640 ;
        RECT 4.400 47.240 1159.530 48.640 ;
        RECT 4.000 45.240 1159.530 47.240 ;
        RECT 4.400 43.840 1159.530 45.240 ;
        RECT 4.000 41.840 1159.530 43.840 ;
        RECT 4.400 40.440 1159.530 41.840 ;
        RECT 4.000 38.440 1159.530 40.440 ;
        RECT 4.400 37.040 1159.530 38.440 ;
        RECT 4.000 35.040 1159.530 37.040 ;
        RECT 4.400 33.640 1159.530 35.040 ;
        RECT 4.000 10.715 1159.530 33.640 ;
      LAYER met4 ;
        RECT 50.000 327.850 174.240 330.305 ;
        RECT 176.640 327.850 177.540 330.305 ;
        RECT 179.940 328.480 327.840 330.305 ;
        RECT 330.240 328.480 331.140 330.305 ;
        RECT 179.940 327.850 331.140 328.480 ;
        RECT 333.540 327.850 481.440 330.305 ;
        RECT 483.840 327.850 484.740 330.305 ;
        RECT 487.140 327.850 635.040 330.305 ;
        RECT 50.000 212.800 635.040 327.850 ;
        RECT 50.000 200.640 577.940 212.800 ;
        RECT 580.340 200.640 635.040 212.800 ;
        RECT 50.000 40.720 635.040 200.640 ;
        RECT 50.000 39.800 177.540 40.720 ;
        RECT 50.000 20.575 174.240 39.800 ;
        RECT 176.640 20.575 177.540 39.800 ;
        RECT 179.940 20.575 327.840 40.720 ;
        RECT 330.240 20.575 331.140 40.720 ;
        RECT 333.540 20.575 481.440 40.720 ;
        RECT 483.840 20.575 484.740 40.720 ;
        RECT 487.140 20.575 635.040 40.720 ;
        RECT 637.440 20.575 638.340 330.305 ;
        RECT 640.740 327.850 788.640 330.305 ;
        RECT 791.040 328.770 791.940 330.305 ;
        RECT 794.340 328.770 942.240 330.305 ;
        RECT 791.040 328.480 942.240 328.770 ;
        RECT 944.640 328.480 945.540 330.305 ;
        RECT 791.040 327.850 945.540 328.480 ;
        RECT 947.940 327.850 1095.840 330.305 ;
        RECT 1098.240 327.850 1099.140 330.305 ;
        RECT 1101.540 327.850 1109.900 330.305 ;
        RECT 640.740 40.720 1109.900 327.850 ;
        RECT 640.740 20.575 788.640 40.720 ;
        RECT 791.040 39.800 942.240 40.720 ;
        RECT 791.040 20.575 791.940 39.800 ;
        RECT 794.340 20.575 942.240 39.800 ;
        RECT 944.640 20.575 945.540 40.720 ;
        RECT 947.940 20.575 1095.840 40.720 ;
        RECT 1098.240 20.575 1099.140 40.720 ;
        RECT 1101.540 20.575 1109.900 40.720 ;
  END
END counter
END LIBRARY

