magic
tech sky130A
magscale 1 2
timestamp 1741102719
<< viali >>
rect 41797 126497 41831 126531
rect 41061 126429 41095 126463
rect 58633 126429 58667 126463
rect 58817 126429 58851 126463
rect 36093 126361 36127 126395
rect 36277 126361 36311 126395
rect 36369 126361 36403 126395
rect 37749 126361 37783 126395
rect 41337 126361 41371 126395
rect 45201 126361 45235 126395
rect 48513 126361 48547 126395
rect 49709 126361 49743 126395
rect 58449 126361 58483 126395
rect 59369 126361 59403 126395
rect 61853 126361 61887 126395
rect 63969 126361 64003 126395
rect 65717 126361 65751 126395
rect 66729 126361 66763 126395
rect 70317 126361 70351 126395
rect 71421 126361 71455 126395
rect 77309 126361 77343 126395
rect 77493 126361 77527 126395
rect 77677 126361 77711 126395
rect 37657 126293 37691 126327
rect 37933 126293 37967 126327
rect 40969 126293 41003 126327
rect 41429 126293 41463 126327
rect 41613 126293 41647 126327
rect 45109 126293 45143 126327
rect 45385 126293 45419 126327
rect 48421 126293 48455 126327
rect 48697 126293 48731 126327
rect 49617 126293 49651 126327
rect 49893 126293 49927 126327
rect 59461 126293 59495 126327
rect 59737 126293 59771 126327
rect 61945 126293 61979 126327
rect 62221 126293 62255 126327
rect 64061 126293 64095 126327
rect 64337 126293 64371 126327
rect 65809 126293 65843 126327
rect 65993 126293 66027 126327
rect 66821 126293 66855 126327
rect 67097 126293 67131 126327
rect 70409 126293 70443 126327
rect 70869 126293 70903 126327
rect 71513 126293 71547 126327
rect 71789 126293 71823 126327
rect 86325 126293 86359 126327
rect 87337 126293 87371 126327
rect 95985 126293 96019 126327
rect 104357 119901 104391 119935
rect 1593 101541 1627 101575
rect 1409 101405 1443 101439
rect 1685 101405 1719 101439
rect 1409 99841 1443 99875
rect 1685 99841 1719 99875
rect 1593 99705 1627 99739
rect 1409 98753 1443 98787
rect 1685 98753 1719 98787
rect 1593 98617 1627 98651
rect 1593 97189 1627 97223
rect 1409 97053 1443 97087
rect 1685 97053 1719 97087
rect 1593 96101 1627 96135
rect 1409 95965 1443 95999
rect 1685 95965 1719 95999
rect 1409 94401 1443 94435
rect 1685 94401 1719 94435
rect 1593 94265 1627 94299
rect 104449 86377 104483 86411
rect 104725 86377 104759 86411
rect 104541 86105 104575 86139
rect 104541 85697 104575 85731
rect 104633 85629 104667 85663
rect 104909 85561 104943 85595
rect 104449 85289 104483 85323
rect 104725 85289 104759 85323
rect 104541 85085 104575 85119
rect 104357 80257 104391 80291
rect 104633 80257 104667 80291
rect 104449 80053 104483 80087
rect 104541 79101 104575 79135
rect 104909 79101 104943 79135
rect 104725 79033 104759 79067
rect 104449 78965 104483 78999
rect 105001 78761 105035 78795
rect 104429 78625 104463 78659
rect 104633 78557 104667 78591
rect 104909 78557 104943 78591
rect 105185 78557 105219 78591
rect 105461 78557 105495 78591
rect 1501 78489 1535 78523
rect 1685 78489 1719 78523
rect 1869 78489 1903 78523
rect 104357 78489 104391 78523
rect 1961 78421 1995 78455
rect 104541 78421 104575 78455
rect 104725 78421 104759 78455
rect 105277 78421 105311 78455
rect 105553 78421 105587 78455
rect 1501 78081 1535 78115
rect 1961 78081 1995 78115
rect 104357 78081 104391 78115
rect 1685 77945 1719 77979
rect 1869 77945 1903 77979
rect 105645 77877 105679 77911
rect 106197 77877 106231 77911
rect 104357 77469 104391 77503
rect 105093 77469 105127 77503
rect 104909 77333 104943 77367
rect 1501 76993 1535 77027
rect 1961 76993 1995 77027
rect 1685 76857 1719 76891
rect 1869 76857 1903 76891
rect 1501 76313 1535 76347
rect 1685 76313 1719 76347
rect 1869 76313 1903 76347
rect 1961 76245 1995 76279
rect 1593 76041 1627 76075
rect 104357 76041 104391 76075
rect 106197 76041 106231 76075
rect 1409 75905 1443 75939
rect 1685 75905 1719 75939
rect 106105 75905 106139 75939
rect 105829 75837 105863 75871
rect 104541 75293 104575 75327
rect 1501 75225 1535 75259
rect 1685 75225 1719 75259
rect 1869 75225 1903 75259
rect 1961 75157 1995 75191
rect 104357 75157 104391 75191
rect 104633 75157 104667 75191
rect 1501 74137 1535 74171
rect 1961 74137 1995 74171
rect 1593 74069 1627 74103
rect 1869 74069 1903 74103
rect 1409 73729 1443 73763
rect 1961 73729 1995 73763
rect 1593 73593 1627 73627
rect 1869 73593 1903 73627
rect 1685 73185 1719 73219
rect 1869 73185 1903 73219
rect 1501 73049 1535 73083
rect 1961 73049 1995 73083
rect 1501 72641 1535 72675
rect 1961 72641 1995 72675
rect 1685 72505 1719 72539
rect 1869 72505 1903 72539
rect 1501 71553 1535 71587
rect 1961 71553 1995 71587
rect 1593 71349 1627 71383
rect 1869 71349 1903 71383
rect 1685 70941 1719 70975
rect 1869 70941 1903 70975
rect 1501 70873 1535 70907
rect 2145 70873 2179 70907
rect 2053 70805 2087 70839
rect 1961 70465 1995 70499
rect 2237 70397 2271 70431
rect 2421 70397 2455 70431
rect 108313 69853 108347 69887
rect 1501 69785 1535 69819
rect 1685 69785 1719 69819
rect 1869 69785 1903 69819
rect 1961 69717 1995 69751
rect 108129 69717 108163 69751
rect 108497 69717 108531 69751
rect 108129 68765 108163 68799
rect 108313 68765 108347 68799
rect 1501 68697 1535 68731
rect 1685 68697 1719 68731
rect 1869 68697 1903 68731
rect 1961 68629 1995 68663
rect 108497 68629 108531 68663
rect 1501 68289 1535 68323
rect 1961 68289 1995 68323
rect 105737 68289 105771 68323
rect 108313 68289 108347 68323
rect 1685 68153 1719 68187
rect 1869 68153 1903 68187
rect 105829 68153 105863 68187
rect 105553 68085 105587 68119
rect 108497 68085 108531 68119
rect 1593 67881 1627 67915
rect 1869 67881 1903 67915
rect 23489 67881 23523 67915
rect 24685 67881 24719 67915
rect 25881 67881 25915 67915
rect 26985 67881 27019 67915
rect 29561 67881 29595 67915
rect 30481 67881 30515 67915
rect 31769 67881 31803 67915
rect 32873 67881 32907 67915
rect 33977 67881 34011 67915
rect 35173 67881 35207 67915
rect 36369 67881 36403 67915
rect 37473 67881 37507 67915
rect 38669 67881 38703 67915
rect 39865 67881 39899 67915
rect 41061 67881 41095 67915
rect 42165 67881 42199 67915
rect 43361 67881 43395 67915
rect 69765 67881 69799 67915
rect 88349 67881 88383 67915
rect 88901 67881 88935 67915
rect 89177 67881 89211 67915
rect 90189 67881 90223 67915
rect 90649 67881 90683 67915
rect 91937 67881 91971 67915
rect 94283 67881 94317 67915
rect 96353 67881 96387 67915
rect 97181 67881 97215 67915
rect 90925 67813 90959 67847
rect 91385 67813 91419 67847
rect 95157 67813 95191 67847
rect 108497 67813 108531 67847
rect 28181 67745 28215 67779
rect 90373 67745 90407 67779
rect 92581 67745 92615 67779
rect 94053 67745 94087 67779
rect 95433 67745 95467 67779
rect 96997 67745 97031 67779
rect 29009 67677 29043 67711
rect 29101 67677 29135 67711
rect 87429 67677 87463 67711
rect 87521 67677 87555 67711
rect 88257 67677 88291 67711
rect 88809 67677 88843 67711
rect 89085 67677 89119 67711
rect 91109 67677 91143 67711
rect 91569 67677 91603 67711
rect 91845 67677 91879 67711
rect 93317 67677 93351 67711
rect 93501 67677 93535 67711
rect 93777 67677 93811 67711
rect 94973 67677 95007 67711
rect 95341 67677 95375 67711
rect 95617 67677 95651 67711
rect 96169 67653 96203 67687
rect 96629 67677 96663 67711
rect 108313 67677 108347 67711
rect 1501 67609 1535 67643
rect 1961 67609 1995 67643
rect 16221 67609 16255 67643
rect 28917 67609 28951 67643
rect 87613 67609 87647 67643
rect 90465 67609 90499 67643
rect 91753 67609 91787 67643
rect 92673 67609 92707 67643
rect 69489 67541 69523 67575
rect 69857 67541 69891 67575
rect 90665 67541 90699 67575
rect 90833 67541 90867 67575
rect 93685 67541 93719 67575
rect 95709 67541 95743 67575
rect 95801 67541 95835 67575
rect 95985 67541 96019 67575
rect 96721 67541 96755 67575
rect 1777 67337 1811 67371
rect 18889 67337 18923 67371
rect 20729 67337 20763 67371
rect 33241 67337 33275 67371
rect 34989 67337 35023 67371
rect 35357 67337 35391 67371
rect 35449 67337 35483 67371
rect 35817 67337 35851 67371
rect 38669 67337 38703 67371
rect 40785 67337 40819 67371
rect 44373 67337 44407 67371
rect 66453 67337 66487 67371
rect 67005 67337 67039 67371
rect 67465 67337 67499 67371
rect 70133 67337 70167 67371
rect 70961 67337 70995 67371
rect 71421 67337 71455 67371
rect 74089 67337 74123 67371
rect 75009 67337 75043 67371
rect 75377 67337 75411 67371
rect 75469 67337 75503 67371
rect 75837 67337 75871 67371
rect 94053 67337 94087 67371
rect 95893 67337 95927 67371
rect 97181 67337 97215 67371
rect 99665 67337 99699 67371
rect 99849 67337 99883 67371
rect 20361 67269 20395 67303
rect 40325 67269 40359 67303
rect 46673 67269 46707 67303
rect 47225 67269 47259 67303
rect 67557 67269 67591 67303
rect 67925 67269 67959 67303
rect 68477 67269 68511 67303
rect 71053 67269 71087 67303
rect 74273 67269 74307 67303
rect 77033 67269 77067 67303
rect 87797 67269 87831 67303
rect 91569 67269 91603 67303
rect 101781 67269 101815 67303
rect 101965 67269 101999 67303
rect 1593 67201 1627 67235
rect 30389 67201 30423 67235
rect 30665 67201 30699 67235
rect 30757 67201 30791 67235
rect 30941 67201 30975 67235
rect 33609 67201 33643 67235
rect 33701 67201 33735 67235
rect 34069 67201 34103 67235
rect 39037 67201 39071 67235
rect 39497 67201 39531 67235
rect 39773 67201 39807 67235
rect 41245 67201 41279 67235
rect 46581 67201 46615 67235
rect 62037 67201 62071 67235
rect 62405 67201 62439 67235
rect 67097 67201 67131 67235
rect 68569 67201 68603 67235
rect 70225 67201 70259 67235
rect 71789 67201 71823 67235
rect 71881 67201 71915 67235
rect 72341 67201 72375 67235
rect 73169 67201 73203 67235
rect 73629 67201 73663 67235
rect 73721 67201 73755 67235
rect 76205 67201 76239 67235
rect 76573 67201 76607 67235
rect 76941 67201 76975 67235
rect 77309 67201 77343 67235
rect 79333 67201 79367 67235
rect 87153 67201 87187 67235
rect 87705 67201 87739 67235
rect 88073 67201 88107 67235
rect 88441 67201 88475 67235
rect 88625 67201 88659 67235
rect 89269 67201 89303 67235
rect 91201 67201 91235 67235
rect 91385 67201 91419 67235
rect 92029 67201 92063 67235
rect 95985 67201 96019 67235
rect 96169 67201 96203 67235
rect 98929 67201 98963 67235
rect 99205 67201 99239 67235
rect 99481 67201 99515 67235
rect 108313 67201 108347 67235
rect 20637 67133 20671 67167
rect 24777 67133 24811 67167
rect 25053 67133 25087 67167
rect 33885 67133 33919 67167
rect 34345 67133 34379 67167
rect 35633 67133 35667 67167
rect 39129 67133 39163 67167
rect 39313 67133 39347 67167
rect 40417 67133 40451 67167
rect 40601 67133 40635 67167
rect 44465 67133 44499 67167
rect 44557 67133 44591 67167
rect 45017 67133 45051 67167
rect 46857 67133 46891 67167
rect 47685 67133 47719 67167
rect 66821 67133 66855 67167
rect 68293 67133 68327 67167
rect 69673 67133 69707 67167
rect 69949 67133 69983 67167
rect 70869 67133 70903 67167
rect 71697 67133 71731 67167
rect 73537 67133 73571 67167
rect 75285 67133 75319 67167
rect 85313 67133 85347 67167
rect 85589 67133 85623 67167
rect 87245 67133 87279 67167
rect 90925 67133 90959 67167
rect 92305 67133 92339 67167
rect 93777 67133 93811 67167
rect 94145 67133 94179 67167
rect 94421 67133 94455 67167
rect 96077 67133 96111 67167
rect 98653 67133 98687 67167
rect 36093 67065 36127 67099
rect 44833 67065 44867 67099
rect 60749 67065 60783 67099
rect 62221 67065 62255 67099
rect 66545 67065 66579 67099
rect 68937 67065 68971 67099
rect 70593 67065 70627 67099
rect 72249 67065 72283 67099
rect 76297 67065 76331 67099
rect 88809 67065 88843 67099
rect 89453 67065 89487 67099
rect 99389 67065 99423 67099
rect 1409 66997 1443 67031
rect 20913 66997 20947 67031
rect 21281 66997 21315 67031
rect 23121 66997 23155 67031
rect 23305 66997 23339 67031
rect 25145 66997 25179 67031
rect 30297 66997 30331 67031
rect 30573 66997 30607 67031
rect 33149 66997 33183 67031
rect 39957 66997 39991 67031
rect 40969 66997 41003 67031
rect 44005 66997 44039 67031
rect 46213 66997 46247 67031
rect 47041 66997 47075 67031
rect 69489 66997 69523 67031
rect 79149 66997 79183 67031
rect 87061 66997 87095 67031
rect 87521 66997 87555 67031
rect 88165 66997 88199 67031
rect 96261 66997 96295 67031
rect 96537 66997 96571 67031
rect 108129 66997 108163 67031
rect 108497 66997 108531 67031
rect 29009 66793 29043 66827
rect 29745 66793 29779 66827
rect 31603 66793 31637 66827
rect 68017 66793 68051 66827
rect 82994 66793 83028 66827
rect 91642 66793 91676 66827
rect 94973 66793 95007 66827
rect 96169 66793 96203 66827
rect 96997 66793 97031 66827
rect 99573 66793 99607 66827
rect 22477 66725 22511 66759
rect 27077 66725 27111 66759
rect 32781 66725 32815 66759
rect 34253 66725 34287 66759
rect 70869 66725 70903 66759
rect 71421 66725 71455 66759
rect 82553 66725 82587 66759
rect 93133 66725 93167 66759
rect 17325 66657 17359 66691
rect 17601 66657 17635 66691
rect 22201 66657 22235 66691
rect 24225 66657 24259 66691
rect 24409 66657 24443 66691
rect 28549 66657 28583 66691
rect 28825 66657 28859 66691
rect 29377 66657 29411 66691
rect 31861 66657 31895 66691
rect 32229 66657 32263 66691
rect 33609 66657 33643 66691
rect 33793 66657 33827 66691
rect 68661 66657 68695 66691
rect 69213 66657 69247 66691
rect 79333 66657 79367 66691
rect 79425 66657 79459 66691
rect 79885 66657 79919 66691
rect 82737 66657 82771 66691
rect 84485 66657 84519 66691
rect 84853 66657 84887 66691
rect 85221 66657 85255 66691
rect 85405 66657 85439 66691
rect 86233 66657 86267 66691
rect 88336 66657 88370 66691
rect 90925 66657 90959 66691
rect 91385 66657 91419 66691
rect 95341 66657 95375 66691
rect 95985 66657 96019 66691
rect 17417 66589 17451 66623
rect 22385 66589 22419 66623
rect 29101 66589 29135 66623
rect 29561 66589 29595 66623
rect 32965 66589 32999 66623
rect 33057 66589 33091 66623
rect 33517 66589 33551 66623
rect 56793 66589 56827 66623
rect 70317 66589 70351 66623
rect 79793 66589 79827 66623
rect 84669 66589 84703 66623
rect 88073 66589 88107 66623
rect 90097 66589 90131 66623
rect 90189 66589 90223 66623
rect 93225 66589 93259 66623
rect 95525 66589 95559 66623
rect 95617 66589 95651 66623
rect 96813 66589 96847 66623
rect 98193 66589 98227 66623
rect 98469 66589 98503 66623
rect 101781 66589 101815 66623
rect 102057 66589 102091 66623
rect 102149 66589 102183 66623
rect 102241 66589 102275 66623
rect 21925 66521 21959 66555
rect 24685 66521 24719 66555
rect 69397 66521 69431 66555
rect 70041 66521 70075 66555
rect 77401 66521 77435 66555
rect 79057 66521 79091 66555
rect 86509 66521 86543 66555
rect 90005 66521 90039 66555
rect 90557 66521 90591 66555
rect 93501 66521 93535 66555
rect 95157 66521 95191 66555
rect 99205 66521 99239 66555
rect 99389 66521 99423 66555
rect 101965 66521 101999 66555
rect 102333 66521 102367 66555
rect 20269 66453 20303 66487
rect 20453 66453 20487 66487
rect 26157 66453 26191 66487
rect 26249 66453 26283 66487
rect 30113 66453 30147 66487
rect 31953 66453 31987 66487
rect 33149 66453 33183 66487
rect 33977 66453 34011 66487
rect 57069 66453 57103 66487
rect 68937 66453 68971 66487
rect 69305 66453 69339 66487
rect 69765 66453 69799 66487
rect 70409 66453 70443 66487
rect 77585 66453 77619 66487
rect 80161 66453 80195 66487
rect 84945 66453 84979 66487
rect 85497 66453 85531 66487
rect 85865 66453 85899 66487
rect 87981 66453 88015 66487
rect 89821 66453 89855 66487
rect 90281 66453 90315 66487
rect 90741 66453 90775 66487
rect 95801 66453 95835 66487
rect 96261 66453 96295 66487
rect 96629 66453 96663 66487
rect 99757 66453 99791 66487
rect 21925 66249 21959 66283
rect 28917 66249 28951 66283
rect 88533 66249 88567 66283
rect 92121 66249 92155 66283
rect 93317 66249 93351 66283
rect 98285 66249 98319 66283
rect 98561 66249 98595 66283
rect 100033 66249 100067 66283
rect 21373 66181 21407 66215
rect 21557 66181 21591 66215
rect 22293 66181 22327 66215
rect 31033 66181 31067 66215
rect 31217 66181 31251 66215
rect 57713 66181 57747 66215
rect 58081 66181 58115 66215
rect 83381 66181 83415 66215
rect 86325 66181 86359 66215
rect 89729 66181 89763 66215
rect 92397 66181 92431 66215
rect 94053 66181 94087 66215
rect 96077 66181 96111 66215
rect 98377 66181 98411 66215
rect 1593 66113 1627 66147
rect 1777 66113 1811 66147
rect 17877 66113 17911 66147
rect 19349 66113 19383 66147
rect 19441 66113 19475 66147
rect 21189 66113 21223 66147
rect 31125 66113 31159 66147
rect 55965 66113 55999 66147
rect 57989 66113 58023 66147
rect 83657 66113 83691 66147
rect 86417 66113 86451 66147
rect 86693 66113 86727 66147
rect 89085 66113 89119 66147
rect 89361 66113 89395 66147
rect 89453 66113 89487 66147
rect 91569 66113 91603 66147
rect 93961 66113 93995 66147
rect 94329 66113 94363 66147
rect 96353 66113 96387 66147
rect 96537 66113 96571 66147
rect 98653 66113 98687 66147
rect 98745 66113 98779 66147
rect 99113 66113 99147 66147
rect 100217 66113 100251 66147
rect 100401 66113 100435 66147
rect 108313 66113 108347 66147
rect 22017 66045 22051 66079
rect 23765 66045 23799 66079
rect 23857 66045 23891 66079
rect 83933 66045 83967 66079
rect 86969 66045 87003 66079
rect 91661 66045 91695 66079
rect 91937 66045 91971 66079
rect 92857 66045 92891 66079
rect 99389 66045 99423 66079
rect 92213 65977 92247 66011
rect 92765 65977 92799 66011
rect 94513 65977 94547 66011
rect 100401 65977 100435 66011
rect 108497 65977 108531 66011
rect 1409 65909 1443 65943
rect 53665 65909 53699 65943
rect 85405 65909 85439 65943
rect 85589 65909 85623 65943
rect 86509 65909 86543 65943
rect 88441 65909 88475 65943
rect 91201 65909 91235 65943
rect 93041 65909 93075 65943
rect 93501 65909 93535 65943
rect 94605 65909 94639 65943
rect 96800 65909 96834 65943
rect 98377 65909 98411 65943
rect 100585 65909 100619 65943
rect 100769 65909 100803 65943
rect 1593 65501 1627 65535
rect 1777 65501 1811 65535
rect 108129 65501 108163 65535
rect 108313 65501 108347 65535
rect 1409 65365 1443 65399
rect 108497 65365 108531 65399
rect 1593 65025 1627 65059
rect 108129 65025 108163 65059
rect 108313 65025 108347 65059
rect 1409 64889 1443 64923
rect 1777 64889 1811 64923
rect 108497 64889 108531 64923
rect 1593 64413 1627 64447
rect 1777 64413 1811 64447
rect 108129 64413 108163 64447
rect 108313 64413 108347 64447
rect 1409 64277 1443 64311
rect 108497 64277 108531 64311
rect 1409 63461 1443 63495
rect 1777 63461 1811 63495
rect 1593 63325 1627 63359
rect 1777 62985 1811 63019
rect 1593 62849 1627 62883
rect 1409 62713 1443 62747
rect 1593 62441 1627 62475
rect 1869 62441 1903 62475
rect 1501 62169 1535 62203
rect 1961 62169 1995 62203
rect 1685 61829 1719 61863
rect 1777 61829 1811 61863
rect 1501 61761 1535 61795
rect 1961 61761 1995 61795
rect 104357 60061 104391 60095
rect 104449 59721 104483 59755
rect 104357 59585 104391 59619
rect 104541 59585 104575 59619
rect 105645 58633 105679 58667
rect 106197 58633 106231 58667
rect 104357 58565 104391 58599
rect 104357 58089 104391 58123
rect 104541 57545 104575 57579
rect 104357 57477 104391 57511
rect 105001 57001 105035 57035
rect 105277 57001 105311 57035
rect 104357 56865 104391 56899
rect 104725 56865 104759 56899
rect 104817 56865 104851 56899
rect 105093 56865 105127 56899
rect 104449 56661 104483 56695
rect 104541 56661 104575 56695
rect 104725 56457 104759 56491
rect 104633 56389 104667 56423
rect 104909 56389 104943 56423
rect 104449 56321 104483 56355
rect 104449 55369 104483 55403
rect 104909 55369 104943 55403
rect 104725 55301 104759 55335
rect 104633 55233 104667 55267
rect 104909 54825 104943 54859
rect 105277 54825 105311 54859
rect 104357 54757 104391 54791
rect 104541 54621 104575 54655
rect 105093 54553 105127 54587
rect 104633 54485 104667 54519
rect 104725 54485 104759 54519
rect 104449 54281 104483 54315
rect 104541 54281 104575 54315
rect 104449 52105 104483 52139
rect 104541 51561 104575 51595
rect 104725 51493 104759 51527
rect 105185 51357 105219 51391
rect 108221 51357 108255 51391
rect 108497 51357 108531 51391
rect 104357 51289 104391 51323
rect 104909 51289 104943 51323
rect 105093 51289 105127 51323
rect 104557 51221 104591 51255
rect 105369 51221 105403 51255
rect 108313 51221 108347 51255
rect 104449 51017 104483 51051
rect 104541 51017 104575 51051
rect 104725 49929 104759 49963
rect 105001 49861 105035 49895
rect 105185 49861 105219 49895
rect 104357 49793 104391 49827
rect 104541 49793 104575 49827
rect 104817 49725 104851 49759
rect 105369 49725 105403 49759
rect 104357 49385 104391 49419
rect 104357 46121 104391 46155
rect 104541 45917 104575 45951
rect 104725 45441 104759 45475
rect 104633 45373 104667 45407
rect 104357 45237 104391 45271
rect 104449 44897 104483 44931
rect 105185 44897 105219 44931
rect 105001 44829 105035 44863
rect 105553 44421 105587 44455
rect 104357 44353 104391 44387
rect 105093 44353 105127 44387
rect 105185 44353 105219 44387
rect 105369 44353 105403 44387
rect 104541 44285 104575 44319
rect 105001 44149 105035 44183
rect 105093 42313 105127 42347
rect 104449 42177 104483 42211
rect 1593 41701 1627 41735
rect 1409 41565 1443 41599
rect 1685 41565 1719 41599
rect 1593 40137 1627 40171
rect 1409 40001 1443 40035
rect 1685 40001 1719 40035
rect 1593 38437 1627 38471
rect 1409 38301 1443 38335
rect 1685 38301 1719 38335
rect 104357 37961 104391 37995
rect 106197 37961 106231 37995
rect 106105 37825 106139 37859
rect 105829 37757 105863 37791
rect 104633 37281 104667 37315
rect 104725 37281 104759 37315
rect 1409 37213 1443 37247
rect 1685 37213 1719 37247
rect 104449 37213 104483 37247
rect 1593 37077 1627 37111
rect 1593 35785 1627 35819
rect 1409 35649 1443 35683
rect 1685 35649 1719 35683
rect 1593 34697 1627 34731
rect 1409 34561 1443 34595
rect 1685 34561 1719 34595
rect 104357 25109 104391 25143
rect 104357 23817 104391 23851
rect 104357 22729 104391 22763
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 1593 15929 1627 15963
rect 16129 7497 16163 7531
rect 90649 7497 90683 7531
rect 90741 7497 90775 7531
rect 91017 7497 91051 7531
rect 23489 2601 23523 2635
rect 24777 2601 24811 2635
rect 25881 2601 25915 2635
rect 27169 2601 27203 2635
rect 28457 2601 28491 2635
rect 29285 2601 29319 2635
rect 30573 2601 30607 2635
rect 31677 2601 31711 2635
rect 32965 2601 32999 2635
rect 34253 2601 34287 2635
rect 35541 2601 35575 2635
rect 36369 2601 36403 2635
rect 37473 2601 37507 2635
rect 38761 2601 38795 2635
rect 40049 2601 40083 2635
rect 41337 2601 41371 2635
rect 42165 2601 42199 2635
rect 43453 2601 43487 2635
rect 23305 2397 23339 2431
rect 24593 2397 24627 2431
rect 26065 2397 26099 2431
rect 27353 2397 27387 2431
rect 28641 2397 28675 2431
rect 29101 2397 29135 2431
rect 30389 2397 30423 2431
rect 31861 2397 31895 2431
rect 33149 2397 33183 2431
rect 34437 2397 34471 2431
rect 35725 2397 35759 2431
rect 36185 2397 36219 2431
rect 37657 2397 37691 2431
rect 38945 2397 38979 2431
rect 40233 2397 40267 2431
rect 41521 2397 41555 2431
rect 41981 2397 42015 2431
rect 43269 2397 43303 2431
rect 23213 2261 23247 2295
rect 24501 2261 24535 2295
rect 25789 2261 25823 2295
rect 27077 2261 27111 2295
rect 28365 2261 28399 2295
rect 29009 2261 29043 2295
rect 30297 2261 30331 2295
rect 31585 2261 31619 2295
rect 32873 2261 32907 2295
rect 34161 2261 34195 2295
rect 35449 2261 35483 2295
rect 36093 2261 36127 2295
rect 37381 2261 37415 2295
rect 38669 2261 38703 2295
rect 39957 2261 39991 2295
rect 41245 2261 41279 2295
rect 41889 2261 41923 2295
rect 43177 2261 43211 2295
<< metal1 >>
rect 98546 128324 98552 128376
rect 98604 128364 98610 128376
rect 102134 128364 102140 128376
rect 98604 128336 102140 128364
rect 98604 128324 98610 128336
rect 102134 128324 102140 128336
rect 102192 128324 102198 128376
rect 1104 127322 108836 127344
rect 1104 127270 4874 127322
rect 4926 127270 4938 127322
rect 4990 127270 5002 127322
rect 5054 127270 5066 127322
rect 5118 127270 5130 127322
rect 5182 127270 35594 127322
rect 35646 127270 35658 127322
rect 35710 127270 35722 127322
rect 35774 127270 35786 127322
rect 35838 127270 35850 127322
rect 35902 127270 66314 127322
rect 66366 127270 66378 127322
rect 66430 127270 66442 127322
rect 66494 127270 66506 127322
rect 66558 127270 66570 127322
rect 66622 127270 97034 127322
rect 97086 127270 97098 127322
rect 97150 127270 97162 127322
rect 97214 127270 97226 127322
rect 97278 127270 97290 127322
rect 97342 127270 108836 127322
rect 1104 127248 108836 127270
rect 1104 126778 108836 126800
rect 1104 126726 4214 126778
rect 4266 126726 4278 126778
rect 4330 126726 4342 126778
rect 4394 126726 4406 126778
rect 4458 126726 4470 126778
rect 4522 126726 34934 126778
rect 34986 126726 34998 126778
rect 35050 126726 35062 126778
rect 35114 126726 35126 126778
rect 35178 126726 35190 126778
rect 35242 126726 65654 126778
rect 65706 126726 65718 126778
rect 65770 126726 65782 126778
rect 65834 126726 65846 126778
rect 65898 126726 65910 126778
rect 65962 126726 96374 126778
rect 96426 126726 96438 126778
rect 96490 126726 96502 126778
rect 96554 126726 96566 126778
rect 96618 126726 96630 126778
rect 96682 126726 105922 126778
rect 105974 126726 105986 126778
rect 106038 126726 106050 126778
rect 106102 126726 106114 126778
rect 106166 126726 106178 126778
rect 106230 126726 108836 126778
rect 1104 126704 108836 126726
rect 41785 126531 41843 126537
rect 41785 126528 41797 126531
rect 40972 126500 41797 126528
rect 36078 126352 36084 126404
rect 36136 126352 36142 126404
rect 36262 126352 36268 126404
rect 36320 126392 36326 126404
rect 36357 126395 36415 126401
rect 36357 126392 36369 126395
rect 36320 126364 36369 126392
rect 36320 126352 36326 126364
rect 36357 126361 36369 126364
rect 36403 126361 36415 126395
rect 36357 126355 36415 126361
rect 37734 126352 37740 126404
rect 37792 126352 37798 126404
rect 40972 126336 41000 126500
rect 41785 126497 41797 126500
rect 41831 126497 41843 126531
rect 41785 126491 41843 126497
rect 41049 126463 41107 126469
rect 41049 126429 41061 126463
rect 41095 126460 41107 126463
rect 42334 126460 42340 126472
rect 41095 126432 42340 126460
rect 41095 126429 41107 126432
rect 41049 126423 41107 126429
rect 42334 126420 42340 126432
rect 42392 126420 42398 126472
rect 58621 126463 58679 126469
rect 58621 126429 58633 126463
rect 58667 126460 58679 126463
rect 58805 126463 58863 126469
rect 58805 126460 58817 126463
rect 58667 126432 58817 126460
rect 58667 126429 58679 126432
rect 58621 126423 58679 126429
rect 58805 126429 58817 126432
rect 58851 126460 58863 126463
rect 102594 126460 102600 126472
rect 58851 126432 102600 126460
rect 58851 126429 58863 126432
rect 58805 126423 58863 126429
rect 102594 126420 102600 126432
rect 102652 126420 102658 126472
rect 41322 126352 41328 126404
rect 41380 126352 41386 126404
rect 45186 126352 45192 126404
rect 45244 126352 45250 126404
rect 48498 126352 48504 126404
rect 48556 126352 48562 126404
rect 49694 126352 49700 126404
rect 49752 126352 49758 126404
rect 56778 126352 56784 126404
rect 56836 126392 56842 126404
rect 58437 126395 58495 126401
rect 58437 126392 58449 126395
rect 56836 126364 58449 126392
rect 56836 126352 56842 126364
rect 58437 126361 58449 126364
rect 58483 126361 58495 126395
rect 58437 126355 58495 126361
rect 59354 126352 59360 126404
rect 59412 126352 59418 126404
rect 61838 126352 61844 126404
rect 61896 126352 61902 126404
rect 63954 126352 63960 126404
rect 64012 126352 64018 126404
rect 64414 126352 64420 126404
rect 64472 126392 64478 126404
rect 65705 126395 65763 126401
rect 65705 126392 65717 126395
rect 64472 126364 65717 126392
rect 64472 126352 64478 126364
rect 65705 126361 65717 126364
rect 65751 126361 65763 126395
rect 65705 126355 65763 126361
rect 66070 126352 66076 126404
rect 66128 126392 66134 126404
rect 66717 126395 66775 126401
rect 66717 126392 66729 126395
rect 66128 126364 66729 126392
rect 66128 126352 66134 126364
rect 66717 126361 66729 126364
rect 66763 126361 66775 126395
rect 66717 126355 66775 126361
rect 68554 126352 68560 126404
rect 68612 126392 68618 126404
rect 70305 126395 70363 126401
rect 70305 126392 70317 126395
rect 68612 126364 70317 126392
rect 68612 126352 68618 126364
rect 70305 126361 70317 126364
rect 70351 126361 70363 126395
rect 70305 126355 70363 126361
rect 71406 126352 71412 126404
rect 71464 126352 71470 126404
rect 77294 126352 77300 126404
rect 77352 126352 77358 126404
rect 77481 126395 77539 126401
rect 77481 126361 77493 126395
rect 77527 126392 77539 126395
rect 77665 126395 77723 126401
rect 77665 126392 77677 126395
rect 77527 126364 77677 126392
rect 77527 126361 77539 126364
rect 77481 126355 77539 126361
rect 77665 126361 77677 126364
rect 77711 126392 77723 126395
rect 102318 126392 102324 126404
rect 77711 126364 102324 126392
rect 77711 126361 77723 126364
rect 77665 126355 77723 126361
rect 102318 126352 102324 126364
rect 102376 126352 102382 126404
rect 37642 126284 37648 126336
rect 37700 126324 37706 126336
rect 37921 126327 37979 126333
rect 37921 126324 37933 126327
rect 37700 126296 37933 126324
rect 37700 126284 37706 126296
rect 37921 126293 37933 126296
rect 37967 126293 37979 126327
rect 37921 126287 37979 126293
rect 40954 126284 40960 126336
rect 41012 126284 41018 126336
rect 41414 126284 41420 126336
rect 41472 126324 41478 126336
rect 41601 126327 41659 126333
rect 41601 126324 41613 126327
rect 41472 126296 41613 126324
rect 41472 126284 41478 126296
rect 41601 126293 41613 126296
rect 41647 126293 41659 126327
rect 41601 126287 41659 126293
rect 45094 126284 45100 126336
rect 45152 126324 45158 126336
rect 45373 126327 45431 126333
rect 45373 126324 45385 126327
rect 45152 126296 45385 126324
rect 45152 126284 45158 126296
rect 45373 126293 45385 126296
rect 45419 126293 45431 126327
rect 45373 126287 45431 126293
rect 48406 126284 48412 126336
rect 48464 126324 48470 126336
rect 48685 126327 48743 126333
rect 48685 126324 48697 126327
rect 48464 126296 48697 126324
rect 48464 126284 48470 126296
rect 48685 126293 48697 126296
rect 48731 126293 48743 126327
rect 48685 126287 48743 126293
rect 49602 126284 49608 126336
rect 49660 126324 49666 126336
rect 49881 126327 49939 126333
rect 49881 126324 49893 126327
rect 49660 126296 49893 126324
rect 49660 126284 49666 126296
rect 49881 126293 49893 126296
rect 49927 126293 49939 126327
rect 49881 126287 49939 126293
rect 59449 126327 59507 126333
rect 59449 126293 59461 126327
rect 59495 126324 59507 126327
rect 59722 126324 59728 126336
rect 59495 126296 59728 126324
rect 59495 126293 59507 126296
rect 59449 126287 59507 126293
rect 59722 126284 59728 126296
rect 59780 126284 59786 126336
rect 61933 126327 61991 126333
rect 61933 126293 61945 126327
rect 61979 126324 61991 126327
rect 62206 126324 62212 126336
rect 61979 126296 62212 126324
rect 61979 126293 61991 126296
rect 61933 126287 61991 126293
rect 62206 126284 62212 126296
rect 62264 126284 62270 126336
rect 64049 126327 64107 126333
rect 64049 126293 64061 126327
rect 64095 126324 64107 126327
rect 64322 126324 64328 126336
rect 64095 126296 64328 126324
rect 64095 126293 64107 126296
rect 64049 126287 64107 126293
rect 64322 126284 64328 126296
rect 64380 126284 64386 126336
rect 65797 126327 65855 126333
rect 65797 126293 65809 126327
rect 65843 126324 65855 126327
rect 65978 126324 65984 126336
rect 65843 126296 65984 126324
rect 65843 126293 65855 126296
rect 65797 126287 65855 126293
rect 65978 126284 65984 126296
rect 66036 126284 66042 126336
rect 66809 126327 66867 126333
rect 66809 126293 66821 126327
rect 66855 126324 66867 126327
rect 67082 126324 67088 126336
rect 66855 126296 67088 126324
rect 66855 126293 66867 126296
rect 66809 126287 66867 126293
rect 67082 126284 67088 126296
rect 67140 126284 67146 126336
rect 70397 126327 70455 126333
rect 70397 126293 70409 126327
rect 70443 126324 70455 126327
rect 70854 126324 70860 126336
rect 70443 126296 70860 126324
rect 70443 126293 70455 126296
rect 70397 126287 70455 126293
rect 70854 126284 70860 126296
rect 70912 126284 70918 126336
rect 71501 126327 71559 126333
rect 71501 126293 71513 126327
rect 71547 126324 71559 126327
rect 71774 126324 71780 126336
rect 71547 126296 71780 126324
rect 71547 126293 71559 126296
rect 71501 126287 71559 126293
rect 71774 126284 71780 126296
rect 71832 126284 71838 126336
rect 86310 126284 86316 126336
rect 86368 126284 86374 126336
rect 87322 126284 87328 126336
rect 87380 126284 87386 126336
rect 95973 126327 96031 126333
rect 95973 126293 95985 126327
rect 96019 126324 96031 126327
rect 96062 126324 96068 126336
rect 96019 126296 96068 126324
rect 96019 126293 96031 126296
rect 95973 126287 96031 126293
rect 96062 126284 96068 126296
rect 96120 126284 96126 126336
rect 1104 126234 108836 126256
rect 1104 126182 4874 126234
rect 4926 126182 4938 126234
rect 4990 126182 5002 126234
rect 5054 126182 5066 126234
rect 5118 126182 5130 126234
rect 5182 126182 35594 126234
rect 35646 126182 35658 126234
rect 35710 126182 35722 126234
rect 35774 126182 35786 126234
rect 35838 126182 35850 126234
rect 35902 126182 66314 126234
rect 66366 126182 66378 126234
rect 66430 126182 66442 126234
rect 66494 126182 66506 126234
rect 66558 126182 66570 126234
rect 66622 126182 97034 126234
rect 97086 126182 97098 126234
rect 97150 126182 97162 126234
rect 97214 126182 97226 126234
rect 97278 126182 97290 126234
rect 97342 126182 106658 126234
rect 106710 126182 106722 126234
rect 106774 126182 106786 126234
rect 106838 126182 106850 126234
rect 106902 126182 106914 126234
rect 106966 126182 108836 126234
rect 1104 126160 108836 126182
rect 9582 126080 9588 126132
rect 9640 126120 9646 126132
rect 49602 126120 49608 126132
rect 9640 126092 49608 126120
rect 9640 126080 9646 126092
rect 49602 126080 49608 126092
rect 49660 126080 49666 126132
rect 59722 126080 59728 126132
rect 59780 126120 59786 126132
rect 103514 126120 103520 126132
rect 59780 126092 103520 126120
rect 59780 126080 59786 126092
rect 103514 126080 103520 126092
rect 103572 126080 103578 126132
rect 8202 126012 8208 126064
rect 8260 126052 8266 126064
rect 45094 126052 45100 126064
rect 8260 126024 45100 126052
rect 8260 126012 8266 126024
rect 45094 126012 45100 126024
rect 45152 126012 45158 126064
rect 62206 126012 62212 126064
rect 62264 126052 62270 126064
rect 102410 126052 102416 126064
rect 62264 126024 102416 126052
rect 62264 126012 62270 126024
rect 102410 126012 102416 126024
rect 102468 126012 102474 126064
rect 8110 125944 8116 125996
rect 8168 125984 8174 125996
rect 41414 125984 41420 125996
rect 8168 125956 41420 125984
rect 8168 125944 8174 125956
rect 41414 125944 41420 125956
rect 41472 125944 41478 125996
rect 64322 125944 64328 125996
rect 64380 125984 64386 125996
rect 102686 125984 102692 125996
rect 64380 125956 102692 125984
rect 64380 125944 64386 125956
rect 102686 125944 102692 125956
rect 102744 125944 102750 125996
rect 7926 125876 7932 125928
rect 7984 125916 7990 125928
rect 40954 125916 40960 125928
rect 7984 125888 40960 125916
rect 7984 125876 7990 125888
rect 40954 125876 40960 125888
rect 41012 125876 41018 125928
rect 65978 125876 65984 125928
rect 66036 125916 66042 125928
rect 103606 125916 103612 125928
rect 66036 125888 103612 125916
rect 66036 125876 66042 125888
rect 103606 125876 103612 125888
rect 103664 125876 103670 125928
rect 7834 125808 7840 125860
rect 7892 125848 7898 125860
rect 37642 125848 37648 125860
rect 7892 125820 37648 125848
rect 7892 125808 7898 125820
rect 37642 125808 37648 125820
rect 37700 125808 37706 125860
rect 67082 125808 67088 125860
rect 67140 125848 67146 125860
rect 102502 125848 102508 125860
rect 67140 125820 102508 125848
rect 67140 125808 67146 125820
rect 102502 125808 102508 125820
rect 102560 125808 102566 125860
rect 9490 125740 9496 125792
rect 9548 125780 9554 125792
rect 36262 125780 36268 125792
rect 9548 125752 36268 125780
rect 9548 125740 9554 125752
rect 36262 125740 36268 125752
rect 36320 125740 36326 125792
rect 71774 125740 71780 125792
rect 71832 125780 71838 125792
rect 103698 125780 103704 125792
rect 71832 125752 103704 125780
rect 71832 125740 71838 125752
rect 103698 125740 103704 125752
rect 103756 125740 103762 125792
rect 1104 125690 7912 125712
rect 1104 125638 4214 125690
rect 4266 125638 4278 125690
rect 4330 125638 4342 125690
rect 4394 125638 4406 125690
rect 4458 125638 4470 125690
rect 4522 125638 7912 125690
rect 8018 125672 8024 125724
rect 8076 125712 8082 125724
rect 48406 125712 48412 125724
rect 8076 125684 48412 125712
rect 8076 125672 8082 125684
rect 48406 125672 48412 125684
rect 48464 125672 48470 125724
rect 70854 125672 70860 125724
rect 70912 125712 70918 125724
rect 102226 125712 102232 125724
rect 70912 125684 102232 125712
rect 70912 125672 70918 125684
rect 102226 125672 102232 125684
rect 102284 125672 102290 125724
rect 104052 125690 108836 125712
rect 1104 125616 7912 125638
rect 104052 125638 105922 125690
rect 105974 125638 105986 125690
rect 106038 125638 106050 125690
rect 106102 125638 106114 125690
rect 106166 125638 106178 125690
rect 106230 125638 108836 125690
rect 104052 125616 108836 125638
rect 1104 125146 7912 125168
rect 1104 125094 4874 125146
rect 4926 125094 4938 125146
rect 4990 125094 5002 125146
rect 5054 125094 5066 125146
rect 5118 125094 5130 125146
rect 5182 125094 7912 125146
rect 1104 125072 7912 125094
rect 104052 125146 108836 125168
rect 104052 125094 106658 125146
rect 106710 125094 106722 125146
rect 106774 125094 106786 125146
rect 106838 125094 106850 125146
rect 106902 125094 106914 125146
rect 106966 125094 108836 125146
rect 104052 125072 108836 125094
rect 1104 124602 7912 124624
rect 1104 124550 4214 124602
rect 4266 124550 4278 124602
rect 4330 124550 4342 124602
rect 4394 124550 4406 124602
rect 4458 124550 4470 124602
rect 4522 124550 7912 124602
rect 1104 124528 7912 124550
rect 104052 124602 108836 124624
rect 104052 124550 105922 124602
rect 105974 124550 105986 124602
rect 106038 124550 106050 124602
rect 106102 124550 106114 124602
rect 106166 124550 106178 124602
rect 106230 124550 108836 124602
rect 104052 124528 108836 124550
rect 1104 124058 7912 124080
rect 1104 124006 4874 124058
rect 4926 124006 4938 124058
rect 4990 124006 5002 124058
rect 5054 124006 5066 124058
rect 5118 124006 5130 124058
rect 5182 124006 7912 124058
rect 1104 123984 7912 124006
rect 104052 124058 108836 124080
rect 104052 124006 106658 124058
rect 106710 124006 106722 124058
rect 106774 124006 106786 124058
rect 106838 124006 106850 124058
rect 106902 124006 106914 124058
rect 106966 124006 108836 124058
rect 104052 123984 108836 124006
rect 87322 123700 87328 123752
rect 87380 123740 87386 123752
rect 104434 123740 104440 123752
rect 87380 123712 104440 123740
rect 87380 123700 87386 123712
rect 104434 123700 104440 123712
rect 104492 123700 104498 123752
rect 1104 123514 7912 123536
rect 1104 123462 4214 123514
rect 4266 123462 4278 123514
rect 4330 123462 4342 123514
rect 4394 123462 4406 123514
rect 4458 123462 4470 123514
rect 4522 123462 7912 123514
rect 1104 123440 7912 123462
rect 104052 123514 108836 123536
rect 104052 123462 105922 123514
rect 105974 123462 105986 123514
rect 106038 123462 106050 123514
rect 106102 123462 106114 123514
rect 106166 123462 106178 123514
rect 106230 123462 108836 123514
rect 104052 123440 108836 123462
rect 1104 122970 7912 122992
rect 1104 122918 4874 122970
rect 4926 122918 4938 122970
rect 4990 122918 5002 122970
rect 5054 122918 5066 122970
rect 5118 122918 5130 122970
rect 5182 122918 7912 122970
rect 1104 122896 7912 122918
rect 104052 122970 108836 122992
rect 104052 122918 106658 122970
rect 106710 122918 106722 122970
rect 106774 122918 106786 122970
rect 106838 122918 106850 122970
rect 106902 122918 106914 122970
rect 106966 122918 108836 122970
rect 104052 122896 108836 122918
rect 1104 122426 7912 122448
rect 1104 122374 4214 122426
rect 4266 122374 4278 122426
rect 4330 122374 4342 122426
rect 4394 122374 4406 122426
rect 4458 122374 4470 122426
rect 4522 122374 7912 122426
rect 1104 122352 7912 122374
rect 104052 122426 108836 122448
rect 104052 122374 105922 122426
rect 105974 122374 105986 122426
rect 106038 122374 106050 122426
rect 106102 122374 106114 122426
rect 106166 122374 106178 122426
rect 106230 122374 108836 122426
rect 104052 122352 108836 122374
rect 1104 121882 7912 121904
rect 1104 121830 4874 121882
rect 4926 121830 4938 121882
rect 4990 121830 5002 121882
rect 5054 121830 5066 121882
rect 5118 121830 5130 121882
rect 5182 121830 7912 121882
rect 1104 121808 7912 121830
rect 104052 121882 108836 121904
rect 104052 121830 106658 121882
rect 106710 121830 106722 121882
rect 106774 121830 106786 121882
rect 106838 121830 106850 121882
rect 106902 121830 106914 121882
rect 106966 121830 108836 121882
rect 104052 121808 108836 121830
rect 1104 121338 7912 121360
rect 1104 121286 4214 121338
rect 4266 121286 4278 121338
rect 4330 121286 4342 121338
rect 4394 121286 4406 121338
rect 4458 121286 4470 121338
rect 4522 121286 7912 121338
rect 1104 121264 7912 121286
rect 104052 121338 108836 121360
rect 104052 121286 105922 121338
rect 105974 121286 105986 121338
rect 106038 121286 106050 121338
rect 106102 121286 106114 121338
rect 106166 121286 106178 121338
rect 106230 121286 108836 121338
rect 104052 121264 108836 121286
rect 1104 120794 7912 120816
rect 1104 120742 4874 120794
rect 4926 120742 4938 120794
rect 4990 120742 5002 120794
rect 5054 120742 5066 120794
rect 5118 120742 5130 120794
rect 5182 120742 7912 120794
rect 1104 120720 7912 120742
rect 104052 120794 108836 120816
rect 104052 120742 106658 120794
rect 106710 120742 106722 120794
rect 106774 120742 106786 120794
rect 106838 120742 106850 120794
rect 106902 120742 106914 120794
rect 106966 120742 108836 120794
rect 104052 120720 108836 120742
rect 1104 120250 7912 120272
rect 1104 120198 4214 120250
rect 4266 120198 4278 120250
rect 4330 120198 4342 120250
rect 4394 120198 4406 120250
rect 4458 120198 4470 120250
rect 4522 120198 7912 120250
rect 1104 120176 7912 120198
rect 104052 120250 108836 120272
rect 104052 120198 105922 120250
rect 105974 120198 105986 120250
rect 106038 120198 106050 120250
rect 106102 120198 106114 120250
rect 106166 120198 106178 120250
rect 106230 120198 108836 120250
rect 104052 120176 108836 120198
rect 104342 119892 104348 119944
rect 104400 119892 104406 119944
rect 1104 119706 7912 119728
rect 1104 119654 4874 119706
rect 4926 119654 4938 119706
rect 4990 119654 5002 119706
rect 5054 119654 5066 119706
rect 5118 119654 5130 119706
rect 5182 119654 7912 119706
rect 1104 119632 7912 119654
rect 104052 119706 108836 119728
rect 104052 119654 106658 119706
rect 106710 119654 106722 119706
rect 106774 119654 106786 119706
rect 106838 119654 106850 119706
rect 106902 119654 106914 119706
rect 106966 119654 108836 119706
rect 104052 119632 108836 119654
rect 1104 119162 7912 119184
rect 1104 119110 4214 119162
rect 4266 119110 4278 119162
rect 4330 119110 4342 119162
rect 4394 119110 4406 119162
rect 4458 119110 4470 119162
rect 4522 119110 7912 119162
rect 1104 119088 7912 119110
rect 104052 119162 108836 119184
rect 104052 119110 105922 119162
rect 105974 119110 105986 119162
rect 106038 119110 106050 119162
rect 106102 119110 106114 119162
rect 106166 119110 106178 119162
rect 106230 119110 108836 119162
rect 104052 119088 108836 119110
rect 1104 118618 7912 118640
rect 1104 118566 4874 118618
rect 4926 118566 4938 118618
rect 4990 118566 5002 118618
rect 5054 118566 5066 118618
rect 5118 118566 5130 118618
rect 5182 118566 7912 118618
rect 1104 118544 7912 118566
rect 104052 118618 108836 118640
rect 104052 118566 106658 118618
rect 106710 118566 106722 118618
rect 106774 118566 106786 118618
rect 106838 118566 106850 118618
rect 106902 118566 106914 118618
rect 106966 118566 108836 118618
rect 104052 118544 108836 118566
rect 1104 118074 7912 118096
rect 1104 118022 4214 118074
rect 4266 118022 4278 118074
rect 4330 118022 4342 118074
rect 4394 118022 4406 118074
rect 4458 118022 4470 118074
rect 4522 118022 7912 118074
rect 1104 118000 7912 118022
rect 104052 118074 108836 118096
rect 104052 118022 105922 118074
rect 105974 118022 105986 118074
rect 106038 118022 106050 118074
rect 106102 118022 106114 118074
rect 106166 118022 106178 118074
rect 106230 118022 108836 118074
rect 104052 118000 108836 118022
rect 1104 117530 7912 117552
rect 1104 117478 4874 117530
rect 4926 117478 4938 117530
rect 4990 117478 5002 117530
rect 5054 117478 5066 117530
rect 5118 117478 5130 117530
rect 5182 117478 7912 117530
rect 1104 117456 7912 117478
rect 104052 117530 108836 117552
rect 104052 117478 106658 117530
rect 106710 117478 106722 117530
rect 106774 117478 106786 117530
rect 106838 117478 106850 117530
rect 106902 117478 106914 117530
rect 106966 117478 108836 117530
rect 104052 117456 108836 117478
rect 1104 116986 7912 117008
rect 1104 116934 4214 116986
rect 4266 116934 4278 116986
rect 4330 116934 4342 116986
rect 4394 116934 4406 116986
rect 4458 116934 4470 116986
rect 4522 116934 7912 116986
rect 1104 116912 7912 116934
rect 104052 116986 108836 117008
rect 104052 116934 105922 116986
rect 105974 116934 105986 116986
rect 106038 116934 106050 116986
rect 106102 116934 106114 116986
rect 106166 116934 106178 116986
rect 106230 116934 108836 116986
rect 104052 116912 108836 116934
rect 1104 116442 7912 116464
rect 1104 116390 4874 116442
rect 4926 116390 4938 116442
rect 4990 116390 5002 116442
rect 5054 116390 5066 116442
rect 5118 116390 5130 116442
rect 5182 116390 7912 116442
rect 1104 116368 7912 116390
rect 104052 116442 108836 116464
rect 104052 116390 106658 116442
rect 106710 116390 106722 116442
rect 106774 116390 106786 116442
rect 106838 116390 106850 116442
rect 106902 116390 106914 116442
rect 106966 116390 108836 116442
rect 104052 116368 108836 116390
rect 1104 115898 7912 115920
rect 1104 115846 4214 115898
rect 4266 115846 4278 115898
rect 4330 115846 4342 115898
rect 4394 115846 4406 115898
rect 4458 115846 4470 115898
rect 4522 115846 7912 115898
rect 1104 115824 7912 115846
rect 104052 115898 108836 115920
rect 104052 115846 105922 115898
rect 105974 115846 105986 115898
rect 106038 115846 106050 115898
rect 106102 115846 106114 115898
rect 106166 115846 106178 115898
rect 106230 115846 108836 115898
rect 104052 115824 108836 115846
rect 1104 115354 7912 115376
rect 1104 115302 4874 115354
rect 4926 115302 4938 115354
rect 4990 115302 5002 115354
rect 5054 115302 5066 115354
rect 5118 115302 5130 115354
rect 5182 115302 7912 115354
rect 1104 115280 7912 115302
rect 104052 115354 108836 115376
rect 104052 115302 106658 115354
rect 106710 115302 106722 115354
rect 106774 115302 106786 115354
rect 106838 115302 106850 115354
rect 106902 115302 106914 115354
rect 106966 115302 108836 115354
rect 104052 115280 108836 115302
rect 1104 114810 7912 114832
rect 1104 114758 4214 114810
rect 4266 114758 4278 114810
rect 4330 114758 4342 114810
rect 4394 114758 4406 114810
rect 4458 114758 4470 114810
rect 4522 114758 7912 114810
rect 1104 114736 7912 114758
rect 104052 114810 108836 114832
rect 104052 114758 105922 114810
rect 105974 114758 105986 114810
rect 106038 114758 106050 114810
rect 106102 114758 106114 114810
rect 106166 114758 106178 114810
rect 106230 114758 108836 114810
rect 104052 114736 108836 114758
rect 1104 114266 7912 114288
rect 1104 114214 4874 114266
rect 4926 114214 4938 114266
rect 4990 114214 5002 114266
rect 5054 114214 5066 114266
rect 5118 114214 5130 114266
rect 5182 114214 7912 114266
rect 1104 114192 7912 114214
rect 104052 114266 108836 114288
rect 104052 114214 106658 114266
rect 106710 114214 106722 114266
rect 106774 114214 106786 114266
rect 106838 114214 106850 114266
rect 106902 114214 106914 114266
rect 106966 114214 108836 114266
rect 104052 114192 108836 114214
rect 1104 113722 7912 113744
rect 1104 113670 4214 113722
rect 4266 113670 4278 113722
rect 4330 113670 4342 113722
rect 4394 113670 4406 113722
rect 4458 113670 4470 113722
rect 4522 113670 7912 113722
rect 1104 113648 7912 113670
rect 104052 113722 108836 113744
rect 104052 113670 105922 113722
rect 105974 113670 105986 113722
rect 106038 113670 106050 113722
rect 106102 113670 106114 113722
rect 106166 113670 106178 113722
rect 106230 113670 108836 113722
rect 104052 113648 108836 113670
rect 1104 113178 7912 113200
rect 1104 113126 4874 113178
rect 4926 113126 4938 113178
rect 4990 113126 5002 113178
rect 5054 113126 5066 113178
rect 5118 113126 5130 113178
rect 5182 113126 7912 113178
rect 1104 113104 7912 113126
rect 104052 113178 108836 113200
rect 104052 113126 106658 113178
rect 106710 113126 106722 113178
rect 106774 113126 106786 113178
rect 106838 113126 106850 113178
rect 106902 113126 106914 113178
rect 106966 113126 108836 113178
rect 104052 113104 108836 113126
rect 1104 112634 7912 112656
rect 1104 112582 4214 112634
rect 4266 112582 4278 112634
rect 4330 112582 4342 112634
rect 4394 112582 4406 112634
rect 4458 112582 4470 112634
rect 4522 112582 7912 112634
rect 1104 112560 7912 112582
rect 104052 112634 108836 112656
rect 104052 112582 105922 112634
rect 105974 112582 105986 112634
rect 106038 112582 106050 112634
rect 106102 112582 106114 112634
rect 106166 112582 106178 112634
rect 106230 112582 108836 112634
rect 104052 112560 108836 112582
rect 1104 112090 7912 112112
rect 1104 112038 4874 112090
rect 4926 112038 4938 112090
rect 4990 112038 5002 112090
rect 5054 112038 5066 112090
rect 5118 112038 5130 112090
rect 5182 112038 7912 112090
rect 1104 112016 7912 112038
rect 104052 112090 108836 112112
rect 104052 112038 106658 112090
rect 106710 112038 106722 112090
rect 106774 112038 106786 112090
rect 106838 112038 106850 112090
rect 106902 112038 106914 112090
rect 106966 112038 108836 112090
rect 104052 112016 108836 112038
rect 1104 111546 7912 111568
rect 1104 111494 4214 111546
rect 4266 111494 4278 111546
rect 4330 111494 4342 111546
rect 4394 111494 4406 111546
rect 4458 111494 4470 111546
rect 4522 111494 7912 111546
rect 1104 111472 7912 111494
rect 104052 111546 108836 111568
rect 104052 111494 105922 111546
rect 105974 111494 105986 111546
rect 106038 111494 106050 111546
rect 106102 111494 106114 111546
rect 106166 111494 106178 111546
rect 106230 111494 108836 111546
rect 104052 111472 108836 111494
rect 1104 111002 7912 111024
rect 1104 110950 4874 111002
rect 4926 110950 4938 111002
rect 4990 110950 5002 111002
rect 5054 110950 5066 111002
rect 5118 110950 5130 111002
rect 5182 110950 7912 111002
rect 1104 110928 7912 110950
rect 104052 111002 108836 111024
rect 104052 110950 106658 111002
rect 106710 110950 106722 111002
rect 106774 110950 106786 111002
rect 106838 110950 106850 111002
rect 106902 110950 106914 111002
rect 106966 110950 108836 111002
rect 104052 110928 108836 110950
rect 1104 110458 7912 110480
rect 1104 110406 4214 110458
rect 4266 110406 4278 110458
rect 4330 110406 4342 110458
rect 4394 110406 4406 110458
rect 4458 110406 4470 110458
rect 4522 110406 7912 110458
rect 1104 110384 7912 110406
rect 104052 110458 108836 110480
rect 104052 110406 105922 110458
rect 105974 110406 105986 110458
rect 106038 110406 106050 110458
rect 106102 110406 106114 110458
rect 106166 110406 106178 110458
rect 106230 110406 108836 110458
rect 104052 110384 108836 110406
rect 1104 109914 7912 109936
rect 1104 109862 4874 109914
rect 4926 109862 4938 109914
rect 4990 109862 5002 109914
rect 5054 109862 5066 109914
rect 5118 109862 5130 109914
rect 5182 109862 7912 109914
rect 1104 109840 7912 109862
rect 104052 109914 108836 109936
rect 104052 109862 106658 109914
rect 106710 109862 106722 109914
rect 106774 109862 106786 109914
rect 106838 109862 106850 109914
rect 106902 109862 106914 109914
rect 106966 109862 108836 109914
rect 104052 109840 108836 109862
rect 1104 109370 7912 109392
rect 1104 109318 4214 109370
rect 4266 109318 4278 109370
rect 4330 109318 4342 109370
rect 4394 109318 4406 109370
rect 4458 109318 4470 109370
rect 4522 109318 7912 109370
rect 1104 109296 7912 109318
rect 104052 109370 108836 109392
rect 104052 109318 105922 109370
rect 105974 109318 105986 109370
rect 106038 109318 106050 109370
rect 106102 109318 106114 109370
rect 106166 109318 106178 109370
rect 106230 109318 108836 109370
rect 104052 109296 108836 109318
rect 1104 108826 7912 108848
rect 1104 108774 4874 108826
rect 4926 108774 4938 108826
rect 4990 108774 5002 108826
rect 5054 108774 5066 108826
rect 5118 108774 5130 108826
rect 5182 108774 7912 108826
rect 1104 108752 7912 108774
rect 104052 108826 108836 108848
rect 104052 108774 106658 108826
rect 106710 108774 106722 108826
rect 106774 108774 106786 108826
rect 106838 108774 106850 108826
rect 106902 108774 106914 108826
rect 106966 108774 108836 108826
rect 104052 108752 108836 108774
rect 1104 108282 7912 108304
rect 1104 108230 4214 108282
rect 4266 108230 4278 108282
rect 4330 108230 4342 108282
rect 4394 108230 4406 108282
rect 4458 108230 4470 108282
rect 4522 108230 7912 108282
rect 1104 108208 7912 108230
rect 104052 108282 108836 108304
rect 104052 108230 105922 108282
rect 105974 108230 105986 108282
rect 106038 108230 106050 108282
rect 106102 108230 106114 108282
rect 106166 108230 106178 108282
rect 106230 108230 108836 108282
rect 104052 108208 108836 108230
rect 1104 107738 7912 107760
rect 1104 107686 4874 107738
rect 4926 107686 4938 107738
rect 4990 107686 5002 107738
rect 5054 107686 5066 107738
rect 5118 107686 5130 107738
rect 5182 107686 7912 107738
rect 1104 107664 7912 107686
rect 104052 107738 108836 107760
rect 104052 107686 106658 107738
rect 106710 107686 106722 107738
rect 106774 107686 106786 107738
rect 106838 107686 106850 107738
rect 106902 107686 106914 107738
rect 106966 107686 108836 107738
rect 104052 107664 108836 107686
rect 1104 107194 7912 107216
rect 1104 107142 4214 107194
rect 4266 107142 4278 107194
rect 4330 107142 4342 107194
rect 4394 107142 4406 107194
rect 4458 107142 4470 107194
rect 4522 107142 7912 107194
rect 1104 107120 7912 107142
rect 104052 107194 108836 107216
rect 104052 107142 105922 107194
rect 105974 107142 105986 107194
rect 106038 107142 106050 107194
rect 106102 107142 106114 107194
rect 106166 107142 106178 107194
rect 106230 107142 108836 107194
rect 104052 107120 108836 107142
rect 1104 106650 7912 106672
rect 1104 106598 4874 106650
rect 4926 106598 4938 106650
rect 4990 106598 5002 106650
rect 5054 106598 5066 106650
rect 5118 106598 5130 106650
rect 5182 106598 7912 106650
rect 1104 106576 7912 106598
rect 104052 106650 108836 106672
rect 104052 106598 106658 106650
rect 106710 106598 106722 106650
rect 106774 106598 106786 106650
rect 106838 106598 106850 106650
rect 106902 106598 106914 106650
rect 106966 106598 108836 106650
rect 104052 106576 108836 106598
rect 1104 106106 7912 106128
rect 1104 106054 4214 106106
rect 4266 106054 4278 106106
rect 4330 106054 4342 106106
rect 4394 106054 4406 106106
rect 4458 106054 4470 106106
rect 4522 106054 7912 106106
rect 1104 106032 7912 106054
rect 104052 106106 108836 106128
rect 104052 106054 105922 106106
rect 105974 106054 105986 106106
rect 106038 106054 106050 106106
rect 106102 106054 106114 106106
rect 106166 106054 106178 106106
rect 106230 106054 108836 106106
rect 104052 106032 108836 106054
rect 1104 105562 7912 105584
rect 1104 105510 4874 105562
rect 4926 105510 4938 105562
rect 4990 105510 5002 105562
rect 5054 105510 5066 105562
rect 5118 105510 5130 105562
rect 5182 105510 7912 105562
rect 1104 105488 7912 105510
rect 104052 105562 108836 105584
rect 104052 105510 106658 105562
rect 106710 105510 106722 105562
rect 106774 105510 106786 105562
rect 106838 105510 106850 105562
rect 106902 105510 106914 105562
rect 106966 105510 108836 105562
rect 104052 105488 108836 105510
rect 1104 105018 7912 105040
rect 1104 104966 4214 105018
rect 4266 104966 4278 105018
rect 4330 104966 4342 105018
rect 4394 104966 4406 105018
rect 4458 104966 4470 105018
rect 4522 104966 7912 105018
rect 1104 104944 7912 104966
rect 104052 105018 108836 105040
rect 104052 104966 105922 105018
rect 105974 104966 105986 105018
rect 106038 104966 106050 105018
rect 106102 104966 106114 105018
rect 106166 104966 106178 105018
rect 106230 104966 108836 105018
rect 104052 104944 108836 104966
rect 1104 104474 7912 104496
rect 1104 104422 4874 104474
rect 4926 104422 4938 104474
rect 4990 104422 5002 104474
rect 5054 104422 5066 104474
rect 5118 104422 5130 104474
rect 5182 104422 7912 104474
rect 1104 104400 7912 104422
rect 104052 104474 108836 104496
rect 104052 104422 106658 104474
rect 106710 104422 106722 104474
rect 106774 104422 106786 104474
rect 106838 104422 106850 104474
rect 106902 104422 106914 104474
rect 106966 104422 108836 104474
rect 104052 104400 108836 104422
rect 1104 103930 7912 103952
rect 1104 103878 4214 103930
rect 4266 103878 4278 103930
rect 4330 103878 4342 103930
rect 4394 103878 4406 103930
rect 4458 103878 4470 103930
rect 4522 103878 7912 103930
rect 1104 103856 7912 103878
rect 104052 103930 108836 103952
rect 104052 103878 105922 103930
rect 105974 103878 105986 103930
rect 106038 103878 106050 103930
rect 106102 103878 106114 103930
rect 106166 103878 106178 103930
rect 106230 103878 108836 103930
rect 104052 103856 108836 103878
rect 1104 103386 7912 103408
rect 1104 103334 4874 103386
rect 4926 103334 4938 103386
rect 4990 103334 5002 103386
rect 5054 103334 5066 103386
rect 5118 103334 5130 103386
rect 5182 103334 7912 103386
rect 1104 103312 7912 103334
rect 104052 103386 108836 103408
rect 104052 103334 106658 103386
rect 106710 103334 106722 103386
rect 106774 103334 106786 103386
rect 106838 103334 106850 103386
rect 106902 103334 106914 103386
rect 106966 103334 108836 103386
rect 104052 103312 108836 103334
rect 1104 102842 7912 102864
rect 1104 102790 4214 102842
rect 4266 102790 4278 102842
rect 4330 102790 4342 102842
rect 4394 102790 4406 102842
rect 4458 102790 4470 102842
rect 4522 102790 7912 102842
rect 1104 102768 7912 102790
rect 104052 102842 108836 102864
rect 104052 102790 105922 102842
rect 105974 102790 105986 102842
rect 106038 102790 106050 102842
rect 106102 102790 106114 102842
rect 106166 102790 106178 102842
rect 106230 102790 108836 102842
rect 104052 102768 108836 102790
rect 1104 102298 7912 102320
rect 1104 102246 4874 102298
rect 4926 102246 4938 102298
rect 4990 102246 5002 102298
rect 5054 102246 5066 102298
rect 5118 102246 5130 102298
rect 5182 102246 7912 102298
rect 1104 102224 7912 102246
rect 104052 102298 108836 102320
rect 104052 102246 106658 102298
rect 106710 102246 106722 102298
rect 106774 102246 106786 102298
rect 106838 102246 106850 102298
rect 106902 102246 106914 102298
rect 106966 102246 108836 102298
rect 104052 102224 108836 102246
rect 1104 101754 7912 101776
rect 1104 101702 4214 101754
rect 4266 101702 4278 101754
rect 4330 101702 4342 101754
rect 4394 101702 4406 101754
rect 4458 101702 4470 101754
rect 4522 101702 7912 101754
rect 1104 101680 7912 101702
rect 104052 101754 108836 101776
rect 104052 101702 105922 101754
rect 105974 101702 105986 101754
rect 106038 101702 106050 101754
rect 106102 101702 106114 101754
rect 106166 101702 106178 101754
rect 106230 101702 108836 101754
rect 104052 101680 108836 101702
rect 1581 101575 1639 101581
rect 1581 101541 1593 101575
rect 1627 101572 1639 101575
rect 8386 101572 8392 101584
rect 1627 101544 8392 101572
rect 1627 101541 1639 101544
rect 1581 101535 1639 101541
rect 8386 101532 8392 101544
rect 8444 101532 8450 101584
rect 1210 101396 1216 101448
rect 1268 101436 1274 101448
rect 1397 101439 1455 101445
rect 1397 101436 1409 101439
rect 1268 101408 1409 101436
rect 1268 101396 1274 101408
rect 1397 101405 1409 101408
rect 1443 101436 1455 101439
rect 1673 101439 1731 101445
rect 1673 101436 1685 101439
rect 1443 101408 1685 101436
rect 1443 101405 1455 101408
rect 1397 101399 1455 101405
rect 1673 101405 1685 101408
rect 1719 101405 1731 101439
rect 1673 101399 1731 101405
rect 1104 101210 7912 101232
rect 1104 101158 4874 101210
rect 4926 101158 4938 101210
rect 4990 101158 5002 101210
rect 5054 101158 5066 101210
rect 5118 101158 5130 101210
rect 5182 101158 7912 101210
rect 1104 101136 7912 101158
rect 104052 101210 108836 101232
rect 104052 101158 106658 101210
rect 106710 101158 106722 101210
rect 106774 101158 106786 101210
rect 106838 101158 106850 101210
rect 106902 101158 106914 101210
rect 106966 101158 108836 101210
rect 104052 101136 108836 101158
rect 1104 100666 7912 100688
rect 1104 100614 4214 100666
rect 4266 100614 4278 100666
rect 4330 100614 4342 100666
rect 4394 100614 4406 100666
rect 4458 100614 4470 100666
rect 4522 100614 7912 100666
rect 1104 100592 7912 100614
rect 104052 100666 108836 100688
rect 104052 100614 105922 100666
rect 105974 100614 105986 100666
rect 106038 100614 106050 100666
rect 106102 100614 106114 100666
rect 106166 100614 106178 100666
rect 106230 100614 108836 100666
rect 104052 100592 108836 100614
rect 1104 100122 7912 100144
rect 1104 100070 4874 100122
rect 4926 100070 4938 100122
rect 4990 100070 5002 100122
rect 5054 100070 5066 100122
rect 5118 100070 5130 100122
rect 5182 100070 7912 100122
rect 1104 100048 7912 100070
rect 104052 100122 108836 100144
rect 104052 100070 106658 100122
rect 106710 100070 106722 100122
rect 106774 100070 106786 100122
rect 106838 100070 106850 100122
rect 106902 100070 106914 100122
rect 106966 100070 108836 100122
rect 104052 100048 108836 100070
rect 1394 99832 1400 99884
rect 1452 99872 1458 99884
rect 1673 99875 1731 99881
rect 1673 99872 1685 99875
rect 1452 99844 1685 99872
rect 1452 99832 1458 99844
rect 1673 99841 1685 99844
rect 1719 99841 1731 99875
rect 1673 99835 1731 99841
rect 1581 99739 1639 99745
rect 1581 99705 1593 99739
rect 1627 99736 1639 99739
rect 8386 99736 8392 99748
rect 1627 99708 8392 99736
rect 1627 99705 1639 99708
rect 1581 99699 1639 99705
rect 8386 99696 8392 99708
rect 8444 99696 8450 99748
rect 1104 99578 7912 99600
rect 1104 99526 4214 99578
rect 4266 99526 4278 99578
rect 4330 99526 4342 99578
rect 4394 99526 4406 99578
rect 4458 99526 4470 99578
rect 4522 99526 7912 99578
rect 1104 99504 7912 99526
rect 104052 99578 108836 99600
rect 104052 99526 105922 99578
rect 105974 99526 105986 99578
rect 106038 99526 106050 99578
rect 106102 99526 106114 99578
rect 106166 99526 106178 99578
rect 106230 99526 108836 99578
rect 104052 99504 108836 99526
rect 1104 99034 7912 99056
rect 1104 98982 4874 99034
rect 4926 98982 4938 99034
rect 4990 98982 5002 99034
rect 5054 98982 5066 99034
rect 5118 98982 5130 99034
rect 5182 98982 7912 99034
rect 1104 98960 7912 98982
rect 104052 99034 108836 99056
rect 104052 98982 106658 99034
rect 106710 98982 106722 99034
rect 106774 98982 106786 99034
rect 106838 98982 106850 99034
rect 106902 98982 106914 99034
rect 106966 98982 108836 99034
rect 104052 98960 108836 98982
rect 1302 98744 1308 98796
rect 1360 98784 1366 98796
rect 1397 98787 1455 98793
rect 1397 98784 1409 98787
rect 1360 98756 1409 98784
rect 1360 98744 1366 98756
rect 1397 98753 1409 98756
rect 1443 98784 1455 98787
rect 1673 98787 1731 98793
rect 1673 98784 1685 98787
rect 1443 98756 1685 98784
rect 1443 98753 1455 98756
rect 1397 98747 1455 98753
rect 1673 98753 1685 98756
rect 1719 98753 1731 98787
rect 1673 98747 1731 98753
rect 1581 98651 1639 98657
rect 1581 98617 1593 98651
rect 1627 98648 1639 98651
rect 8386 98648 8392 98660
rect 1627 98620 8392 98648
rect 1627 98617 1639 98620
rect 1581 98611 1639 98617
rect 8386 98608 8392 98620
rect 8444 98608 8450 98660
rect 1104 98490 7912 98512
rect 1104 98438 4214 98490
rect 4266 98438 4278 98490
rect 4330 98438 4342 98490
rect 4394 98438 4406 98490
rect 4458 98438 4470 98490
rect 4522 98438 7912 98490
rect 1104 98416 7912 98438
rect 104052 98490 108836 98512
rect 104052 98438 105922 98490
rect 105974 98438 105986 98490
rect 106038 98438 106050 98490
rect 106102 98438 106114 98490
rect 106166 98438 106178 98490
rect 106230 98438 108836 98490
rect 104052 98416 108836 98438
rect 1104 97946 7912 97968
rect 1104 97894 4874 97946
rect 4926 97894 4938 97946
rect 4990 97894 5002 97946
rect 5054 97894 5066 97946
rect 5118 97894 5130 97946
rect 5182 97894 7912 97946
rect 1104 97872 7912 97894
rect 104052 97946 108836 97968
rect 104052 97894 106658 97946
rect 106710 97894 106722 97946
rect 106774 97894 106786 97946
rect 106838 97894 106850 97946
rect 106902 97894 106914 97946
rect 106966 97894 108836 97946
rect 104052 97872 108836 97894
rect 1104 97402 7912 97424
rect 1104 97350 4214 97402
rect 4266 97350 4278 97402
rect 4330 97350 4342 97402
rect 4394 97350 4406 97402
rect 4458 97350 4470 97402
rect 4522 97350 7912 97402
rect 1104 97328 7912 97350
rect 104052 97402 108836 97424
rect 104052 97350 105922 97402
rect 105974 97350 105986 97402
rect 106038 97350 106050 97402
rect 106102 97350 106114 97402
rect 106166 97350 106178 97402
rect 106230 97350 108836 97402
rect 104052 97328 108836 97350
rect 1581 97223 1639 97229
rect 1581 97189 1593 97223
rect 1627 97220 1639 97223
rect 8386 97220 8392 97232
rect 1627 97192 8392 97220
rect 1627 97189 1639 97192
rect 1581 97183 1639 97189
rect 8386 97180 8392 97192
rect 8444 97180 8450 97232
rect 1302 97044 1308 97096
rect 1360 97084 1366 97096
rect 1397 97087 1455 97093
rect 1397 97084 1409 97087
rect 1360 97056 1409 97084
rect 1360 97044 1366 97056
rect 1397 97053 1409 97056
rect 1443 97084 1455 97087
rect 1673 97087 1731 97093
rect 1673 97084 1685 97087
rect 1443 97056 1685 97084
rect 1443 97053 1455 97056
rect 1397 97047 1455 97053
rect 1673 97053 1685 97056
rect 1719 97053 1731 97087
rect 1673 97047 1731 97053
rect 1104 96858 7912 96880
rect 1104 96806 4874 96858
rect 4926 96806 4938 96858
rect 4990 96806 5002 96858
rect 5054 96806 5066 96858
rect 5118 96806 5130 96858
rect 5182 96806 7912 96858
rect 1104 96784 7912 96806
rect 104052 96858 108836 96880
rect 104052 96806 106658 96858
rect 106710 96806 106722 96858
rect 106774 96806 106786 96858
rect 106838 96806 106850 96858
rect 106902 96806 106914 96858
rect 106966 96806 108836 96858
rect 104052 96784 108836 96806
rect 1104 96314 7912 96336
rect 1104 96262 4214 96314
rect 4266 96262 4278 96314
rect 4330 96262 4342 96314
rect 4394 96262 4406 96314
rect 4458 96262 4470 96314
rect 4522 96262 7912 96314
rect 1104 96240 7912 96262
rect 104052 96314 108836 96336
rect 104052 96262 105922 96314
rect 105974 96262 105986 96314
rect 106038 96262 106050 96314
rect 106102 96262 106114 96314
rect 106166 96262 106178 96314
rect 106230 96262 108836 96314
rect 104052 96240 108836 96262
rect 1581 96135 1639 96141
rect 1581 96101 1593 96135
rect 1627 96132 1639 96135
rect 8386 96132 8392 96144
rect 1627 96104 8392 96132
rect 1627 96101 1639 96104
rect 1581 96095 1639 96101
rect 8386 96092 8392 96104
rect 8444 96092 8450 96144
rect 1210 95956 1216 96008
rect 1268 95996 1274 96008
rect 1397 95999 1455 96005
rect 1397 95996 1409 95999
rect 1268 95968 1409 95996
rect 1268 95956 1274 95968
rect 1397 95965 1409 95968
rect 1443 95996 1455 95999
rect 1673 95999 1731 96005
rect 1673 95996 1685 95999
rect 1443 95968 1685 95996
rect 1443 95965 1455 95968
rect 1397 95959 1455 95965
rect 1673 95965 1685 95968
rect 1719 95965 1731 95999
rect 1673 95959 1731 95965
rect 1104 95770 7912 95792
rect 1104 95718 4874 95770
rect 4926 95718 4938 95770
rect 4990 95718 5002 95770
rect 5054 95718 5066 95770
rect 5118 95718 5130 95770
rect 5182 95718 7912 95770
rect 1104 95696 7912 95718
rect 104052 95770 108836 95792
rect 104052 95718 106658 95770
rect 106710 95718 106722 95770
rect 106774 95718 106786 95770
rect 106838 95718 106850 95770
rect 106902 95718 106914 95770
rect 106966 95718 108836 95770
rect 104052 95696 108836 95718
rect 1104 95226 7912 95248
rect 1104 95174 4214 95226
rect 4266 95174 4278 95226
rect 4330 95174 4342 95226
rect 4394 95174 4406 95226
rect 4458 95174 4470 95226
rect 4522 95174 7912 95226
rect 1104 95152 7912 95174
rect 104052 95226 108836 95248
rect 104052 95174 105922 95226
rect 105974 95174 105986 95226
rect 106038 95174 106050 95226
rect 106102 95174 106114 95226
rect 106166 95174 106178 95226
rect 106230 95174 108836 95226
rect 104052 95152 108836 95174
rect 1104 94682 7912 94704
rect 1104 94630 4874 94682
rect 4926 94630 4938 94682
rect 4990 94630 5002 94682
rect 5054 94630 5066 94682
rect 5118 94630 5130 94682
rect 5182 94630 7912 94682
rect 1104 94608 7912 94630
rect 104052 94682 108836 94704
rect 104052 94630 106658 94682
rect 106710 94630 106722 94682
rect 106774 94630 106786 94682
rect 106838 94630 106850 94682
rect 106902 94630 106914 94682
rect 106966 94630 108836 94682
rect 104052 94608 108836 94630
rect 1302 94392 1308 94444
rect 1360 94432 1366 94444
rect 1397 94435 1455 94441
rect 1397 94432 1409 94435
rect 1360 94404 1409 94432
rect 1360 94392 1366 94404
rect 1397 94401 1409 94404
rect 1443 94432 1455 94435
rect 1673 94435 1731 94441
rect 1673 94432 1685 94435
rect 1443 94404 1685 94432
rect 1443 94401 1455 94404
rect 1397 94395 1455 94401
rect 1673 94401 1685 94404
rect 1719 94401 1731 94435
rect 1673 94395 1731 94401
rect 1581 94299 1639 94305
rect 1581 94265 1593 94299
rect 1627 94296 1639 94299
rect 8386 94296 8392 94308
rect 1627 94268 8392 94296
rect 1627 94265 1639 94268
rect 1581 94259 1639 94265
rect 8386 94256 8392 94268
rect 8444 94256 8450 94308
rect 1104 94138 7912 94160
rect 1104 94086 4214 94138
rect 4266 94086 4278 94138
rect 4330 94086 4342 94138
rect 4394 94086 4406 94138
rect 4458 94086 4470 94138
rect 4522 94086 7912 94138
rect 1104 94064 7912 94086
rect 104052 94138 108836 94160
rect 104052 94086 105922 94138
rect 105974 94086 105986 94138
rect 106038 94086 106050 94138
rect 106102 94086 106114 94138
rect 106166 94086 106178 94138
rect 106230 94086 108836 94138
rect 104052 94064 108836 94086
rect 1104 93594 7912 93616
rect 1104 93542 4874 93594
rect 4926 93542 4938 93594
rect 4990 93542 5002 93594
rect 5054 93542 5066 93594
rect 5118 93542 5130 93594
rect 5182 93542 7912 93594
rect 1104 93520 7912 93542
rect 104052 93594 108836 93616
rect 104052 93542 106658 93594
rect 106710 93542 106722 93594
rect 106774 93542 106786 93594
rect 106838 93542 106850 93594
rect 106902 93542 106914 93594
rect 106966 93542 108836 93594
rect 104052 93520 108836 93542
rect 1104 93050 7912 93072
rect 1104 92998 4214 93050
rect 4266 92998 4278 93050
rect 4330 92998 4342 93050
rect 4394 92998 4406 93050
rect 4458 92998 4470 93050
rect 4522 92998 7912 93050
rect 1104 92976 7912 92998
rect 104052 93050 108836 93072
rect 104052 92998 105922 93050
rect 105974 92998 105986 93050
rect 106038 92998 106050 93050
rect 106102 92998 106114 93050
rect 106166 92998 106178 93050
rect 106230 92998 108836 93050
rect 104052 92976 108836 92998
rect 1104 92506 7912 92528
rect 1104 92454 4874 92506
rect 4926 92454 4938 92506
rect 4990 92454 5002 92506
rect 5054 92454 5066 92506
rect 5118 92454 5130 92506
rect 5182 92454 7912 92506
rect 1104 92432 7912 92454
rect 104052 92506 108836 92528
rect 104052 92454 106658 92506
rect 106710 92454 106722 92506
rect 106774 92454 106786 92506
rect 106838 92454 106850 92506
rect 106902 92454 106914 92506
rect 106966 92454 108836 92506
rect 104052 92432 108836 92454
rect 1104 91962 7912 91984
rect 1104 91910 4214 91962
rect 4266 91910 4278 91962
rect 4330 91910 4342 91962
rect 4394 91910 4406 91962
rect 4458 91910 4470 91962
rect 4522 91910 7912 91962
rect 1104 91888 7912 91910
rect 104052 91962 108836 91984
rect 104052 91910 105922 91962
rect 105974 91910 105986 91962
rect 106038 91910 106050 91962
rect 106102 91910 106114 91962
rect 106166 91910 106178 91962
rect 106230 91910 108836 91962
rect 104052 91888 108836 91910
rect 1104 91418 7912 91440
rect 1104 91366 4874 91418
rect 4926 91366 4938 91418
rect 4990 91366 5002 91418
rect 5054 91366 5066 91418
rect 5118 91366 5130 91418
rect 5182 91366 7912 91418
rect 1104 91344 7912 91366
rect 104052 91418 108836 91440
rect 104052 91366 106658 91418
rect 106710 91366 106722 91418
rect 106774 91366 106786 91418
rect 106838 91366 106850 91418
rect 106902 91366 106914 91418
rect 106966 91366 108836 91418
rect 104052 91344 108836 91366
rect 1104 90874 7912 90896
rect 1104 90822 4214 90874
rect 4266 90822 4278 90874
rect 4330 90822 4342 90874
rect 4394 90822 4406 90874
rect 4458 90822 4470 90874
rect 4522 90822 7912 90874
rect 1104 90800 7912 90822
rect 104052 90874 108836 90896
rect 104052 90822 105922 90874
rect 105974 90822 105986 90874
rect 106038 90822 106050 90874
rect 106102 90822 106114 90874
rect 106166 90822 106178 90874
rect 106230 90822 108836 90874
rect 104052 90800 108836 90822
rect 1104 90330 7912 90352
rect 1104 90278 4874 90330
rect 4926 90278 4938 90330
rect 4990 90278 5002 90330
rect 5054 90278 5066 90330
rect 5118 90278 5130 90330
rect 5182 90278 7912 90330
rect 1104 90256 7912 90278
rect 104052 90330 108836 90352
rect 104052 90278 106658 90330
rect 106710 90278 106722 90330
rect 106774 90278 106786 90330
rect 106838 90278 106850 90330
rect 106902 90278 106914 90330
rect 106966 90278 108836 90330
rect 104052 90256 108836 90278
rect 1104 89786 7912 89808
rect 1104 89734 4214 89786
rect 4266 89734 4278 89786
rect 4330 89734 4342 89786
rect 4394 89734 4406 89786
rect 4458 89734 4470 89786
rect 4522 89734 7912 89786
rect 1104 89712 7912 89734
rect 104052 89786 108836 89808
rect 104052 89734 105922 89786
rect 105974 89734 105986 89786
rect 106038 89734 106050 89786
rect 106102 89734 106114 89786
rect 106166 89734 106178 89786
rect 106230 89734 108836 89786
rect 104052 89712 108836 89734
rect 1104 89242 7912 89264
rect 1104 89190 4874 89242
rect 4926 89190 4938 89242
rect 4990 89190 5002 89242
rect 5054 89190 5066 89242
rect 5118 89190 5130 89242
rect 5182 89190 7912 89242
rect 1104 89168 7912 89190
rect 104052 89242 108836 89264
rect 104052 89190 106658 89242
rect 106710 89190 106722 89242
rect 106774 89190 106786 89242
rect 106838 89190 106850 89242
rect 106902 89190 106914 89242
rect 106966 89190 108836 89242
rect 104052 89168 108836 89190
rect 1104 88698 7912 88720
rect 1104 88646 4214 88698
rect 4266 88646 4278 88698
rect 4330 88646 4342 88698
rect 4394 88646 4406 88698
rect 4458 88646 4470 88698
rect 4522 88646 7912 88698
rect 1104 88624 7912 88646
rect 104052 88698 108836 88720
rect 104052 88646 105922 88698
rect 105974 88646 105986 88698
rect 106038 88646 106050 88698
rect 106102 88646 106114 88698
rect 106166 88646 106178 88698
rect 106230 88646 108836 88698
rect 104052 88624 108836 88646
rect 1104 88154 7912 88176
rect 1104 88102 4874 88154
rect 4926 88102 4938 88154
rect 4990 88102 5002 88154
rect 5054 88102 5066 88154
rect 5118 88102 5130 88154
rect 5182 88102 7912 88154
rect 1104 88080 7912 88102
rect 104052 88154 108836 88176
rect 104052 88102 106658 88154
rect 106710 88102 106722 88154
rect 106774 88102 106786 88154
rect 106838 88102 106850 88154
rect 106902 88102 106914 88154
rect 106966 88102 108836 88154
rect 104052 88080 108836 88102
rect 1104 87610 7912 87632
rect 1104 87558 4214 87610
rect 4266 87558 4278 87610
rect 4330 87558 4342 87610
rect 4394 87558 4406 87610
rect 4458 87558 4470 87610
rect 4522 87558 7912 87610
rect 1104 87536 7912 87558
rect 104052 87610 108836 87632
rect 104052 87558 105922 87610
rect 105974 87558 105986 87610
rect 106038 87558 106050 87610
rect 106102 87558 106114 87610
rect 106166 87558 106178 87610
rect 106230 87558 108836 87610
rect 104052 87536 108836 87558
rect 1104 87066 7912 87088
rect 1104 87014 4874 87066
rect 4926 87014 4938 87066
rect 4990 87014 5002 87066
rect 5054 87014 5066 87066
rect 5118 87014 5130 87066
rect 5182 87014 7912 87066
rect 1104 86992 7912 87014
rect 104052 87066 108836 87088
rect 104052 87014 106658 87066
rect 106710 87014 106722 87066
rect 106774 87014 106786 87066
rect 106838 87014 106850 87066
rect 106902 87014 106914 87066
rect 106966 87014 108836 87066
rect 104052 86992 108836 87014
rect 1104 86522 7912 86544
rect 1104 86470 4214 86522
rect 4266 86470 4278 86522
rect 4330 86470 4342 86522
rect 4394 86470 4406 86522
rect 4458 86470 4470 86522
rect 4522 86470 7912 86522
rect 1104 86448 7912 86470
rect 104052 86522 108836 86544
rect 104052 86470 105922 86522
rect 105974 86470 105986 86522
rect 106038 86470 106050 86522
rect 106102 86470 106114 86522
rect 106166 86470 106178 86522
rect 106230 86470 108836 86522
rect 104052 86448 108836 86470
rect 104437 86411 104495 86417
rect 104437 86377 104449 86411
rect 104483 86408 104495 86411
rect 104710 86408 104716 86420
rect 104483 86380 104716 86408
rect 104483 86377 104495 86380
rect 104437 86371 104495 86377
rect 104710 86368 104716 86380
rect 104768 86368 104774 86420
rect 104529 86139 104587 86145
rect 104529 86105 104541 86139
rect 104575 86136 104587 86139
rect 104802 86136 104808 86148
rect 104575 86108 104808 86136
rect 104575 86105 104587 86108
rect 104529 86099 104587 86105
rect 104802 86096 104808 86108
rect 104860 86096 104866 86148
rect 1104 85978 7912 86000
rect 1104 85926 4874 85978
rect 4926 85926 4938 85978
rect 4990 85926 5002 85978
rect 5054 85926 5066 85978
rect 5118 85926 5130 85978
rect 5182 85926 7912 85978
rect 1104 85904 7912 85926
rect 104052 85978 108836 86000
rect 104052 85926 106658 85978
rect 106710 85926 106722 85978
rect 106774 85926 106786 85978
rect 106838 85926 106850 85978
rect 106902 85926 106914 85978
rect 106966 85926 108836 85978
rect 104052 85904 108836 85926
rect 104529 85731 104587 85737
rect 104529 85697 104541 85731
rect 104575 85728 104587 85731
rect 104710 85728 104716 85740
rect 104575 85700 104716 85728
rect 104575 85697 104587 85700
rect 104529 85691 104587 85697
rect 104710 85688 104716 85700
rect 104768 85688 104774 85740
rect 104621 85663 104679 85669
rect 104621 85629 104633 85663
rect 104667 85660 104679 85663
rect 104802 85660 104808 85672
rect 104667 85632 104808 85660
rect 104667 85629 104679 85632
rect 104621 85623 104679 85629
rect 104802 85620 104808 85632
rect 104860 85620 104866 85672
rect 104897 85595 104955 85601
rect 104897 85561 104909 85595
rect 104943 85592 104955 85595
rect 105814 85592 105820 85604
rect 104943 85564 105820 85592
rect 104943 85561 104955 85564
rect 104897 85555 104955 85561
rect 105814 85552 105820 85564
rect 105872 85552 105878 85604
rect 1104 85434 7912 85456
rect 1104 85382 4214 85434
rect 4266 85382 4278 85434
rect 4330 85382 4342 85434
rect 4394 85382 4406 85434
rect 4458 85382 4470 85434
rect 4522 85382 7912 85434
rect 1104 85360 7912 85382
rect 104052 85434 108836 85456
rect 104052 85382 105922 85434
rect 105974 85382 105986 85434
rect 106038 85382 106050 85434
rect 106102 85382 106114 85434
rect 106166 85382 106178 85434
rect 106230 85382 108836 85434
rect 104052 85360 108836 85382
rect 104434 85280 104440 85332
rect 104492 85320 104498 85332
rect 104713 85323 104771 85329
rect 104713 85320 104725 85323
rect 104492 85292 104725 85320
rect 104492 85280 104498 85292
rect 104713 85289 104725 85292
rect 104759 85289 104771 85323
rect 104713 85283 104771 85289
rect 104529 85119 104587 85125
rect 104529 85085 104541 85119
rect 104575 85116 104587 85119
rect 104710 85116 104716 85128
rect 104575 85088 104716 85116
rect 104575 85085 104587 85088
rect 104529 85079 104587 85085
rect 104710 85076 104716 85088
rect 104768 85076 104774 85128
rect 1104 84890 7912 84912
rect 1104 84838 4874 84890
rect 4926 84838 4938 84890
rect 4990 84838 5002 84890
rect 5054 84838 5066 84890
rect 5118 84838 5130 84890
rect 5182 84838 7912 84890
rect 1104 84816 7912 84838
rect 104052 84890 108836 84912
rect 104052 84838 106658 84890
rect 106710 84838 106722 84890
rect 106774 84838 106786 84890
rect 106838 84838 106850 84890
rect 106902 84838 106914 84890
rect 106966 84838 108836 84890
rect 104052 84816 108836 84838
rect 1104 84346 7912 84368
rect 1104 84294 4214 84346
rect 4266 84294 4278 84346
rect 4330 84294 4342 84346
rect 4394 84294 4406 84346
rect 4458 84294 4470 84346
rect 4522 84294 7912 84346
rect 1104 84272 7912 84294
rect 104052 84346 108836 84368
rect 104052 84294 105922 84346
rect 105974 84294 105986 84346
rect 106038 84294 106050 84346
rect 106102 84294 106114 84346
rect 106166 84294 106178 84346
rect 106230 84294 108836 84346
rect 104052 84272 108836 84294
rect 1104 83802 7912 83824
rect 1104 83750 4874 83802
rect 4926 83750 4938 83802
rect 4990 83750 5002 83802
rect 5054 83750 5066 83802
rect 5118 83750 5130 83802
rect 5182 83750 7912 83802
rect 1104 83728 7912 83750
rect 104052 83802 108836 83824
rect 104052 83750 106658 83802
rect 106710 83750 106722 83802
rect 106774 83750 106786 83802
rect 106838 83750 106850 83802
rect 106902 83750 106914 83802
rect 106966 83750 108836 83802
rect 104052 83728 108836 83750
rect 1104 83258 7912 83280
rect 1104 83206 4214 83258
rect 4266 83206 4278 83258
rect 4330 83206 4342 83258
rect 4394 83206 4406 83258
rect 4458 83206 4470 83258
rect 4522 83206 7912 83258
rect 1104 83184 7912 83206
rect 104052 83258 108836 83280
rect 104052 83206 105922 83258
rect 105974 83206 105986 83258
rect 106038 83206 106050 83258
rect 106102 83206 106114 83258
rect 106166 83206 106178 83258
rect 106230 83206 108836 83258
rect 104052 83184 108836 83206
rect 1104 82714 7912 82736
rect 1104 82662 4874 82714
rect 4926 82662 4938 82714
rect 4990 82662 5002 82714
rect 5054 82662 5066 82714
rect 5118 82662 5130 82714
rect 5182 82662 7912 82714
rect 1104 82640 7912 82662
rect 104052 82714 108836 82736
rect 104052 82662 106658 82714
rect 106710 82662 106722 82714
rect 106774 82662 106786 82714
rect 106838 82662 106850 82714
rect 106902 82662 106914 82714
rect 106966 82662 108836 82714
rect 104052 82640 108836 82662
rect 1104 82170 7912 82192
rect 1104 82118 4214 82170
rect 4266 82118 4278 82170
rect 4330 82118 4342 82170
rect 4394 82118 4406 82170
rect 4458 82118 4470 82170
rect 4522 82118 7912 82170
rect 1104 82096 7912 82118
rect 104052 82170 108836 82192
rect 104052 82118 105922 82170
rect 105974 82118 105986 82170
rect 106038 82118 106050 82170
rect 106102 82118 106114 82170
rect 106166 82118 106178 82170
rect 106230 82118 108836 82170
rect 104052 82096 108836 82118
rect 1104 81626 7912 81648
rect 1104 81574 4874 81626
rect 4926 81574 4938 81626
rect 4990 81574 5002 81626
rect 5054 81574 5066 81626
rect 5118 81574 5130 81626
rect 5182 81574 7912 81626
rect 1104 81552 7912 81574
rect 104052 81626 108836 81648
rect 104052 81574 106658 81626
rect 106710 81574 106722 81626
rect 106774 81574 106786 81626
rect 106838 81574 106850 81626
rect 106902 81574 106914 81626
rect 106966 81574 108836 81626
rect 104052 81552 108836 81574
rect 1104 81082 7912 81104
rect 1104 81030 4214 81082
rect 4266 81030 4278 81082
rect 4330 81030 4342 81082
rect 4394 81030 4406 81082
rect 4458 81030 4470 81082
rect 4522 81030 7912 81082
rect 1104 81008 7912 81030
rect 104052 81082 108836 81104
rect 104052 81030 105922 81082
rect 105974 81030 105986 81082
rect 106038 81030 106050 81082
rect 106102 81030 106114 81082
rect 106166 81030 106178 81082
rect 106230 81030 108836 81082
rect 104052 81008 108836 81030
rect 1104 80538 7912 80560
rect 1104 80486 4874 80538
rect 4926 80486 4938 80538
rect 4990 80486 5002 80538
rect 5054 80486 5066 80538
rect 5118 80486 5130 80538
rect 5182 80486 7912 80538
rect 1104 80464 7912 80486
rect 104052 80538 108836 80560
rect 104052 80486 106658 80538
rect 106710 80486 106722 80538
rect 106774 80486 106786 80538
rect 106838 80486 106850 80538
rect 106902 80486 106914 80538
rect 106966 80486 108836 80538
rect 104052 80464 108836 80486
rect 104158 80248 104164 80300
rect 104216 80288 104222 80300
rect 104345 80291 104403 80297
rect 104345 80288 104357 80291
rect 104216 80260 104357 80288
rect 104216 80248 104222 80260
rect 104345 80257 104357 80260
rect 104391 80288 104403 80291
rect 104621 80291 104679 80297
rect 104621 80288 104633 80291
rect 104391 80260 104633 80288
rect 104391 80257 104403 80260
rect 104345 80251 104403 80257
rect 104621 80257 104633 80260
rect 104667 80257 104679 80291
rect 104621 80251 104679 80257
rect 104437 80087 104495 80093
rect 104437 80053 104449 80087
rect 104483 80084 104495 80087
rect 104526 80084 104532 80096
rect 104483 80056 104532 80084
rect 104483 80053 104495 80056
rect 104437 80047 104495 80053
rect 104526 80044 104532 80056
rect 104584 80044 104590 80096
rect 1104 79994 7912 80016
rect 1104 79942 4214 79994
rect 4266 79942 4278 79994
rect 4330 79942 4342 79994
rect 4394 79942 4406 79994
rect 4458 79942 4470 79994
rect 4522 79942 7912 79994
rect 1104 79920 7912 79942
rect 104052 79994 108836 80016
rect 104052 79942 105922 79994
rect 105974 79942 105986 79994
rect 106038 79942 106050 79994
rect 106102 79942 106114 79994
rect 106166 79942 106178 79994
rect 106230 79942 108836 79994
rect 104052 79920 108836 79942
rect 1104 79450 7912 79472
rect 1104 79398 4874 79450
rect 4926 79398 4938 79450
rect 4990 79398 5002 79450
rect 5054 79398 5066 79450
rect 5118 79398 5130 79450
rect 5182 79398 7912 79450
rect 1104 79376 7912 79398
rect 104052 79450 108836 79472
rect 104052 79398 106658 79450
rect 106710 79398 106722 79450
rect 106774 79398 106786 79450
rect 106838 79398 106850 79450
rect 106902 79398 106914 79450
rect 106966 79398 108836 79450
rect 104052 79376 108836 79398
rect 104066 79092 104072 79144
rect 104124 79132 104130 79144
rect 104529 79135 104587 79141
rect 104529 79132 104541 79135
rect 104124 79104 104541 79132
rect 104124 79092 104130 79104
rect 104529 79101 104541 79104
rect 104575 79132 104587 79135
rect 104897 79135 104955 79141
rect 104897 79132 104909 79135
rect 104575 79104 104909 79132
rect 104575 79101 104587 79104
rect 104529 79095 104587 79101
rect 104897 79101 104909 79104
rect 104943 79132 104955 79135
rect 105170 79132 105176 79144
rect 104943 79104 105176 79132
rect 104943 79101 104955 79104
rect 104897 79095 104955 79101
rect 105170 79092 105176 79104
rect 105228 79092 105234 79144
rect 104713 79067 104771 79073
rect 104713 79064 104725 79067
rect 104452 79036 104725 79064
rect 103882 78956 103888 79008
rect 103940 78996 103946 79008
rect 104452 79005 104480 79036
rect 104713 79033 104725 79036
rect 104759 79033 104771 79067
rect 104713 79027 104771 79033
rect 104437 78999 104495 79005
rect 104437 78996 104449 78999
rect 103940 78968 104449 78996
rect 103940 78956 103946 78968
rect 104437 78965 104449 78968
rect 104483 78965 104495 78999
rect 104437 78959 104495 78965
rect 1104 78906 7912 78928
rect 1104 78854 4214 78906
rect 4266 78854 4278 78906
rect 4330 78854 4342 78906
rect 4394 78854 4406 78906
rect 4458 78854 4470 78906
rect 4522 78854 7912 78906
rect 1104 78832 7912 78854
rect 104052 78906 108836 78928
rect 104052 78854 105922 78906
rect 105974 78854 105986 78906
rect 106038 78854 106050 78906
rect 106102 78854 106114 78906
rect 106166 78854 106178 78906
rect 106230 78854 108836 78906
rect 104052 78832 108836 78854
rect 104618 78752 104624 78804
rect 104676 78792 104682 78804
rect 104989 78795 105047 78801
rect 104989 78792 105001 78795
rect 104676 78764 105001 78792
rect 104676 78752 104682 78764
rect 104989 78761 105001 78764
rect 105035 78761 105047 78795
rect 104989 78755 105047 78761
rect 104434 78665 104440 78668
rect 104417 78659 104440 78665
rect 104417 78625 104429 78659
rect 104417 78619 104440 78625
rect 104434 78616 104440 78619
rect 104492 78616 104498 78668
rect 104636 78628 105492 78656
rect 104250 78548 104256 78600
rect 104308 78588 104314 78600
rect 104636 78597 104664 78628
rect 104621 78591 104679 78597
rect 104621 78588 104633 78591
rect 104308 78560 104633 78588
rect 104308 78548 104314 78560
rect 104621 78557 104633 78560
rect 104667 78557 104679 78591
rect 104897 78591 104955 78597
rect 104897 78588 104909 78591
rect 104621 78551 104679 78557
rect 104728 78560 104909 78588
rect 1302 78480 1308 78532
rect 1360 78520 1366 78532
rect 1489 78523 1547 78529
rect 1489 78520 1501 78523
rect 1360 78492 1501 78520
rect 1360 78480 1366 78492
rect 1489 78489 1501 78492
rect 1535 78489 1547 78523
rect 1489 78483 1547 78489
rect 1673 78523 1731 78529
rect 1673 78489 1685 78523
rect 1719 78520 1731 78523
rect 1857 78523 1915 78529
rect 1857 78520 1869 78523
rect 1719 78492 1869 78520
rect 1719 78489 1731 78492
rect 1673 78483 1731 78489
rect 1857 78489 1869 78492
rect 1903 78520 1915 78523
rect 7558 78520 7564 78532
rect 1903 78492 7564 78520
rect 1903 78489 1915 78492
rect 1857 78483 1915 78489
rect 1504 78452 1532 78483
rect 7558 78480 7564 78492
rect 7616 78480 7622 78532
rect 104066 78480 104072 78532
rect 104124 78520 104130 78532
rect 104345 78523 104403 78529
rect 104345 78520 104357 78523
rect 104124 78492 104357 78520
rect 104124 78480 104130 78492
rect 104345 78489 104357 78492
rect 104391 78489 104403 78523
rect 104728 78520 104756 78560
rect 104897 78557 104909 78560
rect 104943 78557 104955 78591
rect 104897 78551 104955 78557
rect 105170 78548 105176 78600
rect 105228 78548 105234 78600
rect 105464 78597 105492 78628
rect 105449 78591 105507 78597
rect 105449 78557 105461 78591
rect 105495 78557 105507 78591
rect 105449 78551 105507 78557
rect 104345 78483 104403 78489
rect 104636 78492 104756 78520
rect 1949 78455 2007 78461
rect 1949 78452 1961 78455
rect 1504 78424 1961 78452
rect 1949 78421 1961 78424
rect 1995 78421 2007 78455
rect 1949 78415 2007 78421
rect 103882 78412 103888 78464
rect 103940 78452 103946 78464
rect 104529 78455 104587 78461
rect 104529 78452 104541 78455
rect 103940 78424 104541 78452
rect 103940 78412 103946 78424
rect 104529 78421 104541 78424
rect 104575 78452 104587 78455
rect 104636 78452 104664 78492
rect 104802 78480 104808 78532
rect 104860 78520 104866 78532
rect 104860 78492 105308 78520
rect 104860 78480 104866 78492
rect 104575 78424 104664 78452
rect 104575 78421 104587 78424
rect 104529 78415 104587 78421
rect 104710 78412 104716 78464
rect 104768 78412 104774 78464
rect 105280 78461 105308 78492
rect 105265 78455 105323 78461
rect 105265 78421 105277 78455
rect 105311 78421 105323 78455
rect 105265 78415 105323 78421
rect 105538 78412 105544 78464
rect 105596 78412 105602 78464
rect 1104 78362 7912 78384
rect 1104 78310 4874 78362
rect 4926 78310 4938 78362
rect 4990 78310 5002 78362
rect 5054 78310 5066 78362
rect 5118 78310 5130 78362
rect 5182 78310 7912 78362
rect 1104 78288 7912 78310
rect 104052 78362 108836 78384
rect 104052 78310 106658 78362
rect 106710 78310 106722 78362
rect 106774 78310 106786 78362
rect 106838 78310 106850 78362
rect 106902 78310 106914 78362
rect 106966 78310 108836 78362
rect 104052 78288 108836 78310
rect 104434 78208 104440 78260
rect 104492 78248 104498 78260
rect 104618 78248 104624 78260
rect 104492 78220 104624 78248
rect 104492 78208 104498 78220
rect 104618 78208 104624 78220
rect 104676 78248 104682 78260
rect 105538 78248 105544 78260
rect 104676 78220 105544 78248
rect 104676 78208 104682 78220
rect 105538 78208 105544 78220
rect 105596 78208 105602 78260
rect 1302 78072 1308 78124
rect 1360 78112 1366 78124
rect 1489 78115 1547 78121
rect 1489 78112 1501 78115
rect 1360 78084 1501 78112
rect 1360 78072 1366 78084
rect 1489 78081 1501 78084
rect 1535 78112 1547 78115
rect 1949 78115 2007 78121
rect 1949 78112 1961 78115
rect 1535 78084 1961 78112
rect 1535 78081 1547 78084
rect 1489 78075 1547 78081
rect 1949 78081 1961 78084
rect 1995 78081 2007 78115
rect 1949 78075 2007 78081
rect 104345 78115 104403 78121
rect 104345 78081 104357 78115
rect 104391 78112 104403 78115
rect 104434 78112 104440 78124
rect 104391 78084 104440 78112
rect 104391 78081 104403 78084
rect 104345 78075 104403 78081
rect 104434 78072 104440 78084
rect 104492 78072 104498 78124
rect 1673 77979 1731 77985
rect 1673 77945 1685 77979
rect 1719 77976 1731 77979
rect 1857 77979 1915 77985
rect 1857 77976 1869 77979
rect 1719 77948 1869 77976
rect 1719 77945 1731 77948
rect 1673 77939 1731 77945
rect 1857 77945 1869 77948
rect 1903 77976 1915 77979
rect 7650 77976 7656 77988
rect 1903 77948 7656 77976
rect 1903 77945 1915 77948
rect 1857 77939 1915 77945
rect 7650 77936 7656 77948
rect 7708 77936 7714 77988
rect 105630 77868 105636 77920
rect 105688 77908 105694 77920
rect 106185 77911 106243 77917
rect 106185 77908 106197 77911
rect 105688 77880 106197 77908
rect 105688 77868 105694 77880
rect 106185 77877 106197 77880
rect 106231 77908 106243 77911
rect 106274 77908 106280 77920
rect 106231 77880 106280 77908
rect 106231 77877 106243 77880
rect 106185 77871 106243 77877
rect 106274 77868 106280 77880
rect 106332 77868 106338 77920
rect 1104 77818 7912 77840
rect 1104 77766 4214 77818
rect 4266 77766 4278 77818
rect 4330 77766 4342 77818
rect 4394 77766 4406 77818
rect 4458 77766 4470 77818
rect 4522 77766 7912 77818
rect 1104 77744 7912 77766
rect 104052 77818 108836 77840
rect 104052 77766 105922 77818
rect 105974 77766 105986 77818
rect 106038 77766 106050 77818
rect 106102 77766 106114 77818
rect 106166 77766 106178 77818
rect 106230 77766 108836 77818
rect 104052 77744 108836 77766
rect 102778 77460 102784 77512
rect 102836 77500 102842 77512
rect 104345 77503 104403 77509
rect 104345 77500 104357 77503
rect 102836 77472 104357 77500
rect 102836 77460 102842 77472
rect 104345 77469 104357 77472
rect 104391 77500 104403 77503
rect 105081 77503 105139 77509
rect 105081 77500 105093 77503
rect 104391 77472 105093 77500
rect 104391 77469 104403 77472
rect 104345 77463 104403 77469
rect 105081 77469 105093 77472
rect 105127 77500 105139 77503
rect 105630 77500 105636 77512
rect 105127 77472 105636 77500
rect 105127 77469 105139 77472
rect 105081 77463 105139 77469
rect 105630 77460 105636 77472
rect 105688 77460 105694 77512
rect 104434 77324 104440 77376
rect 104492 77364 104498 77376
rect 104897 77367 104955 77373
rect 104897 77364 104909 77367
rect 104492 77336 104909 77364
rect 104492 77324 104498 77336
rect 104897 77333 104909 77336
rect 104943 77333 104955 77367
rect 104897 77327 104955 77333
rect 1104 77274 7912 77296
rect 1104 77222 4874 77274
rect 4926 77222 4938 77274
rect 4990 77222 5002 77274
rect 5054 77222 5066 77274
rect 5118 77222 5130 77274
rect 5182 77222 7912 77274
rect 1104 77200 7912 77222
rect 104052 77274 108836 77296
rect 104052 77222 106658 77274
rect 106710 77222 106722 77274
rect 106774 77222 106786 77274
rect 106838 77222 106850 77274
rect 106902 77222 106914 77274
rect 106966 77222 108836 77274
rect 104052 77200 108836 77222
rect 1210 76984 1216 77036
rect 1268 77024 1274 77036
rect 1489 77027 1547 77033
rect 1489 77024 1501 77027
rect 1268 76996 1501 77024
rect 1268 76984 1274 76996
rect 1489 76993 1501 76996
rect 1535 77024 1547 77027
rect 1949 77027 2007 77033
rect 1949 77024 1961 77027
rect 1535 76996 1961 77024
rect 1535 76993 1547 76996
rect 1489 76987 1547 76993
rect 1949 76993 1961 76996
rect 1995 76993 2007 77027
rect 1949 76987 2007 76993
rect 1673 76891 1731 76897
rect 1673 76857 1685 76891
rect 1719 76888 1731 76891
rect 1857 76891 1915 76897
rect 1857 76888 1869 76891
rect 1719 76860 1869 76888
rect 1719 76857 1731 76860
rect 1673 76851 1731 76857
rect 1857 76857 1869 76860
rect 1903 76888 1915 76891
rect 8938 76888 8944 76900
rect 1903 76860 8944 76888
rect 1903 76857 1915 76860
rect 1857 76851 1915 76857
rect 8938 76848 8944 76860
rect 8996 76848 9002 76900
rect 1104 76730 7912 76752
rect 1104 76678 4214 76730
rect 4266 76678 4278 76730
rect 4330 76678 4342 76730
rect 4394 76678 4406 76730
rect 4458 76678 4470 76730
rect 4522 76678 7912 76730
rect 1104 76656 7912 76678
rect 104052 76730 108836 76752
rect 104052 76678 105922 76730
rect 105974 76678 105986 76730
rect 106038 76678 106050 76730
rect 106102 76678 106114 76730
rect 106166 76678 106178 76730
rect 106230 76678 108836 76730
rect 104052 76656 108836 76678
rect 1210 76304 1216 76356
rect 1268 76344 1274 76356
rect 1489 76347 1547 76353
rect 1489 76344 1501 76347
rect 1268 76316 1501 76344
rect 1268 76304 1274 76316
rect 1489 76313 1501 76316
rect 1535 76313 1547 76347
rect 1489 76307 1547 76313
rect 1673 76347 1731 76353
rect 1673 76313 1685 76347
rect 1719 76344 1731 76347
rect 1857 76347 1915 76353
rect 1857 76344 1869 76347
rect 1719 76316 1869 76344
rect 1719 76313 1731 76316
rect 1673 76307 1731 76313
rect 1857 76313 1869 76316
rect 1903 76344 1915 76347
rect 8846 76344 8852 76356
rect 1903 76316 8852 76344
rect 1903 76313 1915 76316
rect 1857 76307 1915 76313
rect 1504 76276 1532 76307
rect 8846 76304 8852 76316
rect 8904 76304 8910 76356
rect 1949 76279 2007 76285
rect 1949 76276 1961 76279
rect 1504 76248 1961 76276
rect 1949 76245 1961 76248
rect 1995 76245 2007 76279
rect 1949 76239 2007 76245
rect 1104 76186 7912 76208
rect 1104 76134 4874 76186
rect 4926 76134 4938 76186
rect 4990 76134 5002 76186
rect 5054 76134 5066 76186
rect 5118 76134 5130 76186
rect 5182 76134 7912 76186
rect 1104 76112 7912 76134
rect 104052 76186 108836 76208
rect 104052 76134 106658 76186
rect 106710 76134 106722 76186
rect 106774 76134 106786 76186
rect 106838 76134 106850 76186
rect 106902 76134 106914 76186
rect 106966 76134 108836 76186
rect 104052 76112 108836 76134
rect 1581 76075 1639 76081
rect 1581 76041 1593 76075
rect 1627 76072 1639 76075
rect 5534 76072 5540 76084
rect 1627 76044 5540 76072
rect 1627 76041 1639 76044
rect 1581 76035 1639 76041
rect 5534 76032 5540 76044
rect 5592 76032 5598 76084
rect 104250 76032 104256 76084
rect 104308 76072 104314 76084
rect 104345 76075 104403 76081
rect 104345 76072 104357 76075
rect 104308 76044 104357 76072
rect 104308 76032 104314 76044
rect 104345 76041 104357 76044
rect 104391 76041 104403 76075
rect 104345 76035 104403 76041
rect 106185 76075 106243 76081
rect 106185 76041 106197 76075
rect 106231 76072 106243 76075
rect 106274 76072 106280 76084
rect 106231 76044 106280 76072
rect 106231 76041 106243 76044
rect 106185 76035 106243 76041
rect 104526 75964 104532 76016
rect 104584 76004 104590 76016
rect 104584 75976 104650 76004
rect 104584 75964 104590 75976
rect 1394 75896 1400 75948
rect 1452 75936 1458 75948
rect 1673 75939 1731 75945
rect 1673 75936 1685 75939
rect 1452 75908 1685 75936
rect 1452 75896 1458 75908
rect 1673 75905 1685 75908
rect 1719 75905 1731 75939
rect 1673 75899 1731 75905
rect 106093 75939 106151 75945
rect 106093 75905 106105 75939
rect 106139 75936 106151 75939
rect 106200 75936 106228 76035
rect 106274 76032 106280 76044
rect 106332 76032 106338 76084
rect 106139 75908 106228 75936
rect 106139 75905 106151 75908
rect 106093 75899 106151 75905
rect 105814 75828 105820 75880
rect 105872 75828 105878 75880
rect 1104 75642 7912 75664
rect 1104 75590 4214 75642
rect 4266 75590 4278 75642
rect 4330 75590 4342 75642
rect 4394 75590 4406 75642
rect 4458 75590 4470 75642
rect 4522 75590 7912 75642
rect 1104 75568 7912 75590
rect 104052 75642 108836 75664
rect 104052 75590 105922 75642
rect 105974 75590 105986 75642
rect 106038 75590 106050 75642
rect 106102 75590 106114 75642
rect 106166 75590 106178 75642
rect 106230 75590 108836 75642
rect 104052 75568 108836 75590
rect 104250 75284 104256 75336
rect 104308 75324 104314 75336
rect 104529 75327 104587 75333
rect 104529 75324 104541 75327
rect 104308 75296 104541 75324
rect 104308 75284 104314 75296
rect 104529 75293 104541 75296
rect 104575 75293 104587 75327
rect 104529 75287 104587 75293
rect 1302 75216 1308 75268
rect 1360 75256 1366 75268
rect 1489 75259 1547 75265
rect 1489 75256 1501 75259
rect 1360 75228 1501 75256
rect 1360 75216 1366 75228
rect 1489 75225 1501 75228
rect 1535 75225 1547 75259
rect 1489 75219 1547 75225
rect 1673 75259 1731 75265
rect 1673 75225 1685 75259
rect 1719 75256 1731 75259
rect 1857 75259 1915 75265
rect 1857 75256 1869 75259
rect 1719 75228 1869 75256
rect 1719 75225 1731 75228
rect 1673 75219 1731 75225
rect 1857 75225 1869 75228
rect 1903 75256 1915 75259
rect 6914 75256 6920 75268
rect 1903 75228 6920 75256
rect 1903 75225 1915 75228
rect 1857 75219 1915 75225
rect 1504 75188 1532 75219
rect 6914 75216 6920 75228
rect 6972 75216 6978 75268
rect 1949 75191 2007 75197
rect 1949 75188 1961 75191
rect 1504 75160 1961 75188
rect 1949 75157 1961 75160
rect 1995 75157 2007 75191
rect 1949 75151 2007 75157
rect 102042 75148 102048 75200
rect 102100 75188 102106 75200
rect 104345 75191 104403 75197
rect 104345 75188 104357 75191
rect 102100 75160 104357 75188
rect 102100 75148 102106 75160
rect 104345 75157 104357 75160
rect 104391 75188 104403 75191
rect 104621 75191 104679 75197
rect 104621 75188 104633 75191
rect 104391 75160 104633 75188
rect 104391 75157 104403 75160
rect 104345 75151 104403 75157
rect 104621 75157 104633 75160
rect 104667 75157 104679 75191
rect 104621 75151 104679 75157
rect 1104 75098 7912 75120
rect 1104 75046 4874 75098
rect 4926 75046 4938 75098
rect 4990 75046 5002 75098
rect 5054 75046 5066 75098
rect 5118 75046 5130 75098
rect 5182 75046 7912 75098
rect 1104 75024 7912 75046
rect 104052 75098 108836 75120
rect 104052 75046 106658 75098
rect 106710 75046 106722 75098
rect 106774 75046 106786 75098
rect 106838 75046 106850 75098
rect 106902 75046 106914 75098
rect 106966 75046 108836 75098
rect 104052 75024 108836 75046
rect 1104 74554 7912 74576
rect 1104 74502 4214 74554
rect 4266 74502 4278 74554
rect 4330 74502 4342 74554
rect 4394 74502 4406 74554
rect 4458 74502 4470 74554
rect 4522 74502 7912 74554
rect 1104 74480 7912 74502
rect 104052 74554 108836 74576
rect 104052 74502 105922 74554
rect 105974 74502 105986 74554
rect 106038 74502 106050 74554
rect 106102 74502 106114 74554
rect 106166 74502 106178 74554
rect 106230 74502 108836 74554
rect 104052 74480 108836 74502
rect 1210 74128 1216 74180
rect 1268 74168 1274 74180
rect 1489 74171 1547 74177
rect 1489 74168 1501 74171
rect 1268 74140 1501 74168
rect 1268 74128 1274 74140
rect 1489 74137 1501 74140
rect 1535 74168 1547 74171
rect 1949 74171 2007 74177
rect 1949 74168 1961 74171
rect 1535 74140 1961 74168
rect 1535 74137 1547 74140
rect 1489 74131 1547 74137
rect 1949 74137 1961 74140
rect 1995 74137 2007 74171
rect 1949 74131 2007 74137
rect 1581 74103 1639 74109
rect 1581 74069 1593 74103
rect 1627 74100 1639 74103
rect 1854 74100 1860 74112
rect 1627 74072 1860 74100
rect 1627 74069 1639 74072
rect 1581 74063 1639 74069
rect 1854 74060 1860 74072
rect 1912 74060 1918 74112
rect 1104 74010 7912 74032
rect 1104 73958 4874 74010
rect 4926 73958 4938 74010
rect 4990 73958 5002 74010
rect 5054 73958 5066 74010
rect 5118 73958 5130 74010
rect 5182 73958 7912 74010
rect 1104 73936 7912 73958
rect 104052 74010 108836 74032
rect 104052 73958 106658 74010
rect 106710 73958 106722 74010
rect 106774 73958 106786 74010
rect 106838 73958 106850 74010
rect 106902 73958 106914 74010
rect 106966 73958 108836 74010
rect 104052 73936 108836 73958
rect 1302 73720 1308 73772
rect 1360 73760 1366 73772
rect 1397 73763 1455 73769
rect 1397 73760 1409 73763
rect 1360 73732 1409 73760
rect 1360 73720 1366 73732
rect 1397 73729 1409 73732
rect 1443 73760 1455 73763
rect 1949 73763 2007 73769
rect 1949 73760 1961 73763
rect 1443 73732 1961 73760
rect 1443 73729 1455 73732
rect 1397 73723 1455 73729
rect 1949 73729 1961 73732
rect 1995 73729 2007 73763
rect 1949 73723 2007 73729
rect 9122 73720 9128 73772
rect 9180 73760 9186 73772
rect 9582 73760 9588 73772
rect 9180 73732 9588 73760
rect 9180 73720 9186 73732
rect 9582 73720 9588 73732
rect 9640 73720 9646 73772
rect 1581 73627 1639 73633
rect 1581 73593 1593 73627
rect 1627 73624 1639 73627
rect 1857 73627 1915 73633
rect 1857 73624 1869 73627
rect 1627 73596 1869 73624
rect 1627 73593 1639 73596
rect 1581 73587 1639 73593
rect 1857 73593 1869 73596
rect 1903 73624 1915 73627
rect 9582 73624 9588 73636
rect 1903 73596 9588 73624
rect 1903 73593 1915 73596
rect 1857 73587 1915 73593
rect 9582 73584 9588 73596
rect 9640 73584 9646 73636
rect 1104 73466 7912 73488
rect 1104 73414 4214 73466
rect 4266 73414 4278 73466
rect 4330 73414 4342 73466
rect 4394 73414 4406 73466
rect 4458 73414 4470 73466
rect 4522 73414 7912 73466
rect 1104 73392 7912 73414
rect 104052 73466 108836 73488
rect 104052 73414 105922 73466
rect 105974 73414 105986 73466
rect 106038 73414 106050 73466
rect 106102 73414 106114 73466
rect 106166 73414 106178 73466
rect 106230 73414 108836 73466
rect 104052 73392 108836 73414
rect 1673 73219 1731 73225
rect 1673 73185 1685 73219
rect 1719 73216 1731 73219
rect 1857 73219 1915 73225
rect 1857 73216 1869 73219
rect 1719 73188 1869 73216
rect 1719 73185 1731 73188
rect 1673 73179 1731 73185
rect 1857 73185 1869 73188
rect 1903 73216 1915 73219
rect 9030 73216 9036 73228
rect 1903 73188 9036 73216
rect 1903 73185 1915 73188
rect 1857 73179 1915 73185
rect 9030 73176 9036 73188
rect 9088 73176 9094 73228
rect 1486 73040 1492 73092
rect 1544 73080 1550 73092
rect 1949 73083 2007 73089
rect 1949 73080 1961 73083
rect 1544 73052 1961 73080
rect 1544 73040 1550 73052
rect 1949 73049 1961 73052
rect 1995 73049 2007 73083
rect 1949 73043 2007 73049
rect 1104 72922 7912 72944
rect 1104 72870 4874 72922
rect 4926 72870 4938 72922
rect 4990 72870 5002 72922
rect 5054 72870 5066 72922
rect 5118 72870 5130 72922
rect 5182 72870 7912 72922
rect 1104 72848 7912 72870
rect 104052 72922 108836 72944
rect 104052 72870 106658 72922
rect 106710 72870 106722 72922
rect 106774 72870 106786 72922
rect 106838 72870 106850 72922
rect 106902 72870 106914 72922
rect 106966 72870 108836 72922
rect 104052 72848 108836 72870
rect 1302 72632 1308 72684
rect 1360 72672 1366 72684
rect 1489 72675 1547 72681
rect 1489 72672 1501 72675
rect 1360 72644 1501 72672
rect 1360 72632 1366 72644
rect 1489 72641 1501 72644
rect 1535 72672 1547 72675
rect 1949 72675 2007 72681
rect 1949 72672 1961 72675
rect 1535 72644 1961 72672
rect 1535 72641 1547 72644
rect 1489 72635 1547 72641
rect 1949 72641 1961 72644
rect 1995 72641 2007 72675
rect 1949 72635 2007 72641
rect 1673 72539 1731 72545
rect 1673 72505 1685 72539
rect 1719 72536 1731 72539
rect 1857 72539 1915 72545
rect 1857 72536 1869 72539
rect 1719 72508 1869 72536
rect 1719 72505 1731 72508
rect 1673 72499 1731 72505
rect 1857 72505 1869 72508
rect 1903 72536 1915 72539
rect 9490 72536 9496 72548
rect 1903 72508 9496 72536
rect 1903 72505 1915 72508
rect 1857 72499 1915 72505
rect 9490 72496 9496 72508
rect 9548 72496 9554 72548
rect 1104 72378 7912 72400
rect 1104 72326 4214 72378
rect 4266 72326 4278 72378
rect 4330 72326 4342 72378
rect 4394 72326 4406 72378
rect 4458 72326 4470 72378
rect 4522 72326 7912 72378
rect 1104 72304 7912 72326
rect 104052 72378 108836 72400
rect 104052 72326 105922 72378
rect 105974 72326 105986 72378
rect 106038 72326 106050 72378
rect 106102 72326 106114 72378
rect 106166 72326 106178 72378
rect 106230 72326 108836 72378
rect 104052 72304 108836 72326
rect 1104 71834 7912 71856
rect 1104 71782 4874 71834
rect 4926 71782 4938 71834
rect 4990 71782 5002 71834
rect 5054 71782 5066 71834
rect 5118 71782 5130 71834
rect 5182 71782 7912 71834
rect 1104 71760 7912 71782
rect 104052 71834 108836 71856
rect 104052 71782 106658 71834
rect 106710 71782 106722 71834
rect 106774 71782 106786 71834
rect 106838 71782 106850 71834
rect 106902 71782 106914 71834
rect 106966 71782 108836 71834
rect 104052 71760 108836 71782
rect 1854 71680 1860 71732
rect 1912 71720 1918 71732
rect 9398 71720 9404 71732
rect 1912 71692 9404 71720
rect 1912 71680 1918 71692
rect 9398 71680 9404 71692
rect 9456 71680 9462 71732
rect 1210 71544 1216 71596
rect 1268 71584 1274 71596
rect 1489 71587 1547 71593
rect 1489 71584 1501 71587
rect 1268 71556 1501 71584
rect 1268 71544 1274 71556
rect 1489 71553 1501 71556
rect 1535 71584 1547 71587
rect 1949 71587 2007 71593
rect 1949 71584 1961 71587
rect 1535 71556 1961 71584
rect 1535 71553 1547 71556
rect 1489 71547 1547 71553
rect 1949 71553 1961 71556
rect 1995 71553 2007 71587
rect 1949 71547 2007 71553
rect 1581 71383 1639 71389
rect 1581 71349 1593 71383
rect 1627 71380 1639 71383
rect 1854 71380 1860 71392
rect 1627 71352 1860 71380
rect 1627 71349 1639 71352
rect 1581 71343 1639 71349
rect 1854 71340 1860 71352
rect 1912 71340 1918 71392
rect 1104 71290 7912 71312
rect 1104 71238 4214 71290
rect 4266 71238 4278 71290
rect 4330 71238 4342 71290
rect 4394 71238 4406 71290
rect 4458 71238 4470 71290
rect 4522 71238 7912 71290
rect 1104 71216 7912 71238
rect 104052 71290 108836 71312
rect 104052 71238 105922 71290
rect 105974 71238 105986 71290
rect 106038 71238 106050 71290
rect 106102 71238 106114 71290
rect 106166 71238 106178 71290
rect 106230 71238 108836 71290
rect 104052 71216 108836 71238
rect 1673 70975 1731 70981
rect 1673 70941 1685 70975
rect 1719 70972 1731 70975
rect 1857 70975 1915 70981
rect 1857 70972 1869 70975
rect 1719 70944 1869 70972
rect 1719 70941 1731 70944
rect 1673 70935 1731 70941
rect 1857 70941 1869 70944
rect 1903 70972 1915 70975
rect 9214 70972 9220 70984
rect 1903 70944 9220 70972
rect 1903 70941 1915 70944
rect 1857 70935 1915 70941
rect 9214 70932 9220 70944
rect 9272 70932 9278 70984
rect 1302 70864 1308 70916
rect 1360 70904 1366 70916
rect 1489 70907 1547 70913
rect 1489 70904 1501 70907
rect 1360 70876 1501 70904
rect 1360 70864 1366 70876
rect 1489 70873 1501 70876
rect 1535 70904 1547 70907
rect 2133 70907 2191 70913
rect 2133 70904 2145 70907
rect 1535 70876 2145 70904
rect 1535 70873 1547 70876
rect 1489 70867 1547 70873
rect 2133 70873 2145 70876
rect 2179 70873 2191 70907
rect 2133 70867 2191 70873
rect 2041 70839 2099 70845
rect 2041 70805 2053 70839
rect 2087 70836 2099 70839
rect 2222 70836 2228 70848
rect 2087 70808 2228 70836
rect 2087 70805 2099 70808
rect 2041 70799 2099 70805
rect 2222 70796 2228 70808
rect 2280 70796 2286 70848
rect 1104 70746 7912 70768
rect 1104 70694 4874 70746
rect 4926 70694 4938 70746
rect 4990 70694 5002 70746
rect 5054 70694 5066 70746
rect 5118 70694 5130 70746
rect 5182 70694 7912 70746
rect 1104 70672 7912 70694
rect 104052 70746 108836 70768
rect 104052 70694 106658 70746
rect 106710 70694 106722 70746
rect 106774 70694 106786 70746
rect 106838 70694 106850 70746
rect 106902 70694 106914 70746
rect 106966 70694 108836 70746
rect 104052 70672 108836 70694
rect 1949 70499 2007 70505
rect 1949 70465 1961 70499
rect 1995 70496 2007 70499
rect 1995 70468 2452 70496
rect 1995 70465 2007 70468
rect 1949 70459 2007 70465
rect 2222 70388 2228 70440
rect 2280 70388 2286 70440
rect 2424 70437 2452 70468
rect 2409 70431 2467 70437
rect 2409 70397 2421 70431
rect 2455 70428 2467 70431
rect 8386 70428 8392 70440
rect 2455 70400 8392 70428
rect 2455 70397 2467 70400
rect 2409 70391 2467 70397
rect 8386 70388 8392 70400
rect 8444 70388 8450 70440
rect 1104 70202 7912 70224
rect 1104 70150 4214 70202
rect 4266 70150 4278 70202
rect 4330 70150 4342 70202
rect 4394 70150 4406 70202
rect 4458 70150 4470 70202
rect 4522 70150 7912 70202
rect 1104 70128 7912 70150
rect 104052 70202 108836 70224
rect 104052 70150 105922 70202
rect 105974 70150 105986 70202
rect 106038 70150 106050 70202
rect 106102 70150 106114 70202
rect 106166 70150 106178 70202
rect 106230 70150 108836 70202
rect 104052 70128 108836 70150
rect 1854 69980 1860 70032
rect 1912 70020 1918 70032
rect 38654 70020 38660 70032
rect 1912 69992 38660 70020
rect 1912 69980 1918 69992
rect 38654 69980 38660 69992
rect 38712 69980 38718 70032
rect 73614 69980 73620 70032
rect 73672 70020 73678 70032
rect 103698 70020 103704 70032
rect 73672 69992 103704 70020
rect 73672 69980 73678 69992
rect 103698 69980 103704 69992
rect 103756 69980 103762 70032
rect 9582 69912 9588 69964
rect 9640 69952 9646 69964
rect 43254 69952 43260 69964
rect 9640 69924 43260 69952
rect 9640 69912 9646 69924
rect 43254 69912 43260 69924
rect 43312 69912 43318 69964
rect 71774 69912 71780 69964
rect 71832 69952 71838 69964
rect 102686 69952 102692 69964
rect 71832 69924 102692 69952
rect 71832 69912 71838 69924
rect 102686 69912 102692 69924
rect 102744 69912 102750 69964
rect 9030 69844 9036 69896
rect 9088 69884 9094 69896
rect 40954 69884 40960 69896
rect 9088 69856 40960 69884
rect 9088 69844 9094 69856
rect 40954 69844 40960 69856
rect 41012 69844 41018 69896
rect 70946 69844 70952 69896
rect 71004 69884 71010 69896
rect 103606 69884 103612 69896
rect 71004 69856 103612 69884
rect 71004 69844 71010 69856
rect 103606 69844 103612 69856
rect 103664 69844 103670 69896
rect 108301 69887 108359 69893
rect 108301 69884 108313 69887
rect 108132 69856 108313 69884
rect 1302 69776 1308 69828
rect 1360 69816 1366 69828
rect 1489 69819 1547 69825
rect 1489 69816 1501 69819
rect 1360 69788 1501 69816
rect 1360 69776 1366 69788
rect 1489 69785 1501 69788
rect 1535 69785 1547 69819
rect 1489 69779 1547 69785
rect 1673 69819 1731 69825
rect 1673 69785 1685 69819
rect 1719 69816 1731 69819
rect 1857 69819 1915 69825
rect 1857 69816 1869 69819
rect 1719 69788 1869 69816
rect 1719 69785 1731 69788
rect 1673 69779 1731 69785
rect 1857 69785 1869 69788
rect 1903 69816 1915 69819
rect 1903 69788 6914 69816
rect 1903 69785 1915 69788
rect 1857 69779 1915 69785
rect 1504 69748 1532 69779
rect 1949 69751 2007 69757
rect 1949 69748 1961 69751
rect 1504 69720 1961 69748
rect 1949 69717 1961 69720
rect 1995 69717 2007 69751
rect 6886 69748 6914 69788
rect 9490 69776 9496 69828
rect 9548 69816 9554 69828
rect 39758 69816 39764 69828
rect 9548 69788 39764 69816
rect 9548 69776 9554 69788
rect 39758 69776 39764 69788
rect 39816 69776 39822 69828
rect 69290 69776 69296 69828
rect 69348 69816 69354 69828
rect 102502 69816 102508 69828
rect 69348 69788 102508 69816
rect 69348 69776 69354 69788
rect 102502 69776 102508 69788
rect 102560 69776 102566 69828
rect 37458 69748 37464 69760
rect 6886 69720 37464 69748
rect 1949 69711 2007 69717
rect 37458 69708 37464 69720
rect 37516 69708 37522 69760
rect 68462 69708 68468 69760
rect 68520 69748 68526 69760
rect 102594 69748 102600 69760
rect 68520 69720 102600 69748
rect 68520 69708 68526 69720
rect 102594 69708 102600 69720
rect 102652 69708 102658 69760
rect 107562 69708 107568 69760
rect 107620 69748 107626 69760
rect 108132 69757 108160 69856
rect 108301 69853 108313 69856
rect 108347 69853 108359 69887
rect 108301 69847 108359 69853
rect 108117 69751 108175 69757
rect 108117 69748 108129 69751
rect 107620 69720 108129 69748
rect 107620 69708 107626 69720
rect 108117 69717 108129 69720
rect 108163 69717 108175 69751
rect 108117 69711 108175 69717
rect 108482 69708 108488 69760
rect 108540 69708 108546 69760
rect 1104 69658 7912 69680
rect 1104 69606 4874 69658
rect 4926 69606 4938 69658
rect 4990 69606 5002 69658
rect 5054 69606 5066 69658
rect 5118 69606 5130 69658
rect 5182 69606 7912 69658
rect 66990 69640 66996 69692
rect 67048 69680 67054 69692
rect 103514 69680 103520 69692
rect 67048 69652 103520 69680
rect 67048 69640 67054 69652
rect 103514 69640 103520 69652
rect 103572 69640 103578 69692
rect 104052 69658 108836 69680
rect 1104 69584 7912 69606
rect 104052 69606 106658 69658
rect 106710 69606 106722 69658
rect 106774 69606 106786 69658
rect 106838 69606 106850 69658
rect 106902 69606 106914 69658
rect 106966 69606 108836 69658
rect 104052 69584 108836 69606
rect 7650 69504 7656 69556
rect 7708 69544 7714 69556
rect 32858 69544 32864 69556
rect 7708 69516 32864 69544
rect 7708 69504 7714 69516
rect 32858 69504 32864 69516
rect 32916 69504 32922 69556
rect 7558 69436 7564 69488
rect 7616 69476 7622 69488
rect 36354 69476 36360 69488
rect 7616 69448 36360 69476
rect 7616 69436 7622 69448
rect 36354 69436 36360 69448
rect 36412 69436 36418 69488
rect 6914 69368 6920 69420
rect 6972 69408 6978 69420
rect 35158 69408 35164 69420
rect 6972 69380 35164 69408
rect 6972 69368 6978 69380
rect 35158 69368 35164 69380
rect 35216 69368 35222 69420
rect 1104 69114 7912 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 7912 69114
rect 1104 69040 7912 69062
rect 104052 69114 108836 69136
rect 104052 69062 105922 69114
rect 105974 69062 105986 69114
rect 106038 69062 106050 69114
rect 106102 69062 106114 69114
rect 106166 69062 106178 69114
rect 106230 69062 108836 69114
rect 104052 69040 108836 69062
rect 88610 68756 88616 68808
rect 88668 68796 88674 68808
rect 108117 68799 108175 68805
rect 108117 68796 108129 68799
rect 88668 68768 108129 68796
rect 88668 68756 88674 68768
rect 108117 68765 108129 68768
rect 108163 68796 108175 68799
rect 108301 68799 108359 68805
rect 108301 68796 108313 68799
rect 108163 68768 108313 68796
rect 108163 68765 108175 68768
rect 108117 68759 108175 68765
rect 108301 68765 108313 68768
rect 108347 68765 108359 68799
rect 108301 68759 108359 68765
rect 1210 68688 1216 68740
rect 1268 68728 1274 68740
rect 1489 68731 1547 68737
rect 1489 68728 1501 68731
rect 1268 68700 1501 68728
rect 1268 68688 1274 68700
rect 1489 68697 1501 68700
rect 1535 68697 1547 68731
rect 1489 68691 1547 68697
rect 1673 68731 1731 68737
rect 1673 68697 1685 68731
rect 1719 68728 1731 68731
rect 1857 68731 1915 68737
rect 1857 68728 1869 68731
rect 1719 68700 1869 68728
rect 1719 68697 1731 68700
rect 1673 68691 1731 68697
rect 1857 68697 1869 68700
rect 1903 68728 1915 68731
rect 1903 68700 6914 68728
rect 1903 68697 1915 68700
rect 1857 68691 1915 68697
rect 1504 68660 1532 68691
rect 1949 68663 2007 68669
rect 1949 68660 1961 68663
rect 1504 68632 1961 68660
rect 1949 68629 1961 68632
rect 1995 68629 2007 68663
rect 6886 68660 6914 68700
rect 95878 68688 95884 68740
rect 95936 68728 95942 68740
rect 95936 68700 103836 68728
rect 95936 68688 95942 68700
rect 42150 68660 42156 68672
rect 6886 68632 42156 68660
rect 1949 68623 2007 68629
rect 42150 68620 42156 68632
rect 42208 68620 42214 68672
rect 97166 68620 97172 68672
rect 97224 68660 97230 68672
rect 103698 68660 103704 68672
rect 97224 68632 103704 68660
rect 97224 68620 97230 68632
rect 103698 68620 103704 68632
rect 103756 68620 103762 68672
rect 1104 68570 7912 68592
rect 1104 68518 4874 68570
rect 4926 68518 4938 68570
rect 4990 68518 5002 68570
rect 5054 68518 5066 68570
rect 5118 68518 5130 68570
rect 5182 68518 7912 68570
rect 1104 68496 7912 68518
rect 7834 68416 7840 68468
rect 7892 68456 7898 68468
rect 33594 68456 33600 68468
rect 7892 68428 33600 68456
rect 7892 68416 7898 68428
rect 33594 68416 33600 68428
rect 33652 68416 33658 68468
rect 103808 68456 103836 68700
rect 108482 68620 108488 68672
rect 108540 68620 108546 68672
rect 104052 68570 108836 68592
rect 104052 68518 106658 68570
rect 106710 68518 106722 68570
rect 106774 68518 106786 68570
rect 106838 68518 106850 68570
rect 106902 68518 106914 68570
rect 106966 68518 108836 68570
rect 104052 68496 108836 68518
rect 103808 68428 108344 68456
rect 7926 68348 7932 68400
rect 7984 68388 7990 68400
rect 33686 68388 33692 68400
rect 7984 68360 33692 68388
rect 7984 68348 7990 68360
rect 33686 68348 33692 68360
rect 33744 68348 33750 68400
rect 88334 68348 88340 68400
rect 88392 68388 88398 68400
rect 93578 68388 93584 68400
rect 88392 68360 93584 68388
rect 88392 68348 88398 68360
rect 93578 68348 93584 68360
rect 93636 68348 93642 68400
rect 1302 68280 1308 68332
rect 1360 68320 1366 68332
rect 1489 68323 1547 68329
rect 1489 68320 1501 68323
rect 1360 68292 1501 68320
rect 1360 68280 1366 68292
rect 1489 68289 1501 68292
rect 1535 68320 1547 68323
rect 1949 68323 2007 68329
rect 1949 68320 1961 68323
rect 1535 68292 1961 68320
rect 1535 68289 1547 68292
rect 1489 68283 1547 68289
rect 1949 68289 1961 68292
rect 1995 68289 2007 68323
rect 1949 68283 2007 68289
rect 9306 68280 9312 68332
rect 9364 68320 9370 68332
rect 35986 68320 35992 68332
rect 9364 68292 35992 68320
rect 9364 68280 9370 68292
rect 35986 68280 35992 68292
rect 36044 68280 36050 68332
rect 90634 68280 90640 68332
rect 90692 68320 90698 68332
rect 95694 68320 95700 68332
rect 90692 68292 95700 68320
rect 90692 68280 90698 68292
rect 95694 68280 95700 68292
rect 95752 68280 95758 68332
rect 108316 68329 108344 68428
rect 105725 68323 105783 68329
rect 105725 68289 105737 68323
rect 105771 68320 105783 68323
rect 108301 68323 108359 68329
rect 105771 68292 105952 68320
rect 105771 68289 105783 68292
rect 105725 68283 105783 68289
rect 2038 68212 2044 68264
rect 2096 68252 2102 68264
rect 2096 68224 16574 68252
rect 2096 68212 2102 68224
rect 1673 68187 1731 68193
rect 1673 68153 1685 68187
rect 1719 68184 1731 68187
rect 1857 68187 1915 68193
rect 1857 68184 1869 68187
rect 1719 68156 1869 68184
rect 1719 68153 1731 68156
rect 1673 68147 1731 68153
rect 1857 68153 1869 68156
rect 1903 68184 1915 68187
rect 16546 68184 16574 68224
rect 89162 68212 89168 68264
rect 89220 68252 89226 68264
rect 89220 68224 93716 68252
rect 89220 68212 89226 68224
rect 30466 68184 30472 68196
rect 1903 68156 6914 68184
rect 16546 68156 30472 68184
rect 1903 68153 1915 68156
rect 1857 68147 1915 68153
rect 6886 68116 6914 68156
rect 30466 68144 30472 68156
rect 30524 68144 30530 68196
rect 90726 68144 90732 68196
rect 90784 68184 90790 68196
rect 91554 68184 91560 68196
rect 90784 68156 91560 68184
rect 90784 68144 90790 68156
rect 91554 68144 91560 68156
rect 91612 68184 91618 68196
rect 93688 68184 93716 68224
rect 94038 68212 94044 68264
rect 94096 68252 94102 68264
rect 103790 68252 103796 68264
rect 94096 68224 103796 68252
rect 94096 68212 94102 68224
rect 103790 68212 103796 68224
rect 103848 68212 103854 68264
rect 96062 68184 96068 68196
rect 91612 68156 93624 68184
rect 93688 68156 96068 68184
rect 91612 68144 91618 68156
rect 25774 68116 25780 68128
rect 6886 68088 25780 68116
rect 25774 68076 25780 68088
rect 25832 68076 25838 68128
rect 88886 68076 88892 68128
rect 88944 68116 88950 68128
rect 93486 68116 93492 68128
rect 88944 68088 93492 68116
rect 88944 68076 88950 68088
rect 93486 68076 93492 68088
rect 93544 68076 93550 68128
rect 93596 68116 93624 68156
rect 96062 68144 96068 68156
rect 96120 68144 96126 68196
rect 102594 68144 102600 68196
rect 102652 68184 102658 68196
rect 105817 68187 105875 68193
rect 105817 68184 105829 68187
rect 102652 68156 105829 68184
rect 102652 68144 102658 68156
rect 105817 68153 105829 68156
rect 105863 68153 105875 68187
rect 105817 68147 105875 68153
rect 95602 68116 95608 68128
rect 93596 68088 95608 68116
rect 95602 68076 95608 68088
rect 95660 68076 95666 68128
rect 96154 68076 96160 68128
rect 96212 68116 96218 68128
rect 103698 68116 103704 68128
rect 96212 68088 103704 68116
rect 96212 68076 96218 68088
rect 103698 68076 103704 68088
rect 103756 68116 103762 68128
rect 104158 68116 104164 68128
rect 103756 68088 104164 68116
rect 103756 68076 103762 68088
rect 104158 68076 104164 68088
rect 104216 68116 104222 68128
rect 105541 68119 105599 68125
rect 105541 68116 105553 68119
rect 104216 68088 105553 68116
rect 104216 68076 104222 68088
rect 105541 68085 105553 68088
rect 105587 68116 105599 68119
rect 105924 68116 105952 68292
rect 108301 68289 108313 68323
rect 108347 68289 108359 68323
rect 108301 68283 108359 68289
rect 105587 68088 105952 68116
rect 105587 68085 105599 68088
rect 105541 68079 105599 68085
rect 108482 68076 108488 68128
rect 108540 68076 108546 68128
rect 1104 68026 108836 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 65654 68026
rect 65706 67974 65718 68026
rect 65770 67974 65782 68026
rect 65834 67974 65846 68026
rect 65898 67974 65910 68026
rect 65962 67974 96374 68026
rect 96426 67974 96438 68026
rect 96490 67974 96502 68026
rect 96554 67974 96566 68026
rect 96618 67974 96630 68026
rect 96682 67974 105922 68026
rect 105974 67974 105986 68026
rect 106038 67974 106050 68026
rect 106102 67974 106114 68026
rect 106166 67974 106178 68026
rect 106230 67974 108836 68026
rect 1104 67952 108836 67974
rect 1581 67915 1639 67921
rect 1581 67881 1593 67915
rect 1627 67912 1639 67915
rect 1857 67915 1915 67921
rect 1857 67912 1869 67915
rect 1627 67884 1869 67912
rect 1627 67881 1639 67884
rect 1581 67875 1639 67881
rect 1857 67881 1869 67884
rect 1903 67912 1915 67915
rect 2038 67912 2044 67924
rect 1903 67884 2044 67912
rect 1903 67881 1915 67884
rect 1857 67875 1915 67881
rect 2038 67872 2044 67884
rect 2096 67872 2102 67924
rect 23474 67912 23480 67924
rect 6886 67884 23480 67912
rect 1670 67804 1676 67856
rect 1728 67844 1734 67856
rect 6886 67844 6914 67884
rect 23474 67872 23480 67884
rect 23532 67872 23538 67924
rect 24670 67872 24676 67924
rect 24728 67872 24734 67924
rect 25774 67872 25780 67924
rect 25832 67912 25838 67924
rect 25869 67915 25927 67921
rect 25869 67912 25881 67915
rect 25832 67884 25881 67912
rect 25832 67872 25838 67884
rect 25869 67881 25881 67884
rect 25915 67881 25927 67915
rect 25869 67875 25927 67881
rect 26970 67872 26976 67924
rect 27028 67872 27034 67924
rect 29546 67872 29552 67924
rect 29604 67872 29610 67924
rect 30466 67872 30472 67924
rect 30524 67872 30530 67924
rect 31754 67872 31760 67924
rect 31812 67872 31818 67924
rect 32858 67872 32864 67924
rect 32916 67872 32922 67924
rect 33962 67872 33968 67924
rect 34020 67872 34026 67924
rect 35158 67872 35164 67924
rect 35216 67872 35222 67924
rect 36354 67872 36360 67924
rect 36412 67872 36418 67924
rect 37458 67872 37464 67924
rect 37516 67872 37522 67924
rect 38654 67872 38660 67924
rect 38712 67872 38718 67924
rect 39758 67872 39764 67924
rect 39816 67912 39822 67924
rect 39853 67915 39911 67921
rect 39853 67912 39865 67915
rect 39816 67884 39865 67912
rect 39816 67872 39822 67884
rect 39853 67881 39865 67884
rect 39899 67881 39911 67915
rect 39853 67875 39911 67881
rect 40954 67872 40960 67924
rect 41012 67912 41018 67924
rect 41049 67915 41107 67921
rect 41049 67912 41061 67915
rect 41012 67884 41061 67912
rect 41012 67872 41018 67884
rect 41049 67881 41061 67884
rect 41095 67881 41107 67915
rect 41049 67875 41107 67881
rect 42150 67872 42156 67924
rect 42208 67872 42214 67924
rect 43254 67872 43260 67924
rect 43312 67912 43318 67924
rect 43349 67915 43407 67921
rect 43349 67912 43361 67915
rect 43312 67884 43361 67912
rect 43312 67872 43318 67884
rect 43349 67881 43361 67884
rect 43395 67881 43407 67915
rect 43349 67875 43407 67881
rect 69750 67872 69756 67924
rect 69808 67872 69814 67924
rect 88334 67872 88340 67924
rect 88392 67872 88398 67924
rect 88886 67872 88892 67924
rect 88944 67872 88950 67924
rect 89162 67872 89168 67924
rect 89220 67872 89226 67924
rect 90177 67915 90235 67921
rect 90177 67881 90189 67915
rect 90223 67912 90235 67915
rect 90637 67915 90695 67921
rect 90637 67912 90649 67915
rect 90223 67884 90649 67912
rect 90223 67881 90235 67884
rect 90177 67875 90235 67881
rect 90637 67881 90649 67884
rect 90683 67912 90695 67915
rect 90726 67912 90732 67924
rect 90683 67884 90732 67912
rect 90683 67881 90695 67884
rect 90637 67875 90695 67881
rect 90726 67872 90732 67884
rect 90784 67872 90790 67924
rect 90818 67872 90824 67924
rect 90876 67912 90882 67924
rect 91925 67915 91983 67921
rect 91925 67912 91937 67915
rect 90876 67884 91937 67912
rect 90876 67872 90882 67884
rect 91925 67881 91937 67884
rect 91971 67881 91983 67915
rect 91925 67875 91983 67881
rect 94130 67872 94136 67924
rect 94188 67912 94194 67924
rect 94271 67915 94329 67921
rect 94271 67912 94283 67915
rect 94188 67884 94283 67912
rect 94188 67872 94194 67884
rect 94271 67881 94283 67884
rect 94317 67912 94329 67915
rect 95050 67912 95056 67924
rect 94317 67884 95056 67912
rect 94317 67881 94329 67884
rect 94271 67875 94329 67881
rect 95050 67872 95056 67884
rect 95108 67872 95114 67924
rect 96341 67915 96399 67921
rect 96341 67881 96353 67915
rect 96387 67912 96399 67915
rect 97166 67912 97172 67924
rect 96387 67884 97172 67912
rect 96387 67881 96399 67884
rect 96341 67875 96399 67881
rect 97166 67872 97172 67884
rect 97224 67872 97230 67924
rect 1728 67816 6914 67844
rect 1728 67804 1734 67816
rect 8386 67804 8392 67856
rect 8444 67844 8450 67856
rect 24688 67844 24716 67872
rect 8444 67816 24716 67844
rect 8444 67804 8450 67816
rect 90910 67804 90916 67856
rect 90968 67804 90974 67856
rect 91002 67804 91008 67856
rect 91060 67844 91066 67856
rect 91373 67847 91431 67853
rect 91373 67844 91385 67847
rect 91060 67816 91385 67844
rect 91060 67804 91066 67816
rect 91373 67813 91385 67816
rect 91419 67813 91431 67847
rect 94958 67844 94964 67856
rect 91373 67807 91431 67813
rect 92584 67816 94964 67844
rect 10318 67736 10324 67788
rect 10376 67776 10382 67788
rect 28074 67776 28080 67788
rect 10376 67748 28080 67776
rect 10376 67736 10382 67748
rect 28074 67736 28080 67748
rect 28132 67776 28138 67788
rect 28169 67779 28227 67785
rect 28169 67776 28181 67779
rect 28132 67748 28181 67776
rect 28132 67736 28138 67748
rect 28169 67745 28181 67748
rect 28215 67745 28227 67779
rect 28169 67739 28227 67745
rect 90358 67736 90364 67788
rect 90416 67736 90422 67788
rect 92584 67785 92612 67816
rect 94958 67804 94964 67816
rect 95016 67804 95022 67856
rect 95145 67847 95203 67853
rect 95145 67813 95157 67847
rect 95191 67844 95203 67847
rect 99190 67844 99196 67856
rect 95191 67816 95924 67844
rect 95191 67813 95203 67816
rect 95145 67807 95203 67813
rect 92569 67779 92627 67785
rect 90468 67748 91968 67776
rect 28994 67668 29000 67720
rect 29052 67708 29058 67720
rect 29089 67711 29147 67717
rect 29089 67708 29101 67711
rect 29052 67680 29101 67708
rect 29052 67668 29058 67680
rect 29089 67677 29101 67680
rect 29135 67677 29147 67711
rect 29089 67671 29147 67677
rect 85666 67668 85672 67720
rect 85724 67708 85730 67720
rect 87417 67711 87475 67717
rect 87417 67708 87429 67711
rect 85724 67680 87429 67708
rect 85724 67668 85730 67680
rect 87417 67677 87429 67680
rect 87463 67677 87475 67711
rect 87417 67671 87475 67677
rect 87506 67668 87512 67720
rect 87564 67708 87570 67720
rect 88245 67711 88303 67717
rect 88245 67708 88257 67711
rect 87564 67680 88257 67708
rect 87564 67668 87570 67680
rect 88245 67677 88257 67680
rect 88291 67708 88303 67711
rect 88797 67711 88855 67717
rect 88797 67708 88809 67711
rect 88291 67680 88809 67708
rect 88291 67677 88303 67680
rect 88245 67671 88303 67677
rect 88797 67677 88809 67680
rect 88843 67708 88855 67711
rect 89070 67708 89076 67720
rect 88843 67680 89076 67708
rect 88843 67677 88855 67680
rect 88797 67671 88855 67677
rect 89070 67668 89076 67680
rect 89128 67668 89134 67720
rect 1118 67600 1124 67652
rect 1176 67640 1182 67652
rect 1489 67643 1547 67649
rect 1489 67640 1501 67643
rect 1176 67612 1501 67640
rect 1176 67600 1182 67612
rect 1489 67609 1501 67612
rect 1535 67640 1547 67643
rect 1949 67643 2007 67649
rect 1949 67640 1961 67643
rect 1535 67612 1961 67640
rect 1535 67609 1547 67612
rect 1489 67603 1547 67609
rect 1949 67609 1961 67612
rect 1995 67609 2007 67643
rect 1949 67603 2007 67609
rect 16209 67643 16267 67649
rect 16209 67609 16221 67643
rect 16255 67640 16267 67643
rect 16390 67640 16396 67652
rect 16255 67612 16396 67640
rect 16255 67609 16267 67612
rect 16209 67603 16267 67609
rect 16390 67600 16396 67612
rect 16448 67600 16454 67652
rect 22094 67600 22100 67652
rect 22152 67640 22158 67652
rect 28905 67643 28963 67649
rect 28905 67640 28917 67643
rect 22152 67612 28917 67640
rect 22152 67600 22158 67612
rect 28905 67609 28917 67612
rect 28951 67609 28963 67643
rect 28905 67603 28963 67609
rect 29012 67612 29224 67640
rect 22370 67532 22376 67584
rect 22428 67572 22434 67584
rect 29012 67572 29040 67612
rect 22428 67544 29040 67572
rect 29196 67572 29224 67612
rect 86218 67600 86224 67652
rect 86276 67640 86282 67652
rect 87601 67643 87659 67649
rect 87601 67640 87613 67643
rect 86276 67612 87613 67640
rect 86276 67600 86282 67612
rect 87601 67609 87613 67612
rect 87647 67609 87659 67643
rect 87601 67603 87659 67609
rect 89806 67600 89812 67652
rect 89864 67640 89870 67652
rect 90468 67649 90496 67748
rect 91097 67711 91155 67717
rect 91097 67677 91109 67711
rect 91143 67708 91155 67711
rect 91462 67708 91468 67720
rect 91143 67680 91468 67708
rect 91143 67677 91155 67680
rect 91097 67671 91155 67677
rect 91462 67668 91468 67680
rect 91520 67668 91526 67720
rect 91572 67717 91600 67748
rect 91557 67711 91615 67717
rect 91557 67677 91569 67711
rect 91603 67677 91615 67711
rect 91557 67671 91615 67677
rect 91833 67711 91891 67717
rect 91833 67677 91845 67711
rect 91879 67677 91891 67711
rect 91940 67708 91968 67748
rect 92569 67745 92581 67779
rect 92615 67745 92627 67779
rect 94041 67779 94099 67785
rect 94041 67776 94053 67779
rect 92569 67739 92627 67745
rect 92676 67748 94053 67776
rect 92676 67708 92704 67748
rect 94041 67745 94053 67748
rect 94087 67776 94099 67779
rect 95421 67779 95479 67785
rect 95421 67776 95433 67779
rect 94087 67748 95433 67776
rect 94087 67745 94099 67748
rect 94041 67739 94099 67745
rect 95421 67745 95433 67748
rect 95467 67745 95479 67779
rect 95896 67776 95924 67816
rect 96080 67816 99196 67844
rect 96080 67776 96108 67816
rect 99190 67804 99196 67816
rect 99248 67804 99254 67856
rect 108482 67804 108488 67856
rect 108540 67804 108546 67856
rect 95896 67748 96108 67776
rect 95421 67739 95479 67745
rect 96982 67736 96988 67788
rect 97040 67776 97046 67788
rect 102042 67776 102048 67788
rect 97040 67748 102048 67776
rect 97040 67736 97046 67748
rect 102042 67736 102048 67748
rect 102100 67736 102106 67788
rect 91940 67680 92704 67708
rect 93305 67711 93363 67717
rect 91833 67671 91891 67677
rect 93305 67677 93317 67711
rect 93351 67708 93363 67711
rect 93394 67708 93400 67720
rect 93351 67680 93400 67708
rect 93351 67677 93363 67680
rect 93305 67671 93363 67677
rect 90453 67643 90511 67649
rect 90453 67640 90465 67643
rect 89864 67612 90465 67640
rect 89864 67600 89870 67612
rect 90453 67609 90465 67612
rect 90499 67609 90511 67643
rect 90453 67603 90511 67609
rect 91738 67600 91744 67652
rect 91796 67600 91802 67652
rect 31018 67572 31024 67584
rect 29196 67544 31024 67572
rect 22428 67532 22434 67544
rect 31018 67532 31024 67544
rect 31076 67532 31082 67584
rect 32858 67532 32864 67584
rect 32916 67572 32922 67584
rect 38654 67572 38660 67584
rect 32916 67544 38660 67572
rect 32916 67532 32922 67544
rect 38654 67532 38660 67544
rect 38712 67532 38718 67584
rect 68278 67532 68284 67584
rect 68336 67572 68342 67584
rect 69477 67575 69535 67581
rect 69477 67572 69489 67575
rect 68336 67544 69489 67572
rect 68336 67532 68342 67544
rect 69477 67541 69489 67544
rect 69523 67572 69535 67575
rect 69658 67572 69664 67584
rect 69523 67544 69664 67572
rect 69523 67541 69535 67544
rect 69477 67535 69535 67541
rect 69658 67532 69664 67544
rect 69716 67532 69722 67584
rect 69842 67532 69848 67584
rect 69900 67572 69906 67584
rect 89254 67572 89260 67584
rect 69900 67544 89260 67572
rect 69900 67532 69906 67544
rect 89254 67532 89260 67544
rect 89312 67532 89318 67584
rect 90634 67532 90640 67584
rect 90692 67581 90698 67584
rect 90692 67575 90711 67581
rect 90699 67541 90711 67575
rect 90692 67535 90711 67541
rect 90692 67532 90698 67535
rect 90818 67532 90824 67584
rect 90876 67532 90882 67584
rect 90910 67532 90916 67584
rect 90968 67572 90974 67584
rect 91848 67572 91876 67671
rect 93394 67668 93400 67680
rect 93452 67668 93458 67720
rect 93489 67711 93547 67717
rect 93489 67677 93501 67711
rect 93535 67708 93547 67711
rect 93765 67711 93823 67717
rect 93535 67680 93716 67708
rect 93535 67677 93547 67680
rect 93489 67671 93547 67677
rect 92658 67600 92664 67652
rect 92716 67600 92722 67652
rect 93504 67572 93532 67671
rect 93688 67640 93716 67680
rect 93765 67677 93777 67711
rect 93811 67708 93823 67711
rect 94130 67708 94136 67720
rect 93811 67680 94136 67708
rect 93811 67677 93823 67680
rect 93765 67671 93823 67677
rect 94130 67668 94136 67680
rect 94188 67668 94194 67720
rect 94961 67711 95019 67717
rect 94961 67710 94973 67711
rect 94884 67682 94973 67710
rect 93946 67640 93952 67652
rect 93688 67612 93952 67640
rect 93946 67600 93952 67612
rect 94004 67600 94010 67652
rect 90968 67544 93532 67572
rect 90968 67532 90974 67544
rect 93670 67532 93676 67584
rect 93728 67532 93734 67584
rect 93762 67532 93768 67584
rect 93820 67572 93826 67584
rect 94884 67572 94912 67682
rect 94961 67677 94973 67682
rect 95007 67677 95019 67711
rect 94961 67671 95019 67677
rect 95050 67668 95056 67720
rect 95108 67708 95114 67720
rect 95326 67708 95332 67720
rect 95108 67680 95332 67708
rect 95108 67668 95114 67680
rect 95326 67668 95332 67680
rect 95384 67668 95390 67720
rect 95602 67668 95608 67720
rect 95660 67668 95666 67720
rect 96157 67687 96215 67693
rect 96157 67684 96169 67687
rect 96080 67656 96169 67684
rect 96080 67640 96108 67656
rect 96157 67653 96169 67656
rect 96203 67653 96215 67687
rect 96614 67668 96620 67720
rect 96672 67708 96678 67720
rect 103606 67708 103612 67720
rect 96672 67680 103612 67708
rect 96672 67668 96678 67680
rect 103606 67668 103612 67680
rect 103664 67668 103670 67720
rect 103790 67668 103796 67720
rect 103848 67708 103854 67720
rect 108301 67711 108359 67717
rect 108301 67708 108313 67711
rect 103848 67680 108313 67708
rect 103848 67668 103854 67680
rect 108301 67677 108313 67680
rect 108347 67677 108359 67711
rect 108301 67671 108359 67677
rect 96157 67647 96215 67653
rect 95712 67612 96108 67640
rect 95712 67584 95740 67612
rect 93820 67544 94912 67572
rect 93820 67532 93826 67544
rect 95694 67532 95700 67584
rect 95752 67532 95758 67584
rect 95786 67532 95792 67584
rect 95844 67532 95850 67584
rect 95970 67532 95976 67584
rect 96028 67572 96034 67584
rect 96709 67575 96767 67581
rect 96709 67572 96721 67575
rect 96028 67544 96721 67572
rect 96028 67532 96034 67544
rect 96709 67541 96721 67544
rect 96755 67541 96767 67575
rect 96709 67535 96767 67541
rect 98178 67532 98184 67584
rect 98236 67572 98242 67584
rect 102594 67572 102600 67584
rect 98236 67544 102600 67572
rect 98236 67532 98242 67544
rect 102594 67532 102600 67544
rect 102652 67532 102658 67584
rect 1104 67482 108836 67504
rect 1104 67430 4874 67482
rect 4926 67430 4938 67482
rect 4990 67430 5002 67482
rect 5054 67430 5066 67482
rect 5118 67430 5130 67482
rect 5182 67430 35594 67482
rect 35646 67430 35658 67482
rect 35710 67430 35722 67482
rect 35774 67430 35786 67482
rect 35838 67430 35850 67482
rect 35902 67430 66314 67482
rect 66366 67430 66378 67482
rect 66430 67430 66442 67482
rect 66494 67430 66506 67482
rect 66558 67430 66570 67482
rect 66622 67430 97034 67482
rect 97086 67430 97098 67482
rect 97150 67430 97162 67482
rect 97214 67430 97226 67482
rect 97278 67430 97290 67482
rect 97342 67430 106658 67482
rect 106710 67430 106722 67482
rect 106774 67430 106786 67482
rect 106838 67430 106850 67482
rect 106902 67430 106914 67482
rect 106966 67430 108836 67482
rect 1104 67408 108836 67430
rect 1765 67371 1823 67377
rect 1765 67337 1777 67371
rect 1811 67368 1823 67371
rect 1811 67340 6914 67368
rect 1811 67337 1823 67340
rect 1765 67331 1823 67337
rect 1581 67235 1639 67241
rect 1581 67201 1593 67235
rect 1627 67232 1639 67235
rect 1780 67232 1808 67331
rect 1627 67204 1808 67232
rect 1627 67201 1639 67204
rect 1581 67195 1639 67201
rect 6886 67164 6914 67340
rect 18874 67328 18880 67380
rect 18932 67368 18938 67380
rect 20717 67371 20775 67377
rect 20717 67368 20729 67371
rect 18932 67340 20729 67368
rect 18932 67328 18938 67340
rect 20717 67337 20729 67340
rect 20763 67337 20775 67371
rect 20717 67331 20775 67337
rect 22066 67340 24624 67368
rect 20349 67303 20407 67309
rect 20349 67269 20361 67303
rect 20395 67300 20407 67303
rect 22066 67300 22094 67340
rect 20395 67272 22094 67300
rect 20395 67269 20407 67272
rect 20349 67263 20407 67269
rect 24302 67260 24308 67312
rect 24360 67260 24366 67312
rect 24596 67300 24624 67340
rect 24670 67328 24676 67380
rect 24728 67368 24734 67380
rect 33229 67371 33287 67377
rect 33229 67368 33241 67371
rect 24728 67340 33241 67368
rect 24728 67328 24734 67340
rect 33229 67337 33241 67340
rect 33275 67337 33287 67371
rect 34977 67371 35035 67377
rect 34977 67368 34989 67371
rect 33229 67331 33287 67337
rect 33336 67340 34989 67368
rect 33336 67300 33364 67340
rect 34977 67337 34989 67340
rect 35023 67337 35035 67371
rect 34977 67331 35035 67337
rect 35342 67328 35348 67380
rect 35400 67328 35406 67380
rect 35437 67371 35495 67377
rect 35437 67337 35449 67371
rect 35483 67368 35495 67371
rect 35805 67371 35863 67377
rect 35805 67368 35817 67371
rect 35483 67340 35817 67368
rect 35483 67337 35495 67340
rect 35437 67331 35495 67337
rect 35805 67337 35817 67340
rect 35851 67368 35863 67371
rect 35986 67368 35992 67380
rect 35851 67340 35992 67368
rect 35851 67337 35863 67340
rect 35805 67331 35863 67337
rect 35986 67328 35992 67340
rect 36044 67328 36050 67380
rect 38654 67328 38660 67380
rect 38712 67328 38718 67380
rect 39942 67328 39948 67380
rect 40000 67368 40006 67380
rect 40773 67371 40831 67377
rect 40773 67368 40785 67371
rect 40000 67340 40785 67368
rect 40000 67328 40006 67340
rect 40773 67337 40785 67340
rect 40819 67337 40831 67371
rect 40773 67331 40831 67337
rect 44361 67371 44419 67377
rect 44361 67337 44373 67371
rect 44407 67368 44419 67371
rect 47854 67368 47860 67380
rect 44407 67340 47860 67368
rect 44407 67337 44419 67340
rect 44361 67331 44419 67337
rect 47854 67328 47860 67340
rect 47912 67328 47918 67380
rect 66441 67371 66499 67377
rect 66441 67337 66453 67371
rect 66487 67368 66499 67371
rect 66990 67368 66996 67380
rect 66487 67340 66996 67368
rect 66487 67337 66499 67340
rect 66441 67331 66499 67337
rect 66990 67328 66996 67340
rect 67048 67328 67054 67380
rect 67453 67371 67511 67377
rect 67453 67337 67465 67371
rect 67499 67368 67511 67371
rect 69014 67368 69020 67380
rect 67499 67340 69020 67368
rect 67499 67337 67511 67340
rect 67453 67331 67511 67337
rect 69014 67328 69020 67340
rect 69072 67328 69078 67380
rect 69750 67328 69756 67380
rect 69808 67368 69814 67380
rect 70121 67371 70179 67377
rect 70121 67368 70133 67371
rect 69808 67340 70133 67368
rect 69808 67328 69814 67340
rect 70121 67337 70133 67340
rect 70167 67337 70179 67371
rect 70121 67331 70179 67337
rect 70946 67328 70952 67380
rect 71004 67328 71010 67380
rect 71409 67371 71467 67377
rect 71409 67337 71421 67371
rect 71455 67368 71467 67371
rect 73982 67368 73988 67380
rect 71455 67340 73988 67368
rect 71455 67337 71467 67340
rect 71409 67331 71467 67337
rect 73982 67328 73988 67340
rect 74040 67328 74046 67380
rect 74077 67371 74135 67377
rect 74077 67337 74089 67371
rect 74123 67337 74135 67371
rect 74077 67331 74135 67337
rect 74997 67371 75055 67377
rect 74997 67337 75009 67371
rect 75043 67368 75055 67371
rect 75362 67368 75368 67380
rect 75043 67340 75368 67368
rect 75043 67337 75055 67340
rect 74997 67331 75055 67337
rect 24596 67272 33364 67300
rect 40313 67303 40371 67309
rect 40313 67269 40325 67303
rect 40359 67300 40371 67303
rect 45738 67300 45744 67312
rect 40359 67272 45744 67300
rect 40359 67269 40371 67272
rect 40313 67263 40371 67269
rect 45738 67260 45744 67272
rect 45796 67260 45802 67312
rect 46658 67260 46664 67312
rect 46716 67300 46722 67312
rect 47213 67303 47271 67309
rect 47213 67300 47225 67303
rect 46716 67272 47225 67300
rect 46716 67260 46722 67272
rect 47213 67269 47225 67272
rect 47259 67269 47271 67303
rect 67545 67303 67603 67309
rect 67545 67300 67557 67303
rect 47213 67263 47271 67269
rect 66824 67272 67557 67300
rect 17310 67192 17316 67244
rect 17368 67232 17374 67244
rect 17368 67204 19274 67232
rect 17368 67192 17374 67204
rect 28994 67192 29000 67244
rect 29052 67232 29058 67244
rect 30377 67235 30435 67241
rect 30377 67232 30389 67235
rect 29052 67204 30389 67232
rect 29052 67192 29058 67204
rect 30377 67201 30389 67204
rect 30423 67232 30435 67235
rect 30653 67235 30711 67241
rect 30653 67232 30665 67235
rect 30423 67204 30665 67232
rect 30423 67201 30435 67204
rect 30377 67195 30435 67201
rect 30653 67201 30665 67204
rect 30699 67232 30711 67235
rect 30745 67235 30803 67241
rect 30745 67232 30757 67235
rect 30699 67204 30757 67232
rect 30699 67201 30711 67204
rect 30653 67195 30711 67201
rect 30745 67201 30757 67204
rect 30791 67232 30803 67235
rect 30929 67235 30987 67241
rect 30929 67232 30941 67235
rect 30791 67204 30941 67232
rect 30791 67201 30803 67204
rect 30745 67195 30803 67201
rect 30929 67201 30941 67204
rect 30975 67232 30987 67235
rect 31202 67232 31208 67244
rect 30975 67204 31208 67232
rect 30975 67201 30987 67204
rect 30929 67195 30987 67201
rect 31202 67192 31208 67204
rect 31260 67232 31266 67244
rect 32766 67232 32772 67244
rect 31260 67204 32772 67232
rect 31260 67192 31266 67204
rect 32766 67192 32772 67204
rect 32824 67192 32830 67244
rect 33502 67192 33508 67244
rect 33560 67232 33566 67244
rect 33597 67235 33655 67241
rect 33597 67232 33609 67235
rect 33560 67204 33609 67232
rect 33560 67192 33566 67204
rect 33597 67201 33609 67204
rect 33643 67201 33655 67235
rect 33597 67195 33655 67201
rect 33686 67192 33692 67244
rect 33744 67232 33750 67244
rect 34057 67235 34115 67241
rect 34057 67232 34069 67235
rect 33744 67204 34069 67232
rect 33744 67192 33750 67204
rect 34057 67201 34069 67204
rect 34103 67201 34115 67235
rect 34057 67195 34115 67201
rect 39022 67192 39028 67244
rect 39080 67192 39086 67244
rect 39485 67235 39543 67241
rect 39485 67232 39497 67235
rect 39132 67204 39497 67232
rect 39132 67176 39160 67204
rect 39485 67201 39497 67204
rect 39531 67201 39543 67235
rect 39485 67195 39543 67201
rect 39761 67235 39819 67241
rect 39761 67201 39773 67235
rect 39807 67232 39819 67235
rect 41233 67235 41291 67241
rect 41233 67232 41245 67235
rect 39807 67204 41245 67232
rect 39807 67201 39819 67204
rect 39761 67195 39819 67201
rect 20346 67164 20352 67176
rect 6886 67136 20352 67164
rect 20346 67124 20352 67136
rect 20404 67124 20410 67176
rect 20625 67167 20683 67173
rect 20625 67133 20637 67167
rect 20671 67133 20683 67167
rect 20625 67127 20683 67133
rect 24765 67167 24823 67173
rect 24765 67133 24777 67167
rect 24811 67164 24823 67167
rect 24811 67136 24992 67164
rect 24811 67133 24823 67136
rect 24765 67127 24823 67133
rect 842 66988 848 67040
rect 900 67028 906 67040
rect 1397 67031 1455 67037
rect 1397 67028 1409 67031
rect 900 67000 1409 67028
rect 900 66988 906 67000
rect 1397 66997 1409 67000
rect 1443 66997 1455 67031
rect 1397 66991 1455 66997
rect 20254 66988 20260 67040
rect 20312 67028 20318 67040
rect 20640 67028 20668 67127
rect 24964 67096 24992 67136
rect 25038 67124 25044 67176
rect 25096 67124 25102 67176
rect 29086 67124 29092 67176
rect 29144 67164 29150 67176
rect 32950 67164 32956 67176
rect 29144 67136 32956 67164
rect 29144 67124 29150 67136
rect 32950 67124 32956 67136
rect 33008 67124 33014 67176
rect 33873 67167 33931 67173
rect 33873 67133 33885 67167
rect 33919 67164 33931 67167
rect 34238 67164 34244 67176
rect 33919 67136 34244 67164
rect 33919 67133 33931 67136
rect 33873 67127 33931 67133
rect 34238 67124 34244 67136
rect 34296 67164 34302 67176
rect 34333 67167 34391 67173
rect 34333 67164 34345 67167
rect 34296 67136 34345 67164
rect 34296 67124 34302 67136
rect 34333 67133 34345 67136
rect 34379 67164 34391 67167
rect 35621 67167 35679 67173
rect 35621 67164 35633 67167
rect 34379 67136 35633 67164
rect 34379 67133 34391 67136
rect 34333 67127 34391 67133
rect 35621 67133 35633 67136
rect 35667 67164 35679 67167
rect 35667 67136 36124 67164
rect 35667 67133 35679 67136
rect 35621 67127 35679 67133
rect 32858 67096 32864 67108
rect 24964 67068 32864 67096
rect 32858 67056 32864 67068
rect 32916 67056 32922 67108
rect 36096 67105 36124 67136
rect 39114 67124 39120 67176
rect 39172 67124 39178 67176
rect 39301 67167 39359 67173
rect 39301 67164 39313 67167
rect 39224 67136 39313 67164
rect 36081 67099 36139 67105
rect 33060 67068 33824 67096
rect 20901 67031 20959 67037
rect 20901 67028 20913 67031
rect 20312 67000 20913 67028
rect 20312 66988 20318 67000
rect 20901 66997 20913 67000
rect 20947 66997 20959 67031
rect 20901 66991 20959 66997
rect 21266 66988 21272 67040
rect 21324 66988 21330 67040
rect 22002 66988 22008 67040
rect 22060 67028 22066 67040
rect 23109 67031 23167 67037
rect 23109 67028 23121 67031
rect 22060 67000 23121 67028
rect 22060 66988 22066 67000
rect 23109 66997 23121 67000
rect 23155 66997 23167 67031
rect 23109 66991 23167 66997
rect 23290 66988 23296 67040
rect 23348 67028 23354 67040
rect 25133 67031 25191 67037
rect 25133 67028 25145 67031
rect 23348 67000 25145 67028
rect 23348 66988 23354 67000
rect 25133 66997 25145 67000
rect 25179 66997 25191 67031
rect 25133 66991 25191 66997
rect 25774 66988 25780 67040
rect 25832 67028 25838 67040
rect 30285 67031 30343 67037
rect 30285 67028 30297 67031
rect 25832 67000 30297 67028
rect 25832 66988 25838 67000
rect 30285 66997 30297 67000
rect 30331 66997 30343 67031
rect 30285 66991 30343 66997
rect 30558 66988 30564 67040
rect 30616 66988 30622 67040
rect 31018 66988 31024 67040
rect 31076 67028 31082 67040
rect 33060 67028 33088 67068
rect 31076 67000 33088 67028
rect 33137 67031 33195 67037
rect 31076 66988 31082 67000
rect 33137 66997 33149 67031
rect 33183 67028 33195 67031
rect 33502 67028 33508 67040
rect 33183 67000 33508 67028
rect 33183 66997 33195 67000
rect 33137 66991 33195 66997
rect 33502 66988 33508 67000
rect 33560 66988 33566 67040
rect 33796 67028 33824 67068
rect 36081 67065 36093 67099
rect 36127 67096 36139 67099
rect 39224 67096 39252 67136
rect 39301 67133 39313 67136
rect 39347 67164 39359 67167
rect 39776 67164 39804 67195
rect 39347 67136 39804 67164
rect 39347 67133 39359 67136
rect 39301 67127 39359 67133
rect 40402 67124 40408 67176
rect 40460 67124 40466 67176
rect 40604 67173 40632 67204
rect 41233 67201 41245 67204
rect 41279 67232 41291 67235
rect 46569 67235 46627 67241
rect 41279 67204 44588 67232
rect 41279 67201 41291 67204
rect 41233 67195 41291 67201
rect 40589 67167 40647 67173
rect 40589 67133 40601 67167
rect 40635 67133 40647 67167
rect 40589 67127 40647 67133
rect 44450 67124 44456 67176
rect 44508 67124 44514 67176
rect 44560 67173 44588 67204
rect 46569 67201 46581 67235
rect 46615 67232 46627 67235
rect 47486 67232 47492 67244
rect 46615 67204 47492 67232
rect 46615 67201 46627 67204
rect 46569 67195 46627 67201
rect 47486 67192 47492 67204
rect 47544 67192 47550 67244
rect 62025 67235 62083 67241
rect 62025 67201 62037 67235
rect 62071 67232 62083 67235
rect 62390 67232 62396 67244
rect 62071 67204 62396 67232
rect 62071 67201 62083 67204
rect 62025 67195 62083 67201
rect 62390 67192 62396 67204
rect 62448 67192 62454 67244
rect 66824 67173 66852 67272
rect 67545 67269 67557 67272
rect 67591 67269 67603 67303
rect 67545 67263 67603 67269
rect 67913 67303 67971 67309
rect 67913 67269 67925 67303
rect 67959 67300 67971 67303
rect 68462 67300 68468 67312
rect 67959 67272 68468 67300
rect 67959 67269 67971 67272
rect 67913 67263 67971 67269
rect 67085 67235 67143 67241
rect 67085 67201 67097 67235
rect 67131 67201 67143 67235
rect 67085 67195 67143 67201
rect 44545 67167 44603 67173
rect 44545 67133 44557 67167
rect 44591 67164 44603 67167
rect 45005 67167 45063 67173
rect 45005 67164 45017 67167
rect 44591 67136 45017 67164
rect 44591 67133 44603 67136
rect 44545 67127 44603 67133
rect 45005 67133 45017 67136
rect 45051 67164 45063 67167
rect 46845 67167 46903 67173
rect 46845 67164 46857 67167
rect 45051 67136 46857 67164
rect 45051 67133 45063 67136
rect 45005 67127 45063 67133
rect 46845 67133 46857 67136
rect 46891 67164 46903 67167
rect 47673 67167 47731 67173
rect 47673 67164 47685 67167
rect 46891 67136 47685 67164
rect 46891 67133 46903 67136
rect 46845 67127 46903 67133
rect 47673 67133 47685 67136
rect 47719 67164 47731 67167
rect 66809 67167 66867 67173
rect 66809 67164 66821 67167
rect 47719 67136 66821 67164
rect 47719 67133 47731 67136
rect 47673 67127 47731 67133
rect 66809 67133 66821 67136
rect 66855 67133 66867 67167
rect 66809 67127 66867 67133
rect 36127 67068 39252 67096
rect 36127 67065 36139 67068
rect 36081 67059 36139 67065
rect 39390 67056 39396 67108
rect 39448 67096 39454 67108
rect 44468 67096 44496 67124
rect 44821 67099 44879 67105
rect 44821 67096 44833 67099
rect 39448 67068 44128 67096
rect 44468 67068 44833 67096
rect 39448 67056 39454 67068
rect 39942 67028 39948 67040
rect 33796 67000 39948 67028
rect 39942 66988 39948 67000
rect 40000 66988 40006 67040
rect 40402 66988 40408 67040
rect 40460 67028 40466 67040
rect 40957 67031 41015 67037
rect 40957 67028 40969 67031
rect 40460 67000 40969 67028
rect 40460 66988 40466 67000
rect 40957 66997 40969 67000
rect 41003 66997 41015 67031
rect 40957 66991 41015 66997
rect 43990 66988 43996 67040
rect 44048 66988 44054 67040
rect 44100 67028 44128 67068
rect 44821 67065 44833 67068
rect 44867 67065 44879 67099
rect 44821 67059 44879 67065
rect 60734 67056 60740 67108
rect 60792 67096 60798 67108
rect 62206 67096 62212 67108
rect 60792 67068 62212 67096
rect 60792 67056 60798 67068
rect 62206 67056 62212 67068
rect 62264 67056 62270 67108
rect 63402 67056 63408 67108
rect 63460 67096 63466 67108
rect 66533 67099 66591 67105
rect 66533 67096 66545 67099
rect 63460 67068 66545 67096
rect 63460 67056 63466 67068
rect 66533 67065 66545 67068
rect 66579 67096 66591 67099
rect 67100 67096 67128 67195
rect 67560 67164 67588 67263
rect 68462 67260 68468 67272
rect 68520 67260 68526 67312
rect 71041 67303 71099 67309
rect 71041 67300 71053 67303
rect 69400 67272 71053 67300
rect 68554 67192 68560 67244
rect 68612 67192 68618 67244
rect 68278 67164 68284 67176
rect 67560 67136 68284 67164
rect 68278 67124 68284 67136
rect 68336 67124 68342 67176
rect 69400 67164 69428 67272
rect 71041 67269 71053 67272
rect 71087 67269 71099 67303
rect 74092 67300 74120 67331
rect 75362 67328 75368 67340
rect 75420 67328 75426 67380
rect 75454 67328 75460 67380
rect 75512 67328 75518 67380
rect 75822 67328 75828 67380
rect 75880 67328 75886 67380
rect 89346 67368 89352 67380
rect 76116 67340 89352 67368
rect 74261 67303 74319 67309
rect 74261 67300 74273 67303
rect 74092 67272 74273 67300
rect 71041 67263 71099 67269
rect 74261 67269 74273 67272
rect 74307 67300 74319 67303
rect 76116 67300 76144 67340
rect 89346 67328 89352 67340
rect 89404 67328 89410 67380
rect 89548 67340 92060 67368
rect 74307 67272 76144 67300
rect 77021 67303 77079 67309
rect 74307 67269 74319 67272
rect 74261 67263 74319 67269
rect 77021 67269 77033 67303
rect 77067 67300 77079 67303
rect 87785 67303 87843 67309
rect 77067 67272 86066 67300
rect 77067 67269 77079 67272
rect 77021 67263 77079 67269
rect 87785 67269 87797 67303
rect 87831 67300 87843 67303
rect 89548 67300 89576 67340
rect 87831 67272 89576 67300
rect 89640 67272 89746 67300
rect 87831 67269 87843 67272
rect 87785 67263 87843 67269
rect 69474 67192 69480 67244
rect 69532 67232 69538 67244
rect 70213 67235 70271 67241
rect 70213 67232 70225 67235
rect 69532 67204 70225 67232
rect 69532 67192 69538 67204
rect 70213 67201 70225 67204
rect 70259 67201 70271 67235
rect 70213 67195 70271 67201
rect 71774 67192 71780 67244
rect 71832 67192 71838 67244
rect 71866 67192 71872 67244
rect 71924 67232 71930 67244
rect 72329 67235 72387 67241
rect 72329 67232 72341 67235
rect 71924 67204 72341 67232
rect 71924 67192 71930 67204
rect 72329 67201 72341 67204
rect 72375 67201 72387 67235
rect 72329 67195 72387 67201
rect 73157 67235 73215 67241
rect 73157 67201 73169 67235
rect 73203 67232 73215 67235
rect 73614 67232 73620 67244
rect 73203 67204 73620 67232
rect 73203 67201 73215 67204
rect 73157 67195 73215 67201
rect 73614 67192 73620 67204
rect 73672 67192 73678 67244
rect 73706 67192 73712 67244
rect 73764 67192 73770 67244
rect 75638 67232 75644 67244
rect 75288 67204 75644 67232
rect 69661 67167 69719 67173
rect 69661 67164 69673 67167
rect 68848 67136 69673 67164
rect 66579 67068 67128 67096
rect 66579 67065 66591 67068
rect 66533 67059 66591 67065
rect 67542 67056 67548 67108
rect 67600 67096 67606 67108
rect 68848 67096 68876 67136
rect 69661 67133 69673 67136
rect 69707 67133 69719 67167
rect 69661 67127 69719 67133
rect 69750 67124 69756 67176
rect 69808 67164 69814 67176
rect 69934 67164 69940 67176
rect 69808 67136 69940 67164
rect 69808 67124 69814 67136
rect 69934 67124 69940 67136
rect 69992 67124 69998 67176
rect 70026 67124 70032 67176
rect 70084 67164 70090 67176
rect 75288 67173 75316 67204
rect 75638 67192 75644 67204
rect 75696 67192 75702 67244
rect 76190 67192 76196 67244
rect 76248 67232 76254 67244
rect 76561 67235 76619 67241
rect 76561 67232 76573 67235
rect 76248 67204 76573 67232
rect 76248 67192 76254 67204
rect 76561 67201 76573 67204
rect 76607 67232 76619 67235
rect 76929 67235 76987 67241
rect 76929 67232 76941 67235
rect 76607 67204 76941 67232
rect 76607 67201 76619 67204
rect 76561 67195 76619 67201
rect 76929 67201 76941 67204
rect 76975 67232 76987 67235
rect 77297 67235 77355 67241
rect 77297 67232 77309 67235
rect 76975 67204 77309 67232
rect 76975 67201 76987 67204
rect 76929 67195 76987 67201
rect 77297 67201 77309 67204
rect 77343 67232 77355 67235
rect 77386 67232 77392 67244
rect 77343 67204 77392 67232
rect 77343 67201 77355 67204
rect 77297 67195 77355 67201
rect 77386 67192 77392 67204
rect 77444 67192 77450 67244
rect 77570 67192 77576 67244
rect 77628 67232 77634 67244
rect 79321 67235 79379 67241
rect 79321 67232 79333 67235
rect 77628 67204 79333 67232
rect 77628 67192 77634 67204
rect 79321 67201 79333 67204
rect 79367 67201 79379 67235
rect 79321 67195 79379 67201
rect 86954 67192 86960 67244
rect 87012 67232 87018 67244
rect 87141 67235 87199 67241
rect 87141 67232 87153 67235
rect 87012 67204 87153 67232
rect 87012 67192 87018 67204
rect 87141 67201 87153 67204
rect 87187 67232 87199 67235
rect 87506 67232 87512 67244
rect 87187 67204 87512 67232
rect 87187 67201 87199 67204
rect 87141 67195 87199 67201
rect 87506 67192 87512 67204
rect 87564 67232 87570 67244
rect 87693 67235 87751 67241
rect 87693 67232 87705 67235
rect 87564 67204 87705 67232
rect 87564 67192 87570 67204
rect 87693 67201 87705 67204
rect 87739 67232 87751 67235
rect 88061 67235 88119 67241
rect 88061 67232 88073 67235
rect 87739 67204 88073 67232
rect 87739 67201 87751 67204
rect 87693 67195 87751 67201
rect 88061 67201 88073 67204
rect 88107 67201 88119 67235
rect 88061 67195 88119 67201
rect 88429 67235 88487 67241
rect 88429 67201 88441 67235
rect 88475 67232 88487 67235
rect 88518 67232 88524 67244
rect 88475 67204 88524 67232
rect 88475 67201 88487 67204
rect 88429 67195 88487 67201
rect 88518 67192 88524 67204
rect 88576 67192 88582 67244
rect 88610 67192 88616 67244
rect 88668 67192 88674 67244
rect 89254 67192 89260 67244
rect 89312 67232 89318 67244
rect 89530 67232 89536 67244
rect 89312 67204 89536 67232
rect 89312 67192 89318 67204
rect 89530 67192 89536 67204
rect 89588 67192 89594 67244
rect 70857 67167 70915 67173
rect 70857 67164 70869 67167
rect 70084 67136 70869 67164
rect 70084 67124 70090 67136
rect 70857 67133 70869 67136
rect 70903 67164 70915 67167
rect 71685 67167 71743 67173
rect 71685 67164 71697 67167
rect 70903 67136 71697 67164
rect 70903 67133 70915 67136
rect 70857 67127 70915 67133
rect 71685 67133 71697 67136
rect 71731 67164 71743 67167
rect 73525 67167 73583 67173
rect 73525 67164 73537 67167
rect 71731 67136 73537 67164
rect 71731 67133 71743 67136
rect 71685 67127 71743 67133
rect 73525 67133 73537 67136
rect 73571 67164 73583 67167
rect 75273 67167 75331 67173
rect 75273 67164 75285 67167
rect 73571 67136 75285 67164
rect 73571 67133 73583 67136
rect 73525 67127 73583 67133
rect 75273 67133 75285 67136
rect 75319 67133 75331 67167
rect 85206 67164 85212 67176
rect 75273 67127 75331 67133
rect 75380 67136 85212 67164
rect 67600 67068 68876 67096
rect 68925 67099 68983 67105
rect 67600 67056 67606 67068
rect 68925 67065 68937 67099
rect 68971 67096 68983 67099
rect 70394 67096 70400 67108
rect 68971 67068 70400 67096
rect 68971 67065 68983 67068
rect 68925 67059 68983 67065
rect 70394 67056 70400 67068
rect 70452 67056 70458 67108
rect 70578 67056 70584 67108
rect 70636 67056 70642 67108
rect 72237 67099 72295 67105
rect 72237 67065 72249 67099
rect 72283 67096 72295 67099
rect 75380 67096 75408 67136
rect 85206 67124 85212 67136
rect 85264 67124 85270 67176
rect 85301 67167 85359 67173
rect 85301 67133 85313 67167
rect 85347 67133 85359 67167
rect 85301 67127 85359 67133
rect 72283 67068 75408 67096
rect 76285 67099 76343 67105
rect 72283 67065 72295 67068
rect 72237 67059 72295 67065
rect 76285 67065 76297 67099
rect 76331 67096 76343 67099
rect 77938 67096 77944 67108
rect 76331 67068 77944 67096
rect 76331 67065 76343 67068
rect 76285 67059 76343 67065
rect 77938 67056 77944 67068
rect 77996 67056 78002 67108
rect 46201 67031 46259 67037
rect 46201 67028 46213 67031
rect 44100 67000 46213 67028
rect 46201 66997 46213 67000
rect 46247 67028 46259 67031
rect 47029 67031 47087 67037
rect 47029 67028 47041 67031
rect 46247 67000 47041 67028
rect 46247 66997 46259 67000
rect 46201 66991 46259 66997
rect 47029 66997 47041 67000
rect 47075 66997 47087 67031
rect 47029 66991 47087 66997
rect 66162 66988 66168 67040
rect 66220 67028 66226 67040
rect 69474 67028 69480 67040
rect 66220 67000 69480 67028
rect 66220 66988 66226 67000
rect 69474 66988 69480 67000
rect 69532 66988 69538 67040
rect 75638 66988 75644 67040
rect 75696 67028 75702 67040
rect 79137 67031 79195 67037
rect 79137 67028 79149 67031
rect 75696 67000 79149 67028
rect 75696 66988 75702 67000
rect 79137 66997 79149 67000
rect 79183 67028 79195 67031
rect 79778 67028 79784 67040
rect 79183 67000 79784 67028
rect 79183 66997 79195 67000
rect 79137 66991 79195 66997
rect 79778 66988 79784 67000
rect 79836 66988 79842 67040
rect 79870 66988 79876 67040
rect 79928 67028 79934 67040
rect 83090 67028 83096 67040
rect 79928 67000 83096 67028
rect 79928 66988 79934 67000
rect 83090 66988 83096 67000
rect 83148 66988 83154 67040
rect 85316 67028 85344 67127
rect 85574 67124 85580 67176
rect 85632 67124 85638 67176
rect 87233 67167 87291 67173
rect 87233 67133 87245 67167
rect 87279 67164 87291 67167
rect 89640 67164 89668 67272
rect 91554 67260 91560 67312
rect 91612 67260 91618 67312
rect 92032 67300 92060 67340
rect 92106 67328 92112 67380
rect 92164 67368 92170 67380
rect 93302 67368 93308 67380
rect 92164 67340 93308 67368
rect 92164 67328 92170 67340
rect 93302 67328 93308 67340
rect 93360 67368 93366 67380
rect 94041 67371 94099 67377
rect 94041 67368 94053 67371
rect 93360 67340 94053 67368
rect 93360 67328 93366 67340
rect 94041 67337 94053 67340
rect 94087 67368 94099 67371
rect 95786 67368 95792 67380
rect 94087 67340 95792 67368
rect 94087 67337 94099 67340
rect 94041 67331 94099 67337
rect 95786 67328 95792 67340
rect 95844 67328 95850 67380
rect 95878 67328 95884 67380
rect 95936 67328 95942 67380
rect 96706 67328 96712 67380
rect 96764 67368 96770 67380
rect 97169 67371 97227 67377
rect 97169 67368 97181 67371
rect 96764 67340 97181 67368
rect 96764 67328 96770 67340
rect 97169 67337 97181 67340
rect 97215 67368 97227 67371
rect 99653 67371 99711 67377
rect 97215 67340 99512 67368
rect 97215 67337 97227 67340
rect 97169 67331 97227 67337
rect 92032 67272 92782 67300
rect 93578 67260 93584 67312
rect 93636 67300 93642 67312
rect 93636 67272 94898 67300
rect 95988 67272 96936 67300
rect 93636 67260 93642 67272
rect 91189 67235 91247 67241
rect 91189 67201 91201 67235
rect 91235 67232 91247 67235
rect 91373 67235 91431 67241
rect 91373 67232 91385 67235
rect 91235 67204 91385 67232
rect 91235 67201 91247 67204
rect 91189 67195 91247 67201
rect 91373 67201 91385 67204
rect 91419 67232 91431 67235
rect 92014 67232 92020 67244
rect 91419 67204 92020 67232
rect 91419 67201 91431 67204
rect 91373 67195 91431 67201
rect 92014 67192 92020 67204
rect 92072 67192 92078 67244
rect 95988 67241 96016 67272
rect 95973 67235 96031 67241
rect 95973 67201 95985 67235
rect 96019 67201 96031 67235
rect 95973 67195 96031 67201
rect 96157 67235 96215 67241
rect 96157 67201 96169 67235
rect 96203 67232 96215 67235
rect 96706 67232 96712 67244
rect 96203 67204 96712 67232
rect 96203 67201 96215 67204
rect 96157 67195 96215 67201
rect 87279 67136 89668 67164
rect 90913 67167 90971 67173
rect 87279 67133 87291 67136
rect 87233 67127 87291 67133
rect 90913 67133 90925 67167
rect 90959 67164 90971 67167
rect 90959 67136 92152 67164
rect 90959 67133 90971 67136
rect 90913 67127 90971 67133
rect 88426 67096 88432 67108
rect 86972 67068 88432 67096
rect 86218 67028 86224 67040
rect 85316 67000 86224 67028
rect 86218 66988 86224 67000
rect 86276 67028 86282 67040
rect 86972 67028 87000 67068
rect 88426 67056 88432 67068
rect 88484 67096 88490 67108
rect 88797 67099 88855 67105
rect 88797 67096 88809 67099
rect 88484 67068 88809 67096
rect 88484 67056 88490 67068
rect 88797 67065 88809 67068
rect 88843 67065 88855 67099
rect 88797 67059 88855 67065
rect 89441 67099 89499 67105
rect 89441 67065 89453 67099
rect 89487 67096 89499 67099
rect 89806 67096 89812 67108
rect 89487 67068 89812 67096
rect 89487 67065 89499 67068
rect 89441 67059 89499 67065
rect 89806 67056 89812 67068
rect 89864 67056 89870 67108
rect 91388 67068 92060 67096
rect 86276 67000 87000 67028
rect 87049 67031 87107 67037
rect 86276 66988 86282 67000
rect 87049 66997 87061 67031
rect 87095 67028 87107 67031
rect 87509 67031 87567 67037
rect 87509 67028 87521 67031
rect 87095 67000 87521 67028
rect 87095 66997 87107 67000
rect 87049 66991 87107 66997
rect 87509 66997 87521 67000
rect 87555 67028 87567 67031
rect 87598 67028 87604 67040
rect 87555 67000 87604 67028
rect 87555 66997 87567 67000
rect 87509 66991 87567 66997
rect 87598 66988 87604 67000
rect 87656 66988 87662 67040
rect 87782 66988 87788 67040
rect 87840 67028 87846 67040
rect 88153 67031 88211 67037
rect 88153 67028 88165 67031
rect 87840 67000 88165 67028
rect 87840 66988 87846 67000
rect 88153 66997 88165 67000
rect 88199 66997 88211 67031
rect 88153 66991 88211 66997
rect 89346 66988 89352 67040
rect 89404 67028 89410 67040
rect 91388 67028 91416 67068
rect 92032 67040 92060 67068
rect 89404 67000 91416 67028
rect 89404 66988 89410 67000
rect 92014 66988 92020 67040
rect 92072 66988 92078 67040
rect 92124 67028 92152 67136
rect 92290 67124 92296 67176
rect 92348 67124 92354 67176
rect 93762 67124 93768 67176
rect 93820 67124 93826 67176
rect 94133 67167 94191 67173
rect 94133 67133 94145 67167
rect 94179 67164 94191 67167
rect 94409 67167 94467 67173
rect 94179 67136 94268 67164
rect 94179 67133 94191 67136
rect 94133 67127 94191 67133
rect 93394 67056 93400 67108
rect 93452 67096 93458 67108
rect 93780 67096 93808 67124
rect 93452 67068 93808 67096
rect 93452 67056 93458 67068
rect 93670 67028 93676 67040
rect 92124 67000 93676 67028
rect 93670 66988 93676 67000
rect 93728 66988 93734 67040
rect 94240 67028 94268 67136
rect 94409 67133 94421 67167
rect 94455 67164 94467 67167
rect 94498 67164 94504 67176
rect 94455 67136 94504 67164
rect 94455 67133 94467 67136
rect 94409 67127 94467 67133
rect 94498 67124 94504 67136
rect 94556 67124 94562 67176
rect 94774 67124 94780 67176
rect 94832 67164 94838 67176
rect 95988 67164 96016 67195
rect 96706 67192 96712 67204
rect 96764 67192 96770 67244
rect 94832 67136 96016 67164
rect 96065 67167 96123 67173
rect 94832 67124 94838 67136
rect 96065 67133 96077 67167
rect 96111 67164 96123 67167
rect 96798 67164 96804 67176
rect 96111 67136 96804 67164
rect 96111 67133 96123 67136
rect 96065 67127 96123 67133
rect 96798 67124 96804 67136
rect 96856 67124 96862 67176
rect 95528 67068 96292 67096
rect 95528 67028 95556 67068
rect 96264 67040 96292 67068
rect 94240 67000 95556 67028
rect 96246 66988 96252 67040
rect 96304 66988 96310 67040
rect 96525 67031 96583 67037
rect 96525 66997 96537 67031
rect 96571 67028 96583 67031
rect 96706 67028 96712 67040
rect 96571 67000 96712 67028
rect 96571 66997 96583 67000
rect 96525 66991 96583 66997
rect 96706 66988 96712 67000
rect 96764 66988 96770 67040
rect 96908 67028 96936 67272
rect 98178 67260 98184 67312
rect 98236 67260 98242 67312
rect 99374 67300 99380 67312
rect 98932 67272 99380 67300
rect 98932 67241 98960 67272
rect 99374 67260 99380 67272
rect 99432 67260 99438 67312
rect 98917 67235 98975 67241
rect 98917 67201 98929 67235
rect 98963 67201 98975 67235
rect 98917 67195 98975 67201
rect 99190 67192 99196 67244
rect 99248 67192 99254 67244
rect 99484 67241 99512 67340
rect 99653 67337 99665 67371
rect 99699 67337 99711 67371
rect 99653 67331 99711 67337
rect 99668 67300 99696 67331
rect 99742 67328 99748 67380
rect 99800 67368 99806 67380
rect 99837 67371 99895 67377
rect 99837 67368 99849 67371
rect 99800 67340 99849 67368
rect 99800 67328 99806 67340
rect 99837 67337 99849 67340
rect 99883 67368 99895 67371
rect 102778 67368 102784 67380
rect 99883 67340 102784 67368
rect 99883 67337 99895 67340
rect 99837 67331 99895 67337
rect 102778 67328 102784 67340
rect 102836 67328 102842 67380
rect 101766 67300 101772 67312
rect 99668 67272 101772 67300
rect 101766 67260 101772 67272
rect 101824 67260 101830 67312
rect 101950 67260 101956 67312
rect 102008 67260 102014 67312
rect 99469 67235 99527 67241
rect 99469 67201 99481 67235
rect 99515 67201 99527 67235
rect 108301 67235 108359 67241
rect 108301 67232 108313 67235
rect 99469 67195 99527 67201
rect 108132 67204 108313 67232
rect 98641 67167 98699 67173
rect 98641 67133 98653 67167
rect 98687 67164 98699 67167
rect 99558 67164 99564 67176
rect 98687 67136 99564 67164
rect 98687 67133 98699 67136
rect 98641 67127 98699 67133
rect 99558 67124 99564 67136
rect 99616 67124 99622 67176
rect 99377 67099 99435 67105
rect 99377 67065 99389 67099
rect 99423 67096 99435 67099
rect 103054 67096 103060 67108
rect 99423 67068 103060 67096
rect 99423 67065 99435 67068
rect 99377 67059 99435 67065
rect 103054 67056 103060 67068
rect 103112 67056 103118 67108
rect 101858 67028 101864 67040
rect 96908 67000 101864 67028
rect 101858 66988 101864 67000
rect 101916 66988 101922 67040
rect 106182 66988 106188 67040
rect 106240 67028 106246 67040
rect 108132 67037 108160 67204
rect 108301 67201 108313 67204
rect 108347 67201 108359 67235
rect 108301 67195 108359 67201
rect 108117 67031 108175 67037
rect 108117 67028 108129 67031
rect 106240 67000 108129 67028
rect 106240 66988 106246 67000
rect 108117 66997 108129 67000
rect 108163 66997 108175 67031
rect 108117 66991 108175 66997
rect 108482 66988 108488 67040
rect 108540 66988 108546 67040
rect 1104 66938 108836 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 96374 66938
rect 96426 66886 96438 66938
rect 96490 66886 96502 66938
rect 96554 66886 96566 66938
rect 96618 66886 96630 66938
rect 96682 66886 108836 66938
rect 1104 66864 108836 66886
rect 2774 66784 2780 66836
rect 2832 66824 2838 66836
rect 23290 66824 23296 66836
rect 2832 66796 23296 66824
rect 2832 66784 2838 66796
rect 23290 66784 23296 66796
rect 23348 66784 23354 66836
rect 24302 66784 24308 66836
rect 24360 66824 24366 66836
rect 28997 66827 29055 66833
rect 28997 66824 29009 66827
rect 24360 66796 29009 66824
rect 24360 66784 24366 66796
rect 28997 66793 29009 66796
rect 29043 66793 29055 66827
rect 28997 66787 29055 66793
rect 29730 66784 29736 66836
rect 29788 66784 29794 66836
rect 31591 66827 31649 66833
rect 31591 66793 31603 66827
rect 31637 66824 31649 66827
rect 43990 66824 43996 66836
rect 31637 66796 43996 66824
rect 31637 66793 31649 66796
rect 31591 66787 31649 66793
rect 43990 66784 43996 66796
rect 44048 66784 44054 66836
rect 68005 66827 68063 66833
rect 68005 66824 68017 66827
rect 60706 66796 68017 66824
rect 3418 66716 3424 66768
rect 3476 66756 3482 66768
rect 18874 66756 18880 66768
rect 3476 66728 18880 66756
rect 3476 66716 3482 66728
rect 18874 66716 18880 66728
rect 18932 66716 18938 66768
rect 22465 66759 22523 66765
rect 22465 66756 22477 66759
rect 22112 66728 22477 66756
rect 17310 66648 17316 66700
rect 17368 66648 17374 66700
rect 17589 66691 17647 66697
rect 17589 66657 17601 66691
rect 17635 66688 17647 66691
rect 19334 66688 19340 66700
rect 17635 66660 19340 66688
rect 17635 66657 17647 66660
rect 17589 66651 17647 66657
rect 17405 66623 17463 66629
rect 17405 66589 17417 66623
rect 17451 66620 17463 66623
rect 17604 66620 17632 66651
rect 19334 66648 19340 66660
rect 19392 66648 19398 66700
rect 22112 66688 22140 66728
rect 22465 66725 22477 66728
rect 22511 66725 22523 66759
rect 22465 66719 22523 66725
rect 27062 66716 27068 66768
rect 27120 66716 27126 66768
rect 29086 66756 29092 66768
rect 28736 66728 29092 66756
rect 20456 66660 22140 66688
rect 22189 66691 22247 66697
rect 17451 66592 17632 66620
rect 17451 66589 17463 66592
rect 17405 66583 17463 66589
rect 20456 66496 20484 66660
rect 22189 66657 22201 66691
rect 22235 66688 22247 66691
rect 24213 66691 24271 66697
rect 24213 66688 24225 66691
rect 22235 66660 24225 66688
rect 22235 66657 22247 66660
rect 22189 66651 22247 66657
rect 24213 66657 24225 66660
rect 24259 66688 24271 66691
rect 24397 66691 24455 66697
rect 24397 66688 24409 66691
rect 24259 66660 24409 66688
rect 24259 66657 24271 66660
rect 24213 66651 24271 66657
rect 24397 66657 24409 66660
rect 24443 66688 24455 66691
rect 25038 66688 25044 66700
rect 24443 66660 25044 66688
rect 24443 66657 24455 66660
rect 24397 66651 24455 66657
rect 21818 66552 21824 66564
rect 21482 66524 21824 66552
rect 21818 66512 21824 66524
rect 21876 66512 21882 66564
rect 21913 66555 21971 66561
rect 21913 66521 21925 66555
rect 21959 66521 21971 66555
rect 21913 66515 21971 66521
rect 20254 66444 20260 66496
rect 20312 66444 20318 66496
rect 20438 66444 20444 66496
rect 20496 66444 20502 66496
rect 21928 66484 21956 66515
rect 22002 66512 22008 66564
rect 22060 66552 22066 66564
rect 22204 66552 22232 66651
rect 25038 66648 25044 66660
rect 25096 66648 25102 66700
rect 28537 66691 28595 66697
rect 28537 66657 28549 66691
rect 28583 66688 28595 66691
rect 28736 66688 28764 66728
rect 29086 66716 29092 66728
rect 29144 66716 29150 66768
rect 32766 66716 32772 66768
rect 32824 66756 32830 66768
rect 33042 66756 33048 66768
rect 32824 66728 33048 66756
rect 32824 66716 32830 66728
rect 33042 66716 33048 66728
rect 33100 66716 33106 66768
rect 34238 66756 34244 66768
rect 33796 66728 34244 66756
rect 28583 66660 28764 66688
rect 28813 66691 28871 66697
rect 28583 66657 28595 66660
rect 28537 66651 28595 66657
rect 28813 66657 28825 66691
rect 28859 66688 28871 66691
rect 29365 66691 29423 66697
rect 29365 66688 29377 66691
rect 28859 66660 29377 66688
rect 28859 66657 28871 66660
rect 28813 66651 28871 66657
rect 29365 66657 29377 66660
rect 29411 66688 29423 66691
rect 31849 66691 31907 66697
rect 31849 66688 31861 66691
rect 29411 66660 31861 66688
rect 29411 66657 29423 66660
rect 29365 66651 29423 66657
rect 31849 66657 31861 66660
rect 31895 66688 31907 66691
rect 32217 66691 32275 66697
rect 32217 66688 32229 66691
rect 31895 66660 32229 66688
rect 31895 66657 31907 66660
rect 31849 66651 31907 66657
rect 32217 66657 32229 66660
rect 32263 66688 32275 66691
rect 32263 66660 33180 66688
rect 32263 66657 32275 66660
rect 32217 66651 32275 66657
rect 22370 66580 22376 66632
rect 22428 66580 22434 66632
rect 25774 66580 25780 66632
rect 25832 66580 25838 66632
rect 28994 66580 29000 66632
rect 29052 66620 29058 66632
rect 29089 66623 29147 66629
rect 29089 66620 29101 66623
rect 29052 66592 29101 66620
rect 29052 66580 29058 66592
rect 29089 66589 29101 66592
rect 29135 66620 29147 66623
rect 29549 66623 29607 66629
rect 29549 66620 29561 66623
rect 29135 66592 29561 66620
rect 29135 66589 29147 66592
rect 29089 66583 29147 66589
rect 29549 66589 29561 66592
rect 29595 66589 29607 66623
rect 32953 66623 33011 66629
rect 32953 66622 32965 66623
rect 32876 66620 32965 66622
rect 29549 66583 29607 66589
rect 31864 66594 32965 66620
rect 31864 66592 32904 66594
rect 22060 66524 22232 66552
rect 22060 66512 22066 66524
rect 22388 66484 22416 66580
rect 24670 66512 24676 66564
rect 24728 66512 24734 66564
rect 28106 66524 28488 66552
rect 21928 66456 22416 66484
rect 26142 66444 26148 66496
rect 26200 66484 26206 66496
rect 26237 66487 26295 66493
rect 26237 66484 26249 66487
rect 26200 66456 26249 66484
rect 26200 66444 26206 66456
rect 26237 66453 26249 66456
rect 26283 66453 26295 66487
rect 28460 66484 28488 66524
rect 28644 66524 30236 66552
rect 28644 66484 28672 66524
rect 28460 66456 28672 66484
rect 26237 66447 26295 66453
rect 30098 66444 30104 66496
rect 30156 66444 30162 66496
rect 30208 66484 30236 66524
rect 31018 66512 31024 66564
rect 31076 66512 31082 66564
rect 31864 66484 31892 66592
rect 32953 66589 32965 66594
rect 32999 66589 33011 66623
rect 32953 66583 33011 66589
rect 33042 66580 33048 66632
rect 33100 66580 33106 66632
rect 33152 66552 33180 66660
rect 33594 66648 33600 66700
rect 33652 66648 33658 66700
rect 33796 66697 33824 66728
rect 34238 66716 34244 66728
rect 34296 66716 34302 66768
rect 53650 66716 53656 66768
rect 53708 66756 53714 66768
rect 60706 66756 60734 66796
rect 68005 66793 68017 66796
rect 68051 66824 68063 66827
rect 68554 66824 68560 66836
rect 68051 66796 68560 66824
rect 68051 66793 68063 66796
rect 68005 66787 68063 66793
rect 68554 66784 68560 66796
rect 68612 66784 68618 66836
rect 75822 66784 75828 66836
rect 75880 66824 75886 66836
rect 79870 66824 79876 66836
rect 75880 66796 79876 66824
rect 75880 66784 75886 66796
rect 79870 66784 79876 66796
rect 79928 66784 79934 66836
rect 80146 66784 80152 66836
rect 80204 66824 80210 66836
rect 82982 66827 83040 66833
rect 82982 66824 82994 66827
rect 80204 66796 82994 66824
rect 80204 66784 80210 66796
rect 82982 66793 82994 66796
rect 83028 66793 83040 66827
rect 82982 66787 83040 66793
rect 83090 66784 83096 66836
rect 83148 66824 83154 66836
rect 83148 66796 88196 66824
rect 83148 66784 83154 66796
rect 70857 66759 70915 66765
rect 53708 66728 60734 66756
rect 65536 66728 70394 66756
rect 53708 66716 53714 66728
rect 33781 66691 33839 66697
rect 33781 66657 33793 66691
rect 33827 66657 33839 66691
rect 33781 66651 33839 66657
rect 33870 66648 33876 66700
rect 33928 66688 33934 66700
rect 65536 66688 65564 66728
rect 33928 66660 65564 66688
rect 33928 66648 33934 66660
rect 68278 66648 68284 66700
rect 68336 66688 68342 66700
rect 68649 66691 68707 66697
rect 68649 66688 68661 66691
rect 68336 66660 68661 66688
rect 68336 66648 68342 66660
rect 68649 66657 68661 66660
rect 68695 66657 68707 66691
rect 68649 66651 68707 66657
rect 69201 66691 69259 66697
rect 69201 66657 69213 66691
rect 69247 66688 69259 66691
rect 70026 66688 70032 66700
rect 69247 66660 70032 66688
rect 69247 66657 69259 66660
rect 69201 66651 69259 66657
rect 70026 66648 70032 66660
rect 70084 66648 70090 66700
rect 70366 66688 70394 66728
rect 70857 66725 70869 66759
rect 70903 66756 70915 66759
rect 70946 66756 70952 66768
rect 70903 66728 70952 66756
rect 70903 66725 70915 66728
rect 70857 66719 70915 66725
rect 70946 66716 70952 66728
rect 71004 66716 71010 66768
rect 71409 66759 71467 66765
rect 71409 66725 71421 66759
rect 71455 66756 71467 66759
rect 71774 66756 71780 66768
rect 71455 66728 71780 66756
rect 71455 66725 71467 66728
rect 71409 66719 71467 66725
rect 71774 66716 71780 66728
rect 71832 66716 71838 66768
rect 82541 66759 82599 66765
rect 82541 66756 82553 66759
rect 79336 66728 82553 66756
rect 76190 66688 76196 66700
rect 70366 66660 76196 66688
rect 76190 66648 76196 66660
rect 76248 66648 76254 66700
rect 79336 66697 79364 66728
rect 82541 66725 82553 66728
rect 82587 66756 82599 66759
rect 85666 66756 85672 66768
rect 82587 66728 82768 66756
rect 82587 66725 82599 66728
rect 82541 66719 82599 66725
rect 79321 66691 79379 66697
rect 79321 66688 79333 66691
rect 77404 66660 79333 66688
rect 33505 66623 33563 66629
rect 33505 66589 33517 66623
rect 33551 66620 33563 66623
rect 35986 66620 35992 66632
rect 33551 66592 35992 66620
rect 33551 66589 33563 66592
rect 33505 66583 33563 66589
rect 35986 66580 35992 66592
rect 36044 66580 36050 66632
rect 56781 66623 56839 66629
rect 56781 66589 56793 66623
rect 56827 66620 56839 66623
rect 56827 66592 57100 66620
rect 56827 66589 56839 66592
rect 56781 66583 56839 66589
rect 33152 66524 41414 66552
rect 30208 66456 31892 66484
rect 31938 66444 31944 66496
rect 31996 66444 32002 66496
rect 32766 66444 32772 66496
rect 32824 66484 32830 66496
rect 33137 66487 33195 66493
rect 33137 66484 33149 66487
rect 32824 66456 33149 66484
rect 32824 66444 32830 66456
rect 33137 66453 33149 66456
rect 33183 66453 33195 66487
rect 33137 66447 33195 66453
rect 33594 66444 33600 66496
rect 33652 66484 33658 66496
rect 33965 66487 34023 66493
rect 33965 66484 33977 66487
rect 33652 66456 33977 66484
rect 33652 66444 33658 66456
rect 33965 66453 33977 66456
rect 34011 66453 34023 66487
rect 41386 66484 41414 66524
rect 57072 66493 57100 66592
rect 60706 66592 70164 66620
rect 57057 66487 57115 66493
rect 57057 66484 57069 66487
rect 41386 66456 57069 66484
rect 33965 66447 34023 66453
rect 57057 66453 57069 66456
rect 57103 66484 57115 66487
rect 57882 66484 57888 66496
rect 57103 66456 57888 66484
rect 57103 66453 57115 66456
rect 57057 66447 57115 66453
rect 57882 66444 57888 66456
rect 57940 66484 57946 66496
rect 60706 66484 60734 66592
rect 67634 66512 67640 66564
rect 67692 66552 67698 66564
rect 69385 66555 69443 66561
rect 69385 66552 69397 66555
rect 67692 66524 69397 66552
rect 67692 66512 67698 66524
rect 69385 66521 69397 66524
rect 69431 66521 69443 66555
rect 69385 66515 69443 66521
rect 69934 66512 69940 66564
rect 69992 66552 69998 66564
rect 70029 66555 70087 66561
rect 70029 66552 70041 66555
rect 69992 66524 70041 66552
rect 69992 66512 69998 66524
rect 70029 66521 70041 66524
rect 70075 66521 70087 66555
rect 70136 66552 70164 66592
rect 70302 66580 70308 66632
rect 70360 66580 70366 66632
rect 70578 66580 70584 66632
rect 70636 66620 70642 66632
rect 75914 66620 75920 66632
rect 70636 66592 75920 66620
rect 70636 66580 70642 66592
rect 75914 66580 75920 66592
rect 75972 66580 75978 66632
rect 77404 66561 77432 66660
rect 79321 66657 79333 66660
rect 79367 66657 79379 66691
rect 79321 66651 79379 66657
rect 79413 66691 79471 66697
rect 79413 66657 79425 66691
rect 79459 66657 79471 66691
rect 79413 66651 79471 66657
rect 79873 66691 79931 66697
rect 79873 66657 79885 66691
rect 79919 66688 79931 66691
rect 79962 66688 79968 66700
rect 79919 66660 79968 66688
rect 79919 66657 79931 66660
rect 79873 66651 79931 66657
rect 77938 66580 77944 66632
rect 77996 66580 78002 66632
rect 77389 66555 77447 66561
rect 77389 66552 77401 66555
rect 70136 66524 77401 66552
rect 70029 66515 70087 66521
rect 77389 66521 77401 66524
rect 77435 66521 77447 66555
rect 77389 66515 77447 66521
rect 79045 66555 79103 66561
rect 79045 66521 79057 66555
rect 79091 66552 79103 66555
rect 79428 66552 79456 66651
rect 79962 66648 79968 66660
rect 80020 66648 80026 66700
rect 82740 66697 82768 66728
rect 84120 66728 85672 66756
rect 82725 66691 82783 66697
rect 82725 66657 82737 66691
rect 82771 66688 82783 66691
rect 83366 66688 83372 66700
rect 82771 66660 83372 66688
rect 82771 66657 82783 66660
rect 82725 66651 82783 66657
rect 83366 66648 83372 66660
rect 83424 66648 83430 66700
rect 79778 66580 79784 66632
rect 79836 66620 79842 66632
rect 79836 66592 82676 66620
rect 84120 66606 84148 66728
rect 85666 66716 85672 66728
rect 85724 66716 85730 66768
rect 84473 66691 84531 66697
rect 84473 66657 84485 66691
rect 84519 66657 84531 66691
rect 84473 66651 84531 66657
rect 84488 66620 84516 66651
rect 84838 66648 84844 66700
rect 84896 66648 84902 66700
rect 85209 66691 85267 66697
rect 85209 66657 85221 66691
rect 85255 66657 85267 66691
rect 85209 66651 85267 66657
rect 84654 66620 84660 66632
rect 84488 66592 84660 66620
rect 79836 66580 79842 66592
rect 79091 66524 79456 66552
rect 79091 66521 79103 66524
rect 79045 66515 79103 66521
rect 57940 66456 60734 66484
rect 68925 66487 68983 66493
rect 57940 66444 57946 66456
rect 68925 66453 68937 66487
rect 68971 66484 68983 66487
rect 69290 66484 69296 66496
rect 68971 66456 69296 66484
rect 68971 66453 68983 66456
rect 68925 66447 68983 66453
rect 69290 66444 69296 66456
rect 69348 66444 69354 66496
rect 69753 66487 69811 66493
rect 69753 66453 69765 66487
rect 69799 66484 69811 66487
rect 69842 66484 69848 66496
rect 69799 66456 69848 66484
rect 69799 66453 69811 66456
rect 69753 66447 69811 66453
rect 69842 66444 69848 66456
rect 69900 66444 69906 66496
rect 70044 66484 70072 66515
rect 70397 66487 70455 66493
rect 70397 66484 70409 66487
rect 70044 66456 70409 66484
rect 70397 66453 70409 66456
rect 70443 66453 70455 66487
rect 70397 66447 70455 66453
rect 77570 66444 77576 66496
rect 77628 66444 77634 66496
rect 80146 66444 80152 66496
rect 80204 66444 80210 66496
rect 82648 66484 82676 66592
rect 84654 66580 84660 66592
rect 84712 66580 84718 66632
rect 85224 66552 85252 66651
rect 85390 66648 85396 66700
rect 85448 66648 85454 66700
rect 86218 66648 86224 66700
rect 86276 66688 86282 66700
rect 88168 66688 88196 66796
rect 88334 66784 88340 66836
rect 88392 66824 88398 66836
rect 91630 66827 91688 66833
rect 91630 66824 91642 66827
rect 88392 66796 91642 66824
rect 88392 66784 88398 66796
rect 91630 66793 91642 66796
rect 91676 66793 91688 66827
rect 91630 66787 91688 66793
rect 92014 66784 92020 66836
rect 92072 66824 92078 66836
rect 94498 66824 94504 66836
rect 92072 66796 94504 66824
rect 92072 66784 92078 66796
rect 94498 66784 94504 66796
rect 94556 66784 94562 66836
rect 94958 66784 94964 66836
rect 95016 66784 95022 66836
rect 96154 66784 96160 66836
rect 96212 66784 96218 66836
rect 96246 66784 96252 66836
rect 96304 66824 96310 66836
rect 96985 66827 97043 66833
rect 96985 66824 96997 66827
rect 96304 66796 96997 66824
rect 96304 66784 96310 66796
rect 96985 66793 96997 66796
rect 97031 66824 97043 66827
rect 99374 66824 99380 66836
rect 97031 66796 99380 66824
rect 97031 66793 97043 66796
rect 96985 66787 97043 66793
rect 99374 66784 99380 66796
rect 99432 66784 99438 66836
rect 99466 66784 99472 66836
rect 99524 66824 99530 66836
rect 99561 66827 99619 66833
rect 99561 66824 99573 66827
rect 99524 66796 99573 66824
rect 99524 66784 99530 66796
rect 99561 66793 99573 66796
rect 99607 66824 99619 66827
rect 104250 66824 104256 66836
rect 99607 66796 104256 66824
rect 99607 66793 99619 66796
rect 99561 66787 99619 66793
rect 104250 66784 104256 66796
rect 104308 66784 104314 66836
rect 93121 66759 93179 66765
rect 93121 66725 93133 66759
rect 93167 66756 93179 66759
rect 93167 66728 93348 66756
rect 93167 66725 93179 66728
rect 93121 66719 93179 66725
rect 88324 66691 88382 66697
rect 88324 66688 88336 66691
rect 86276 66660 87828 66688
rect 88168 66660 88336 66688
rect 86276 66648 86282 66660
rect 87800 66620 87828 66660
rect 88324 66657 88336 66660
rect 88370 66657 88382 66691
rect 88324 66651 88382 66657
rect 88426 66648 88432 66700
rect 88484 66688 88490 66700
rect 90913 66691 90971 66697
rect 90913 66688 90925 66691
rect 88484 66660 90925 66688
rect 88484 66648 88490 66660
rect 90913 66657 90925 66660
rect 90959 66688 90971 66691
rect 91373 66691 91431 66697
rect 91373 66688 91385 66691
rect 90959 66660 91385 66688
rect 90959 66657 90971 66660
rect 90913 66651 90971 66657
rect 91373 66657 91385 66660
rect 91419 66688 91431 66691
rect 93320 66688 93348 66728
rect 96062 66716 96068 66768
rect 96120 66756 96126 66768
rect 96430 66756 96436 66768
rect 96120 66728 96436 66756
rect 96120 66716 96126 66728
rect 96430 66716 96436 66728
rect 96488 66716 96494 66768
rect 96706 66716 96712 66768
rect 96764 66756 96770 66768
rect 104618 66756 104624 66768
rect 96764 66728 104624 66756
rect 96764 66716 96770 66728
rect 104618 66716 104624 66728
rect 104676 66716 104682 66768
rect 94038 66688 94044 66700
rect 91419 66660 93256 66688
rect 93320 66660 94044 66688
rect 91419 66657 91431 66660
rect 91373 66651 91431 66657
rect 93228 66632 93256 66660
rect 94038 66648 94044 66660
rect 94096 66648 94102 66700
rect 95329 66691 95387 66697
rect 95329 66657 95341 66691
rect 95375 66688 95387 66691
rect 95973 66691 96031 66697
rect 95973 66688 95985 66691
rect 95375 66660 95985 66688
rect 95375 66657 95387 66660
rect 95329 66651 95387 66657
rect 95973 66657 95985 66660
rect 96019 66688 96031 66691
rect 96019 66660 101720 66688
rect 96019 66657 96031 66660
rect 95973 66651 96031 66657
rect 88061 66623 88119 66629
rect 88061 66620 88073 66623
rect 87800 66592 88073 66620
rect 88061 66589 88073 66592
rect 88107 66589 88119 66623
rect 88061 66583 88119 66589
rect 89622 66580 89628 66632
rect 89680 66620 89686 66632
rect 90085 66623 90143 66629
rect 90085 66620 90097 66623
rect 89680 66592 90097 66620
rect 89680 66580 89686 66592
rect 90085 66589 90097 66592
rect 90131 66620 90143 66623
rect 90177 66623 90235 66629
rect 90177 66620 90189 66623
rect 90131 66592 90189 66620
rect 90131 66589 90143 66592
rect 90085 66583 90143 66589
rect 90177 66589 90189 66592
rect 90223 66589 90235 66623
rect 90177 66583 90235 66589
rect 93210 66580 93216 66632
rect 93268 66580 93274 66632
rect 95513 66623 95571 66629
rect 95513 66620 95525 66623
rect 94792 66592 95525 66620
rect 84304 66524 85252 66552
rect 84304 66484 84332 66524
rect 85298 66512 85304 66564
rect 85356 66552 85362 66564
rect 86497 66555 86555 66561
rect 86497 66552 86509 66555
rect 85356 66524 86509 66552
rect 85356 66512 85362 66524
rect 86497 66521 86509 66524
rect 86543 66521 86555 66555
rect 87722 66524 88288 66552
rect 86497 66515 86555 66521
rect 82648 66456 84332 66484
rect 84930 66444 84936 66496
rect 84988 66484 84994 66496
rect 85485 66487 85543 66493
rect 85485 66484 85497 66487
rect 84988 66456 85497 66484
rect 84988 66444 84994 66456
rect 85485 66453 85497 66456
rect 85531 66453 85543 66487
rect 85485 66447 85543 66453
rect 85853 66487 85911 66493
rect 85853 66453 85865 66487
rect 85899 66484 85911 66487
rect 87874 66484 87880 66496
rect 85899 66456 87880 66484
rect 85899 66453 85911 66456
rect 85853 66447 85911 66453
rect 87874 66444 87880 66456
rect 87932 66444 87938 66496
rect 87966 66444 87972 66496
rect 88024 66444 88030 66496
rect 88260 66484 88288 66524
rect 88334 66512 88340 66564
rect 88392 66552 88398 66564
rect 89993 66555 90051 66561
rect 89993 66552 90005 66555
rect 88392 66524 88826 66552
rect 89686 66524 90005 66552
rect 88392 66512 88398 66524
rect 89686 66484 89714 66524
rect 89993 66521 90005 66524
rect 90039 66521 90051 66555
rect 90545 66555 90603 66561
rect 90545 66552 90557 66555
rect 89993 66515 90051 66521
rect 90192 66524 90557 66552
rect 88260 66456 89714 66484
rect 89809 66487 89867 66493
rect 89809 66453 89821 66487
rect 89855 66484 89867 66487
rect 90192 66484 90220 66524
rect 90545 66521 90557 66524
rect 90591 66552 90603 66555
rect 90591 66524 92060 66552
rect 92874 66524 93440 66552
rect 90591 66521 90603 66524
rect 90545 66515 90603 66521
rect 89855 66456 90220 66484
rect 89855 66453 89867 66456
rect 89809 66447 89867 66453
rect 90266 66444 90272 66496
rect 90324 66444 90330 66496
rect 90729 66487 90787 66493
rect 90729 66453 90741 66487
rect 90775 66484 90787 66487
rect 90910 66484 90916 66496
rect 90775 66456 90916 66484
rect 90775 66453 90787 66456
rect 90729 66447 90787 66453
rect 90910 66444 90916 66456
rect 90968 66444 90974 66496
rect 92032 66484 92060 66524
rect 93026 66484 93032 66496
rect 92032 66456 93032 66484
rect 93026 66444 93032 66456
rect 93084 66444 93090 66496
rect 93412 66484 93440 66524
rect 93486 66512 93492 66564
rect 93544 66512 93550 66564
rect 93578 66512 93584 66564
rect 93636 66552 93642 66564
rect 93636 66524 93978 66552
rect 93636 66512 93642 66524
rect 94792 66484 94820 66592
rect 95513 66589 95525 66592
rect 95559 66589 95571 66623
rect 95513 66583 95571 66589
rect 95605 66623 95663 66629
rect 95605 66589 95617 66623
rect 95651 66620 95663 66623
rect 96154 66620 96160 66632
rect 95651 66592 96160 66620
rect 95651 66589 95663 66592
rect 95605 66583 95663 66589
rect 94958 66512 94964 66564
rect 95016 66552 95022 66564
rect 95145 66555 95203 66561
rect 95145 66552 95157 66555
rect 95016 66524 95157 66552
rect 95016 66512 95022 66524
rect 95145 66521 95157 66524
rect 95191 66521 95203 66555
rect 95145 66515 95203 66521
rect 93412 66456 94820 66484
rect 94866 66444 94872 66496
rect 94924 66484 94930 66496
rect 95620 66484 95648 66583
rect 96154 66580 96160 66592
rect 96212 66580 96218 66632
rect 96614 66580 96620 66632
rect 96672 66620 96678 66632
rect 96801 66623 96859 66629
rect 96801 66620 96813 66623
rect 96672 66592 96813 66620
rect 96672 66580 96678 66592
rect 96801 66589 96813 66592
rect 96847 66620 96859 66623
rect 98181 66623 98239 66629
rect 98181 66620 98193 66623
rect 96847 66592 98193 66620
rect 96847 66589 96859 66592
rect 96801 66583 96859 66589
rect 98181 66589 98193 66592
rect 98227 66620 98239 66623
rect 98362 66620 98368 66632
rect 98227 66592 98368 66620
rect 98227 66589 98239 66592
rect 98181 66583 98239 66589
rect 98362 66580 98368 66592
rect 98420 66580 98426 66632
rect 98457 66623 98515 66629
rect 98457 66589 98469 66623
rect 98503 66620 98515 66623
rect 99466 66620 99472 66632
rect 98503 66592 99472 66620
rect 98503 66589 98515 66592
rect 98457 66583 98515 66589
rect 99466 66580 99472 66592
rect 99524 66580 99530 66632
rect 95694 66512 95700 66564
rect 95752 66552 95758 66564
rect 98270 66552 98276 66564
rect 95752 66524 98276 66552
rect 95752 66512 95758 66524
rect 98270 66512 98276 66524
rect 98328 66552 98334 66564
rect 99193 66555 99251 66561
rect 99193 66552 99205 66555
rect 98328 66524 99205 66552
rect 98328 66512 98334 66524
rect 99193 66521 99205 66524
rect 99239 66521 99251 66555
rect 99193 66515 99251 66521
rect 99377 66555 99435 66561
rect 99377 66521 99389 66555
rect 99423 66552 99435 66555
rect 99423 66524 99788 66552
rect 99423 66521 99435 66524
rect 99377 66515 99435 66521
rect 99760 66496 99788 66524
rect 94924 66456 95648 66484
rect 94924 66444 94930 66456
rect 95786 66444 95792 66496
rect 95844 66484 95850 66496
rect 96154 66484 96160 66496
rect 95844 66456 96160 66484
rect 95844 66444 95850 66456
rect 96154 66444 96160 66456
rect 96212 66484 96218 66496
rect 96249 66487 96307 66493
rect 96249 66484 96261 66487
rect 96212 66456 96261 66484
rect 96212 66444 96218 66456
rect 96249 66453 96261 66456
rect 96295 66453 96307 66487
rect 96249 66447 96307 66453
rect 96617 66487 96675 66493
rect 96617 66453 96629 66487
rect 96663 66484 96675 66487
rect 96890 66484 96896 66496
rect 96663 66456 96896 66484
rect 96663 66453 96675 66456
rect 96617 66447 96675 66453
rect 96890 66444 96896 66456
rect 96948 66444 96954 66496
rect 99742 66444 99748 66496
rect 99800 66444 99806 66496
rect 101692 66484 101720 66660
rect 101784 66660 102272 66688
rect 101784 66632 101812 66660
rect 101766 66580 101772 66632
rect 101824 66580 101830 66632
rect 101858 66580 101864 66632
rect 101916 66620 101922 66632
rect 102045 66623 102103 66629
rect 102045 66620 102057 66623
rect 101916 66592 102057 66620
rect 101916 66580 101922 66592
rect 102045 66589 102057 66592
rect 102091 66589 102103 66623
rect 102045 66583 102103 66589
rect 102134 66580 102140 66632
rect 102192 66580 102198 66632
rect 102244 66629 102272 66660
rect 102229 66623 102287 66629
rect 102229 66589 102241 66623
rect 102275 66589 102287 66623
rect 102229 66583 102287 66589
rect 101950 66512 101956 66564
rect 102008 66552 102014 66564
rect 102321 66555 102379 66561
rect 102321 66552 102333 66555
rect 102008 66524 102333 66552
rect 102008 66512 102014 66524
rect 102321 66521 102333 66524
rect 102367 66521 102379 66555
rect 102321 66515 102379 66521
rect 104802 66484 104808 66496
rect 101692 66456 104808 66484
rect 104802 66444 104808 66456
rect 104860 66444 104866 66496
rect 1104 66394 108836 66416
rect 1104 66342 4874 66394
rect 4926 66342 4938 66394
rect 4990 66342 5002 66394
rect 5054 66342 5066 66394
rect 5118 66342 5130 66394
rect 5182 66342 35594 66394
rect 35646 66342 35658 66394
rect 35710 66342 35722 66394
rect 35774 66342 35786 66394
rect 35838 66342 35850 66394
rect 35902 66342 66314 66394
rect 66366 66342 66378 66394
rect 66430 66342 66442 66394
rect 66494 66342 66506 66394
rect 66558 66342 66570 66394
rect 66622 66342 97034 66394
rect 97086 66342 97098 66394
rect 97150 66342 97162 66394
rect 97214 66342 97226 66394
rect 97278 66342 97290 66394
rect 97342 66342 106658 66394
rect 106710 66342 106722 66394
rect 106774 66342 106786 66394
rect 106838 66342 106850 66394
rect 106902 66342 106914 66394
rect 106966 66342 108836 66394
rect 1104 66320 108836 66342
rect 9582 66240 9588 66292
rect 9640 66280 9646 66292
rect 16390 66280 16396 66292
rect 9640 66252 16396 66280
rect 9640 66240 9646 66252
rect 16390 66240 16396 66252
rect 16448 66240 16454 66292
rect 20438 66280 20444 66292
rect 16500 66252 20444 66280
rect 16500 66212 16528 66252
rect 20438 66240 20444 66252
rect 20496 66240 20502 66292
rect 21913 66283 21971 66289
rect 21913 66249 21925 66283
rect 21959 66280 21971 66283
rect 28905 66283 28963 66289
rect 21959 66252 22140 66280
rect 21959 66249 21971 66252
rect 21913 66243 21971 66249
rect 21361 66215 21419 66221
rect 21361 66212 21373 66215
rect 6886 66184 16528 66212
rect 20272 66184 21373 66212
rect 1581 66147 1639 66153
rect 1581 66113 1593 66147
rect 1627 66144 1639 66147
rect 1765 66147 1823 66153
rect 1765 66144 1777 66147
rect 1627 66116 1777 66144
rect 1627 66113 1639 66116
rect 1581 66107 1639 66113
rect 1765 66113 1777 66116
rect 1811 66144 1823 66147
rect 6886 66144 6914 66184
rect 20272 66156 20300 66184
rect 21361 66181 21373 66184
rect 21407 66212 21419 66215
rect 21545 66215 21603 66221
rect 21545 66212 21557 66215
rect 21407 66184 21557 66212
rect 21407 66181 21419 66184
rect 21361 66175 21419 66181
rect 21545 66181 21557 66184
rect 21591 66212 21603 66215
rect 22002 66212 22008 66224
rect 21591 66184 22008 66212
rect 21591 66181 21603 66184
rect 21545 66175 21603 66181
rect 22002 66172 22008 66184
rect 22060 66172 22066 66224
rect 22112 66212 22140 66252
rect 22664 66252 23704 66280
rect 22281 66215 22339 66221
rect 22281 66212 22293 66215
rect 22112 66184 22293 66212
rect 22281 66181 22293 66184
rect 22327 66212 22339 66215
rect 22664 66212 22692 66252
rect 22327 66184 22692 66212
rect 22327 66181 22339 66184
rect 22281 66175 22339 66181
rect 1811 66116 6914 66144
rect 1811 66113 1823 66116
rect 1765 66107 1823 66113
rect 16574 66104 16580 66156
rect 16632 66144 16638 66156
rect 17865 66147 17923 66153
rect 17865 66144 17877 66147
rect 16632 66116 17877 66144
rect 16632 66104 16638 66116
rect 17865 66113 17877 66116
rect 17911 66144 17923 66147
rect 19337 66147 19395 66153
rect 19337 66144 19349 66147
rect 17911 66116 19349 66144
rect 17911 66113 17923 66116
rect 17865 66107 17923 66113
rect 19337 66113 19349 66116
rect 19383 66144 19395 66147
rect 19429 66147 19487 66153
rect 19429 66144 19441 66147
rect 19383 66116 19441 66144
rect 19383 66113 19395 66116
rect 19337 66107 19395 66113
rect 19429 66113 19441 66116
rect 19475 66144 19487 66147
rect 20254 66144 20260 66156
rect 19475 66116 20260 66144
rect 19475 66113 19487 66116
rect 19429 66107 19487 66113
rect 20254 66104 20260 66116
rect 20312 66104 20318 66156
rect 21177 66147 21235 66153
rect 21177 66113 21189 66147
rect 21223 66144 21235 66147
rect 21266 66144 21272 66156
rect 21223 66116 21272 66144
rect 21223 66113 21235 66116
rect 21177 66107 21235 66113
rect 21266 66104 21272 66116
rect 21324 66144 21330 66156
rect 21324 66116 21956 66144
rect 21324 66104 21330 66116
rect 842 65900 848 65952
rect 900 65940 906 65952
rect 1397 65943 1455 65949
rect 1397 65940 1409 65943
rect 900 65912 1409 65940
rect 900 65900 906 65912
rect 1397 65909 1409 65912
rect 1443 65909 1455 65943
rect 21928 65940 21956 66116
rect 22020 66085 22048 66172
rect 23566 66144 23572 66156
rect 23414 66116 23572 66144
rect 23566 66104 23572 66116
rect 23624 66104 23630 66156
rect 23676 66144 23704 66252
rect 28905 66249 28917 66283
rect 28951 66280 28963 66283
rect 29086 66280 29092 66292
rect 28951 66252 29092 66280
rect 28951 66249 28963 66252
rect 28905 66243 28963 66249
rect 29086 66240 29092 66252
rect 29144 66240 29150 66292
rect 30098 66240 30104 66292
rect 30156 66280 30162 66292
rect 31938 66280 31944 66292
rect 30156 66252 31944 66280
rect 30156 66240 30162 66252
rect 31938 66240 31944 66252
rect 31996 66240 32002 66292
rect 32950 66240 32956 66292
rect 33008 66280 33014 66292
rect 39390 66280 39396 66292
rect 33008 66252 39396 66280
rect 33008 66240 33014 66252
rect 39390 66240 39396 66252
rect 39448 66240 39454 66292
rect 70302 66240 70308 66292
rect 70360 66280 70366 66292
rect 77570 66280 77576 66292
rect 70360 66252 77576 66280
rect 70360 66240 70366 66252
rect 77570 66240 77576 66252
rect 77628 66240 77634 66292
rect 80146 66240 80152 66292
rect 80204 66280 80210 66292
rect 86954 66280 86960 66292
rect 80204 66252 86960 66280
rect 80204 66240 80210 66252
rect 86954 66240 86960 66252
rect 87012 66240 87018 66292
rect 88334 66280 88340 66292
rect 87340 66252 88340 66280
rect 23750 66172 23756 66224
rect 23808 66212 23814 66224
rect 30558 66212 30564 66224
rect 23808 66184 30564 66212
rect 23808 66172 23814 66184
rect 30558 66172 30564 66184
rect 30616 66172 30622 66224
rect 31018 66172 31024 66224
rect 31076 66172 31082 66224
rect 31202 66212 31208 66224
rect 31128 66184 31208 66212
rect 31128 66153 31156 66184
rect 31202 66172 31208 66184
rect 31260 66172 31266 66224
rect 57701 66215 57759 66221
rect 57701 66181 57713 66215
rect 57747 66212 57759 66215
rect 57882 66212 57888 66224
rect 57747 66184 57888 66212
rect 57747 66181 57759 66184
rect 57701 66175 57759 66181
rect 57882 66172 57888 66184
rect 57940 66212 57946 66224
rect 58069 66215 58127 66221
rect 58069 66212 58081 66215
rect 57940 66184 58081 66212
rect 57940 66172 57946 66184
rect 58069 66181 58081 66184
rect 58115 66181 58127 66215
rect 58069 66175 58127 66181
rect 83366 66172 83372 66224
rect 83424 66172 83430 66224
rect 86313 66215 86371 66221
rect 86313 66181 86325 66215
rect 86359 66212 86371 66215
rect 87340 66212 87368 66252
rect 88334 66240 88340 66252
rect 88392 66240 88398 66292
rect 88426 66240 88432 66292
rect 88484 66280 88490 66292
rect 88521 66283 88579 66289
rect 88521 66280 88533 66283
rect 88484 66252 88533 66280
rect 88484 66240 88490 66252
rect 88521 66249 88533 66252
rect 88567 66249 88579 66283
rect 88521 66243 88579 66249
rect 86359 66184 87368 66212
rect 88536 66212 88564 66243
rect 89622 66240 89628 66292
rect 89680 66240 89686 66292
rect 92109 66283 92167 66289
rect 92109 66249 92121 66283
rect 92155 66280 92167 66283
rect 93302 66280 93308 66292
rect 92155 66252 93308 66280
rect 92155 66249 92167 66252
rect 92109 66243 92167 66249
rect 93302 66240 93308 66252
rect 93360 66240 93366 66292
rect 96706 66280 96712 66292
rect 93412 66252 96712 66280
rect 89640 66212 89668 66240
rect 89717 66215 89775 66221
rect 89717 66212 89729 66215
rect 88536 66184 89484 66212
rect 89640 66184 89729 66212
rect 86359 66181 86371 66184
rect 86313 66175 86371 66181
rect 31113 66147 31171 66153
rect 23676 66116 25360 66144
rect 22005 66079 22063 66085
rect 22005 66045 22017 66079
rect 22051 66045 22063 66079
rect 22005 66039 22063 66045
rect 22370 66036 22376 66088
rect 22428 66076 22434 66088
rect 23753 66079 23811 66085
rect 23753 66076 23765 66079
rect 22428 66048 23765 66076
rect 22428 66036 22434 66048
rect 23753 66045 23765 66048
rect 23799 66076 23811 66079
rect 23845 66079 23903 66085
rect 23845 66076 23857 66079
rect 23799 66048 23857 66076
rect 23799 66045 23811 66048
rect 23753 66039 23811 66045
rect 23845 66045 23857 66048
rect 23891 66045 23903 66079
rect 25332 66076 25360 66116
rect 31113 66113 31125 66147
rect 31159 66113 31171 66147
rect 55953 66147 56011 66153
rect 55953 66144 55965 66147
rect 31113 66107 31171 66113
rect 41386 66116 55965 66144
rect 32766 66076 32772 66088
rect 25332 66048 32772 66076
rect 23845 66039 23903 66045
rect 32766 66036 32772 66048
rect 32824 66036 32830 66088
rect 41386 66008 41414 66116
rect 55953 66113 55965 66116
rect 55999 66144 56011 66147
rect 57977 66147 58035 66153
rect 57977 66144 57989 66147
rect 55999 66116 57989 66144
rect 55999 66113 56011 66116
rect 55953 66107 56011 66113
rect 57977 66113 57989 66116
rect 58023 66144 58035 66147
rect 60734 66144 60740 66156
rect 58023 66116 60740 66144
rect 58023 66113 58035 66116
rect 57977 66107 58035 66113
rect 60734 66104 60740 66116
rect 60792 66104 60798 66156
rect 83384 66144 83412 66172
rect 83645 66147 83703 66153
rect 83645 66144 83657 66147
rect 83384 66116 83657 66144
rect 83645 66113 83657 66116
rect 83691 66113 83703 66147
rect 86405 66147 86463 66153
rect 83645 66107 83703 66113
rect 73982 66036 73988 66088
rect 74040 66076 74046 66088
rect 83921 66079 83979 66085
rect 83921 66076 83933 66079
rect 74040 66048 83933 66076
rect 74040 66036 74046 66048
rect 83921 66045 83933 66048
rect 83967 66045 83979 66079
rect 83921 66039 83979 66045
rect 23676 65980 41414 66008
rect 85040 66008 85068 66130
rect 86405 66113 86417 66147
rect 86451 66144 86463 66147
rect 86494 66144 86500 66156
rect 86451 66116 86500 66144
rect 86451 66113 86463 66116
rect 86405 66107 86463 66113
rect 86494 66104 86500 66116
rect 86552 66104 86558 66156
rect 86681 66147 86739 66153
rect 86681 66144 86693 66147
rect 86604 66116 86693 66144
rect 86218 66036 86224 66088
rect 86276 66076 86282 66088
rect 86604 66076 86632 66116
rect 86681 66113 86693 66116
rect 86727 66113 86739 66147
rect 86681 66107 86739 66113
rect 88058 66104 88064 66156
rect 88116 66104 88122 66156
rect 88426 66104 88432 66156
rect 88484 66144 88490 66156
rect 88610 66144 88616 66156
rect 88484 66116 88616 66144
rect 88484 66104 88490 66116
rect 88610 66104 88616 66116
rect 88668 66104 88674 66156
rect 89070 66104 89076 66156
rect 89128 66104 89134 66156
rect 89456 66153 89484 66184
rect 89717 66181 89729 66184
rect 89763 66181 89775 66215
rect 89717 66175 89775 66181
rect 89806 66172 89812 66224
rect 89864 66212 89870 66224
rect 92385 66215 92443 66221
rect 89864 66184 90206 66212
rect 89864 66172 89870 66184
rect 92385 66181 92397 66215
rect 92431 66212 92443 66215
rect 92934 66212 92940 66224
rect 92431 66184 92940 66212
rect 92431 66181 92443 66184
rect 92385 66175 92443 66181
rect 92934 66172 92940 66184
rect 92992 66172 92998 66224
rect 93026 66172 93032 66224
rect 93084 66212 93090 66224
rect 93412 66212 93440 66252
rect 96706 66240 96712 66252
rect 96764 66240 96770 66292
rect 98270 66240 98276 66292
rect 98328 66240 98334 66292
rect 98549 66283 98607 66289
rect 98549 66249 98561 66283
rect 98595 66280 98607 66283
rect 99190 66280 99196 66292
rect 98595 66252 99196 66280
rect 98595 66249 98607 66252
rect 98549 66243 98607 66249
rect 93084 66184 93440 66212
rect 94041 66215 94099 66221
rect 93084 66172 93090 66184
rect 94041 66181 94053 66215
rect 94087 66212 94099 66215
rect 94087 66184 94898 66212
rect 94087 66181 94099 66184
rect 94041 66175 94099 66181
rect 96062 66172 96068 66224
rect 96120 66172 96126 66224
rect 96430 66172 96436 66224
rect 96488 66212 96494 66224
rect 96488 66184 97290 66212
rect 96488 66172 96494 66184
rect 98362 66172 98368 66224
rect 98420 66172 98426 66224
rect 89349 66147 89407 66153
rect 89349 66113 89361 66147
rect 89395 66113 89407 66147
rect 89349 66107 89407 66113
rect 89441 66147 89499 66153
rect 89441 66113 89453 66147
rect 89487 66113 89499 66147
rect 89441 66107 89499 66113
rect 91557 66147 91615 66153
rect 91557 66113 91569 66147
rect 91603 66144 91615 66147
rect 92658 66144 92664 66156
rect 91603 66116 92664 66144
rect 91603 66113 91615 66116
rect 91557 66107 91615 66113
rect 86957 66079 87015 66085
rect 86957 66076 86969 66079
rect 86276 66048 86632 66076
rect 86788 66048 86969 66076
rect 86276 66036 86282 66048
rect 86586 66008 86592 66020
rect 85040 65980 86592 66008
rect 23676 65940 23704 65980
rect 86586 65968 86592 65980
rect 86644 65968 86650 66020
rect 86788 66008 86816 66048
rect 86957 66045 86969 66048
rect 87003 66045 87015 66079
rect 89364 66076 89392 66107
rect 92658 66104 92664 66116
rect 92716 66104 92722 66156
rect 92768 66116 93900 66144
rect 90910 66076 90916 66088
rect 89364 66048 90916 66076
rect 86957 66039 87015 66045
rect 90910 66036 90916 66048
rect 90968 66036 90974 66088
rect 91649 66079 91707 66085
rect 91649 66045 91661 66079
rect 91695 66045 91707 66079
rect 91649 66039 91707 66045
rect 91925 66079 91983 66085
rect 91925 66045 91937 66079
rect 91971 66076 91983 66079
rect 92290 66076 92296 66088
rect 91971 66048 92296 66076
rect 91971 66045 91983 66048
rect 91925 66039 91983 66045
rect 91664 66008 91692 66039
rect 92290 66036 92296 66048
rect 92348 66036 92354 66088
rect 92768 66076 92796 66116
rect 92676 66048 92796 66076
rect 92845 66079 92903 66085
rect 92201 66011 92259 66017
rect 92201 66008 92213 66011
rect 86696 65980 86816 66008
rect 88352 65980 88564 66008
rect 91664 65980 92213 66008
rect 21928 65912 23704 65940
rect 1397 65903 1455 65909
rect 53650 65900 53656 65952
rect 53708 65900 53714 65952
rect 85393 65943 85451 65949
rect 85393 65909 85405 65943
rect 85439 65940 85451 65943
rect 85574 65940 85580 65952
rect 85439 65912 85580 65940
rect 85439 65909 85451 65912
rect 85393 65903 85451 65909
rect 85574 65900 85580 65912
rect 85632 65900 85638 65952
rect 86494 65900 86500 65952
rect 86552 65940 86558 65952
rect 86696 65940 86724 65980
rect 86552 65912 86724 65940
rect 86552 65900 86558 65912
rect 86770 65900 86776 65952
rect 86828 65940 86834 65952
rect 88352 65940 88380 65980
rect 86828 65912 88380 65940
rect 86828 65900 86834 65912
rect 88426 65900 88432 65952
rect 88484 65900 88490 65952
rect 88536 65940 88564 65980
rect 92201 65977 92213 65980
rect 92247 66008 92259 66011
rect 92676 66008 92704 66048
rect 92845 66045 92857 66079
rect 92891 66076 92903 66079
rect 93486 66076 93492 66088
rect 92891 66048 93492 66076
rect 92891 66045 92903 66048
rect 92845 66039 92903 66045
rect 93486 66036 93492 66048
rect 93544 66036 93550 66088
rect 93872 66076 93900 66116
rect 93946 66104 93952 66156
rect 94004 66104 94010 66156
rect 94317 66147 94375 66153
rect 94317 66113 94329 66147
rect 94363 66144 94375 66147
rect 94498 66144 94504 66156
rect 94363 66116 94504 66144
rect 94363 66113 94375 66116
rect 94317 66107 94375 66113
rect 94498 66104 94504 66116
rect 94556 66104 94562 66156
rect 96338 66104 96344 66156
rect 96396 66144 96402 66156
rect 99116 66153 99144 66252
rect 99190 66240 99196 66252
rect 99248 66240 99254 66292
rect 99374 66240 99380 66292
rect 99432 66280 99438 66292
rect 100021 66283 100079 66289
rect 100021 66280 100033 66283
rect 99432 66252 100033 66280
rect 99432 66240 99438 66252
rect 100021 66249 100033 66252
rect 100067 66249 100079 66283
rect 100021 66243 100079 66249
rect 99742 66172 99748 66224
rect 99800 66212 99806 66224
rect 102134 66212 102140 66224
rect 99800 66184 102140 66212
rect 99800 66172 99806 66184
rect 102134 66172 102140 66184
rect 102192 66172 102198 66224
rect 96525 66147 96583 66153
rect 96525 66144 96537 66147
rect 96396 66116 96537 66144
rect 96396 66104 96402 66116
rect 96525 66113 96537 66116
rect 96571 66113 96583 66147
rect 96525 66107 96583 66113
rect 98641 66147 98699 66153
rect 98641 66113 98653 66147
rect 98687 66144 98699 66147
rect 98733 66147 98791 66153
rect 98733 66144 98745 66147
rect 98687 66116 98745 66144
rect 98687 66113 98699 66116
rect 98641 66107 98699 66113
rect 98733 66113 98745 66116
rect 98779 66113 98791 66147
rect 98733 66107 98791 66113
rect 99101 66147 99159 66153
rect 99101 66113 99113 66147
rect 99147 66113 99159 66147
rect 99101 66107 99159 66113
rect 95970 66076 95976 66088
rect 93872 66048 95976 66076
rect 95970 66036 95976 66048
rect 96028 66076 96034 66088
rect 98656 66076 98684 66107
rect 100202 66104 100208 66156
rect 100260 66104 100266 66156
rect 100389 66147 100447 66153
rect 100389 66113 100401 66147
rect 100435 66144 100447 66147
rect 102042 66144 102048 66156
rect 100435 66116 102048 66144
rect 100435 66113 100447 66116
rect 100389 66107 100447 66113
rect 102042 66104 102048 66116
rect 102100 66104 102106 66156
rect 108298 66104 108304 66156
rect 108356 66104 108362 66156
rect 96028 66048 98684 66076
rect 96028 66036 96034 66048
rect 92247 65980 92704 66008
rect 92753 66011 92811 66017
rect 92247 65977 92259 65980
rect 92201 65971 92259 65977
rect 92753 65977 92765 66011
rect 92799 66008 92811 66011
rect 92799 65980 93532 66008
rect 92799 65977 92811 65980
rect 92753 65971 92811 65977
rect 93504 65952 93532 65980
rect 93946 65968 93952 66020
rect 94004 66008 94010 66020
rect 94501 66011 94559 66017
rect 94501 66008 94513 66011
rect 94004 65980 94513 66008
rect 94004 65968 94010 65980
rect 94501 65977 94513 65980
rect 94547 66008 94559 66011
rect 94866 66008 94872 66020
rect 94547 65980 94872 66008
rect 94547 65977 94559 65980
rect 94501 65971 94559 65977
rect 94866 65968 94872 65980
rect 94924 65968 94930 66020
rect 98656 66008 98684 66048
rect 99377 66079 99435 66085
rect 99377 66045 99389 66079
rect 99423 66076 99435 66079
rect 99423 66048 100892 66076
rect 99423 66045 99435 66048
rect 99377 66039 99435 66045
rect 98656 65980 99374 66008
rect 90266 65940 90272 65952
rect 88536 65912 90272 65940
rect 90266 65900 90272 65912
rect 90324 65900 90330 65952
rect 91186 65900 91192 65952
rect 91244 65900 91250 65952
rect 93026 65900 93032 65952
rect 93084 65900 93090 65952
rect 93486 65900 93492 65952
rect 93544 65900 93550 65952
rect 94593 65943 94651 65949
rect 94593 65909 94605 65943
rect 94639 65940 94651 65943
rect 96614 65940 96620 65952
rect 94639 65912 96620 65940
rect 94639 65909 94651 65912
rect 94593 65903 94651 65909
rect 96614 65900 96620 65912
rect 96672 65900 96678 65952
rect 96798 65949 96804 65952
rect 96788 65943 96804 65949
rect 96788 65909 96800 65943
rect 96788 65903 96804 65909
rect 96798 65900 96804 65903
rect 96856 65900 96862 65952
rect 98362 65900 98368 65952
rect 98420 65900 98426 65952
rect 99346 65940 99374 65980
rect 99558 65968 99564 66020
rect 99616 66008 99622 66020
rect 100389 66011 100447 66017
rect 100389 66008 100401 66011
rect 99616 65980 100401 66008
rect 99616 65968 99622 65980
rect 100389 65977 100401 65980
rect 100435 65977 100447 66011
rect 100389 65971 100447 65977
rect 100202 65940 100208 65952
rect 99346 65912 100208 65940
rect 100202 65900 100208 65912
rect 100260 65940 100266 65952
rect 100570 65940 100576 65952
rect 100260 65912 100576 65940
rect 100260 65900 100266 65912
rect 100570 65900 100576 65912
rect 100628 65900 100634 65952
rect 100757 65943 100815 65949
rect 100757 65909 100769 65943
rect 100803 65940 100815 65943
rect 100864 65940 100892 66048
rect 108482 65968 108488 66020
rect 108540 65968 108546 66020
rect 103790 65940 103796 65952
rect 100803 65912 103796 65940
rect 100803 65909 100815 65912
rect 100757 65903 100815 65909
rect 103790 65900 103796 65912
rect 103848 65900 103854 65952
rect 1104 65850 108836 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 96374 65850
rect 96426 65798 96438 65850
rect 96490 65798 96502 65850
rect 96554 65798 96566 65850
rect 96618 65798 96630 65850
rect 96682 65798 105922 65850
rect 105974 65798 105986 65850
rect 106038 65798 106050 65850
rect 106102 65798 106114 65850
rect 106166 65798 106178 65850
rect 106230 65798 108836 65850
rect 1104 65776 108836 65798
rect 86954 65696 86960 65748
rect 87012 65736 87018 65748
rect 93026 65736 93032 65748
rect 87012 65708 93032 65736
rect 87012 65696 87018 65708
rect 93026 65696 93032 65708
rect 93084 65736 93090 65748
rect 103882 65736 103888 65748
rect 93084 65708 103888 65736
rect 93084 65696 93090 65708
rect 103882 65696 103888 65708
rect 103940 65696 103946 65748
rect 87782 65628 87788 65680
rect 87840 65668 87846 65680
rect 89622 65668 89628 65680
rect 87840 65640 89628 65668
rect 87840 65628 87846 65640
rect 89622 65628 89628 65640
rect 89680 65628 89686 65680
rect 91186 65628 91192 65680
rect 91244 65668 91250 65680
rect 108298 65668 108304 65680
rect 91244 65640 108304 65668
rect 91244 65628 91250 65640
rect 108298 65628 108304 65640
rect 108356 65628 108362 65680
rect 75914 65560 75920 65612
rect 75972 65600 75978 65612
rect 86494 65600 86500 65612
rect 75972 65572 86500 65600
rect 75972 65560 75978 65572
rect 86494 65560 86500 65572
rect 86552 65560 86558 65612
rect 88058 65560 88064 65612
rect 88116 65600 88122 65612
rect 91738 65600 91744 65612
rect 88116 65572 91744 65600
rect 88116 65560 88122 65572
rect 91738 65560 91744 65572
rect 91796 65560 91802 65612
rect 100570 65560 100576 65612
rect 100628 65600 100634 65612
rect 104158 65600 104164 65612
rect 100628 65572 104164 65600
rect 100628 65560 100634 65572
rect 104158 65560 104164 65572
rect 104216 65560 104222 65612
rect 1581 65535 1639 65541
rect 1581 65501 1593 65535
rect 1627 65532 1639 65535
rect 1765 65535 1823 65541
rect 1765 65532 1777 65535
rect 1627 65504 1777 65532
rect 1627 65501 1639 65504
rect 1581 65495 1639 65501
rect 1765 65501 1777 65504
rect 1811 65532 1823 65535
rect 30098 65532 30104 65544
rect 1811 65504 30104 65532
rect 1811 65501 1823 65504
rect 1765 65495 1823 65501
rect 30098 65492 30104 65504
rect 30156 65492 30162 65544
rect 96706 65492 96712 65544
rect 96764 65532 96770 65544
rect 108117 65535 108175 65541
rect 108117 65532 108129 65535
rect 96764 65504 108129 65532
rect 96764 65492 96770 65504
rect 108117 65501 108129 65504
rect 108163 65532 108175 65535
rect 108301 65535 108359 65541
rect 108301 65532 108313 65535
rect 108163 65504 108313 65532
rect 108163 65501 108175 65504
rect 108117 65495 108175 65501
rect 108301 65501 108313 65504
rect 108347 65501 108359 65535
rect 108301 65495 108359 65501
rect 85574 65424 85580 65476
rect 85632 65464 85638 65476
rect 107562 65464 107568 65476
rect 85632 65436 107568 65464
rect 85632 65424 85638 65436
rect 107562 65424 107568 65436
rect 107620 65424 107626 65476
rect 842 65356 848 65408
rect 900 65396 906 65408
rect 1397 65399 1455 65405
rect 1397 65396 1409 65399
rect 900 65368 1409 65396
rect 900 65356 906 65368
rect 1397 65365 1409 65368
rect 1443 65365 1455 65399
rect 1397 65359 1455 65365
rect 93486 65356 93492 65408
rect 93544 65396 93550 65408
rect 104986 65396 104992 65408
rect 93544 65368 104992 65396
rect 93544 65356 93550 65368
rect 104986 65356 104992 65368
rect 105044 65356 105050 65408
rect 108482 65356 108488 65408
rect 108540 65356 108546 65408
rect 1104 65306 7912 65328
rect 1104 65254 4874 65306
rect 4926 65254 4938 65306
rect 4990 65254 5002 65306
rect 5054 65254 5066 65306
rect 5118 65254 5130 65306
rect 5182 65254 7912 65306
rect 98362 65288 98368 65340
rect 98420 65328 98426 65340
rect 103422 65328 103428 65340
rect 98420 65300 103428 65328
rect 98420 65288 98426 65300
rect 103422 65288 103428 65300
rect 103480 65288 103486 65340
rect 104052 65306 108836 65328
rect 1104 65232 7912 65254
rect 104052 65254 106658 65306
rect 106710 65254 106722 65306
rect 106774 65254 106786 65306
rect 106838 65254 106850 65306
rect 106902 65254 106914 65306
rect 106966 65254 108836 65306
rect 104052 65232 108836 65254
rect 96062 65152 96068 65204
rect 96120 65192 96126 65204
rect 104434 65192 104440 65204
rect 96120 65164 104440 65192
rect 96120 65152 96126 65164
rect 104434 65152 104440 65164
rect 104492 65152 104498 65204
rect 1581 65059 1639 65065
rect 1581 65025 1593 65059
rect 1627 65056 1639 65059
rect 1627 65028 1808 65056
rect 1627 65025 1639 65028
rect 1581 65019 1639 65025
rect 1394 64880 1400 64932
rect 1452 64880 1458 64932
rect 1780 64929 1808 65028
rect 87598 65016 87604 65068
rect 87656 65056 87662 65068
rect 108117 65059 108175 65065
rect 108117 65056 108129 65059
rect 87656 65028 108129 65056
rect 87656 65016 87662 65028
rect 108117 65025 108129 65028
rect 108163 65056 108175 65059
rect 108301 65059 108359 65065
rect 108301 65056 108313 65059
rect 108163 65028 108313 65056
rect 108163 65025 108175 65028
rect 108117 65019 108175 65025
rect 108301 65025 108313 65028
rect 108347 65025 108359 65059
rect 108301 65019 108359 65025
rect 1765 64923 1823 64929
rect 1765 64889 1777 64923
rect 1811 64920 1823 64923
rect 26142 64920 26148 64932
rect 1811 64892 26148 64920
rect 1811 64889 1823 64892
rect 1765 64883 1823 64889
rect 26142 64880 26148 64892
rect 26200 64880 26206 64932
rect 108482 64880 108488 64932
rect 108540 64880 108546 64932
rect 1104 64762 7912 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 7912 64762
rect 1104 64688 7912 64710
rect 104052 64762 108836 64784
rect 104052 64710 105922 64762
rect 105974 64710 105986 64762
rect 106038 64710 106050 64762
rect 106102 64710 106114 64762
rect 106166 64710 106178 64762
rect 106230 64710 108836 64762
rect 104052 64688 108836 64710
rect 1581 64447 1639 64453
rect 1581 64413 1593 64447
rect 1627 64444 1639 64447
rect 1765 64447 1823 64453
rect 1765 64444 1777 64447
rect 1627 64416 1777 64444
rect 1627 64413 1639 64416
rect 1581 64407 1639 64413
rect 1765 64413 1777 64416
rect 1811 64444 1823 64447
rect 22002 64444 22008 64456
rect 1811 64416 22008 64444
rect 1811 64413 1823 64416
rect 1765 64407 1823 64413
rect 22002 64404 22008 64416
rect 22060 64404 22066 64456
rect 88518 64404 88524 64456
rect 88576 64444 88582 64456
rect 108117 64447 108175 64453
rect 108117 64444 108129 64447
rect 88576 64416 108129 64444
rect 88576 64404 88582 64416
rect 108117 64413 108129 64416
rect 108163 64444 108175 64447
rect 108301 64447 108359 64453
rect 108301 64444 108313 64447
rect 108163 64416 108313 64444
rect 108163 64413 108175 64416
rect 108117 64407 108175 64413
rect 108301 64413 108313 64416
rect 108347 64413 108359 64447
rect 108301 64407 108359 64413
rect 842 64268 848 64320
rect 900 64308 906 64320
rect 1397 64311 1455 64317
rect 1397 64308 1409 64311
rect 900 64280 1409 64308
rect 900 64268 906 64280
rect 1397 64277 1409 64280
rect 1443 64277 1455 64311
rect 1397 64271 1455 64277
rect 1854 64268 1860 64320
rect 1912 64308 1918 64320
rect 10318 64308 10324 64320
rect 1912 64280 10324 64308
rect 1912 64268 1918 64280
rect 10318 64268 10324 64280
rect 10376 64268 10382 64320
rect 108482 64268 108488 64320
rect 108540 64268 108546 64320
rect 1104 64218 7912 64240
rect 1104 64166 4874 64218
rect 4926 64166 4938 64218
rect 4990 64166 5002 64218
rect 5054 64166 5066 64218
rect 5118 64166 5130 64218
rect 5182 64166 7912 64218
rect 104052 64218 108836 64240
rect 1104 64144 7912 64166
rect 77386 64132 77392 64184
rect 77444 64172 77450 64184
rect 102778 64172 102784 64184
rect 77444 64144 102784 64172
rect 77444 64132 77450 64144
rect 102778 64132 102784 64144
rect 102836 64132 102842 64184
rect 104052 64166 106658 64218
rect 106710 64166 106722 64218
rect 106774 64166 106786 64218
rect 106838 64166 106850 64218
rect 106902 64166 106914 64218
rect 106966 64166 108836 64218
rect 104052 64144 108836 64166
rect 1104 63674 7912 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 7912 63674
rect 1104 63600 7912 63622
rect 104052 63674 108836 63696
rect 104052 63622 105922 63674
rect 105974 63622 105986 63674
rect 106038 63622 106050 63674
rect 106102 63622 106114 63674
rect 106166 63622 106178 63674
rect 106230 63622 108836 63674
rect 104052 63600 108836 63622
rect 842 63452 848 63504
rect 900 63492 906 63504
rect 1397 63495 1455 63501
rect 1397 63492 1409 63495
rect 900 63464 1409 63492
rect 900 63452 906 63464
rect 1397 63461 1409 63464
rect 1443 63461 1455 63495
rect 1397 63455 1455 63461
rect 1765 63495 1823 63501
rect 1765 63461 1777 63495
rect 1811 63492 1823 63495
rect 2774 63492 2780 63504
rect 1811 63464 2780 63492
rect 1811 63461 1823 63464
rect 1765 63455 1823 63461
rect 1581 63359 1639 63365
rect 1581 63325 1593 63359
rect 1627 63356 1639 63359
rect 1780 63356 1808 63455
rect 2774 63452 2780 63464
rect 2832 63452 2838 63504
rect 1627 63328 1808 63356
rect 1627 63325 1639 63328
rect 1581 63319 1639 63325
rect 1104 63130 7912 63152
rect 1104 63078 4874 63130
rect 4926 63078 4938 63130
rect 4990 63078 5002 63130
rect 5054 63078 5066 63130
rect 5118 63078 5130 63130
rect 5182 63078 7912 63130
rect 1104 63056 7912 63078
rect 104052 63130 108836 63152
rect 104052 63078 106658 63130
rect 106710 63078 106722 63130
rect 106774 63078 106786 63130
rect 106838 63078 106850 63130
rect 106902 63078 106914 63130
rect 106966 63078 108836 63130
rect 104052 63056 108836 63078
rect 1765 63019 1823 63025
rect 1765 62985 1777 63019
rect 1811 63016 1823 63019
rect 3418 63016 3424 63028
rect 1811 62988 3424 63016
rect 1811 62985 1823 62988
rect 1765 62979 1823 62985
rect 1581 62883 1639 62889
rect 1581 62849 1593 62883
rect 1627 62880 1639 62883
rect 1780 62880 1808 62979
rect 3418 62976 3424 62988
rect 3476 62976 3482 63028
rect 1627 62852 1808 62880
rect 1627 62849 1639 62852
rect 1581 62843 1639 62849
rect 842 62704 848 62756
rect 900 62744 906 62756
rect 1397 62747 1455 62753
rect 1397 62744 1409 62747
rect 900 62716 1409 62744
rect 900 62704 906 62716
rect 1397 62713 1409 62716
rect 1443 62713 1455 62747
rect 1397 62707 1455 62713
rect 1104 62586 7912 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 7912 62586
rect 1104 62512 7912 62534
rect 104052 62586 108836 62608
rect 104052 62534 105922 62586
rect 105974 62534 105986 62586
rect 106038 62534 106050 62586
rect 106102 62534 106114 62586
rect 106166 62534 106178 62586
rect 106230 62534 108836 62586
rect 104052 62512 108836 62534
rect 1581 62475 1639 62481
rect 1581 62441 1593 62475
rect 1627 62472 1639 62475
rect 1854 62472 1860 62484
rect 1627 62444 1860 62472
rect 1627 62441 1639 62444
rect 1581 62435 1639 62441
rect 1854 62432 1860 62444
rect 1912 62432 1918 62484
rect 1486 62160 1492 62212
rect 1544 62200 1550 62212
rect 1949 62203 2007 62209
rect 1949 62200 1961 62203
rect 1544 62172 1961 62200
rect 1544 62160 1550 62172
rect 1949 62169 1961 62172
rect 1995 62169 2007 62203
rect 1949 62163 2007 62169
rect 1104 62042 7912 62064
rect 1104 61990 4874 62042
rect 4926 61990 4938 62042
rect 4990 61990 5002 62042
rect 5054 61990 5066 62042
rect 5118 61990 5130 62042
rect 5182 61990 7912 62042
rect 1104 61968 7912 61990
rect 104052 62042 108836 62064
rect 104052 61990 106658 62042
rect 106710 61990 106722 62042
rect 106774 61990 106786 62042
rect 106838 61990 106850 62042
rect 106902 61990 106914 62042
rect 106966 61990 108836 62042
rect 104052 61968 108836 61990
rect 1670 61820 1676 61872
rect 1728 61860 1734 61872
rect 1765 61863 1823 61869
rect 1765 61860 1777 61863
rect 1728 61832 1777 61860
rect 1728 61820 1734 61832
rect 1765 61829 1777 61832
rect 1811 61829 1823 61863
rect 1765 61823 1823 61829
rect 1302 61752 1308 61804
rect 1360 61792 1366 61804
rect 1489 61795 1547 61801
rect 1489 61792 1501 61795
rect 1360 61764 1501 61792
rect 1360 61752 1366 61764
rect 1489 61761 1501 61764
rect 1535 61792 1547 61795
rect 1949 61795 2007 61801
rect 1949 61792 1961 61795
rect 1535 61764 1961 61792
rect 1535 61761 1547 61764
rect 1489 61755 1547 61761
rect 1949 61761 1961 61764
rect 1995 61761 2007 61795
rect 1949 61755 2007 61761
rect 1104 61498 7912 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 7912 61498
rect 1104 61424 7912 61446
rect 104052 61498 108836 61520
rect 104052 61446 105922 61498
rect 105974 61446 105986 61498
rect 106038 61446 106050 61498
rect 106102 61446 106114 61498
rect 106166 61446 106178 61498
rect 106230 61446 108836 61498
rect 104052 61424 108836 61446
rect 1104 60954 7912 60976
rect 1104 60902 4874 60954
rect 4926 60902 4938 60954
rect 4990 60902 5002 60954
rect 5054 60902 5066 60954
rect 5118 60902 5130 60954
rect 5182 60902 7912 60954
rect 1104 60880 7912 60902
rect 104052 60954 108836 60976
rect 104052 60902 106658 60954
rect 106710 60902 106722 60954
rect 106774 60902 106786 60954
rect 106838 60902 106850 60954
rect 106902 60902 106914 60954
rect 106966 60902 108836 60954
rect 104052 60880 108836 60902
rect 1104 60410 7912 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 7912 60410
rect 1104 60336 7912 60358
rect 104052 60410 108836 60432
rect 104052 60358 105922 60410
rect 105974 60358 105986 60410
rect 106038 60358 106050 60410
rect 106102 60358 106114 60410
rect 106166 60358 106178 60410
rect 106230 60358 108836 60410
rect 104052 60336 108836 60358
rect 103974 60052 103980 60104
rect 104032 60092 104038 60104
rect 104345 60095 104403 60101
rect 104345 60092 104357 60095
rect 104032 60064 104357 60092
rect 104032 60052 104038 60064
rect 104345 60061 104357 60064
rect 104391 60061 104403 60095
rect 104345 60055 104403 60061
rect 1104 59866 7912 59888
rect 1104 59814 4874 59866
rect 4926 59814 4938 59866
rect 4990 59814 5002 59866
rect 5054 59814 5066 59866
rect 5118 59814 5130 59866
rect 5182 59814 7912 59866
rect 1104 59792 7912 59814
rect 104052 59866 108836 59888
rect 104052 59814 106658 59866
rect 106710 59814 106722 59866
rect 106774 59814 106786 59866
rect 106838 59814 106850 59866
rect 106902 59814 106914 59866
rect 106966 59814 108836 59866
rect 104052 59792 108836 59814
rect 104434 59712 104440 59764
rect 104492 59712 104498 59764
rect 103422 59576 103428 59628
rect 103480 59616 103486 59628
rect 104345 59619 104403 59625
rect 104345 59616 104357 59619
rect 103480 59588 104357 59616
rect 103480 59576 103486 59588
rect 104345 59585 104357 59588
rect 104391 59585 104403 59619
rect 104345 59579 104403 59585
rect 104529 59619 104587 59625
rect 104529 59585 104541 59619
rect 104575 59585 104587 59619
rect 104529 59579 104587 59585
rect 103974 59508 103980 59560
rect 104032 59548 104038 59560
rect 104544 59548 104572 59579
rect 104032 59520 104572 59548
rect 104032 59508 104038 59520
rect 1104 59322 7912 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 7912 59322
rect 1104 59248 7912 59270
rect 104052 59322 108836 59344
rect 104052 59270 105922 59322
rect 105974 59270 105986 59322
rect 106038 59270 106050 59322
rect 106102 59270 106114 59322
rect 106166 59270 106178 59322
rect 106230 59270 108836 59322
rect 104052 59248 108836 59270
rect 1104 58778 7912 58800
rect 1104 58726 4874 58778
rect 4926 58726 4938 58778
rect 4990 58726 5002 58778
rect 5054 58726 5066 58778
rect 5118 58726 5130 58778
rect 5182 58726 7912 58778
rect 1104 58704 7912 58726
rect 104052 58778 108836 58800
rect 104052 58726 106658 58778
rect 106710 58726 106722 58778
rect 106774 58726 106786 58778
rect 106838 58726 106850 58778
rect 106902 58726 106914 58778
rect 106966 58726 108836 58778
rect 104052 58704 108836 58726
rect 105630 58624 105636 58676
rect 105688 58664 105694 58676
rect 105814 58664 105820 58676
rect 105688 58636 105820 58664
rect 105688 58624 105694 58636
rect 105814 58624 105820 58636
rect 105872 58664 105878 58676
rect 106185 58667 106243 58673
rect 106185 58664 106197 58667
rect 105872 58636 106197 58664
rect 105872 58624 105878 58636
rect 106185 58633 106197 58636
rect 106231 58633 106243 58667
rect 106185 58627 106243 58633
rect 104342 58556 104348 58608
rect 104400 58556 104406 58608
rect 1104 58234 7912 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 7912 58234
rect 1104 58160 7912 58182
rect 104052 58234 108836 58256
rect 104052 58182 105922 58234
rect 105974 58182 105986 58234
rect 106038 58182 106050 58234
rect 106102 58182 106114 58234
rect 106166 58182 106178 58234
rect 106230 58182 108836 58234
rect 104052 58160 108836 58182
rect 104342 58080 104348 58132
rect 104400 58080 104406 58132
rect 1104 57690 7912 57712
rect 1104 57638 4874 57690
rect 4926 57638 4938 57690
rect 4990 57638 5002 57690
rect 5054 57638 5066 57690
rect 5118 57638 5130 57690
rect 5182 57638 7912 57690
rect 1104 57616 7912 57638
rect 104052 57690 108836 57712
rect 104052 57638 106658 57690
rect 106710 57638 106722 57690
rect 106774 57638 106786 57690
rect 106838 57638 106850 57690
rect 106902 57638 106914 57690
rect 106966 57638 108836 57690
rect 104052 57616 108836 57638
rect 104250 57536 104256 57588
rect 104308 57576 104314 57588
rect 104526 57576 104532 57588
rect 104308 57548 104532 57576
rect 104308 57536 104314 57548
rect 104526 57536 104532 57548
rect 104584 57536 104590 57588
rect 103790 57468 103796 57520
rect 103848 57508 103854 57520
rect 104345 57511 104403 57517
rect 104345 57508 104357 57511
rect 103848 57480 104357 57508
rect 103848 57468 103854 57480
rect 104345 57477 104357 57480
rect 104391 57508 104403 57511
rect 104710 57508 104716 57520
rect 104391 57480 104716 57508
rect 104391 57477 104403 57480
rect 104345 57471 104403 57477
rect 104710 57468 104716 57480
rect 104768 57468 104774 57520
rect 1104 57146 7912 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 7912 57146
rect 1104 57072 7912 57094
rect 104052 57146 108836 57168
rect 104052 57094 105922 57146
rect 105974 57094 105986 57146
rect 106038 57094 106050 57146
rect 106102 57094 106114 57146
rect 106166 57094 106178 57146
rect 106230 57094 108836 57146
rect 104052 57072 108836 57094
rect 104986 56992 104992 57044
rect 105044 57032 105050 57044
rect 105265 57035 105323 57041
rect 105265 57032 105277 57035
rect 105044 57004 105277 57032
rect 105044 56992 105050 57004
rect 105265 57001 105277 57004
rect 105311 57001 105323 57035
rect 105265 56995 105323 57001
rect 104158 56856 104164 56908
rect 104216 56896 104222 56908
rect 104345 56899 104403 56905
rect 104345 56896 104357 56899
rect 104216 56868 104357 56896
rect 104216 56856 104222 56868
rect 104345 56865 104357 56868
rect 104391 56865 104403 56899
rect 104345 56859 104403 56865
rect 104434 56856 104440 56908
rect 104492 56896 104498 56908
rect 104710 56896 104716 56908
rect 104492 56868 104716 56896
rect 104492 56856 104498 56868
rect 104710 56856 104716 56868
rect 104768 56856 104774 56908
rect 104802 56856 104808 56908
rect 104860 56896 104866 56908
rect 105081 56899 105139 56905
rect 105081 56896 105093 56899
rect 104860 56868 105093 56896
rect 104860 56856 104866 56868
rect 105081 56865 105093 56868
rect 105127 56865 105139 56899
rect 105081 56859 105139 56865
rect 104250 56788 104256 56840
rect 104308 56828 104314 56840
rect 104820 56828 104848 56856
rect 104308 56800 104848 56828
rect 104308 56788 104314 56800
rect 104342 56652 104348 56704
rect 104400 56692 104406 56704
rect 104437 56695 104495 56701
rect 104437 56692 104449 56695
rect 104400 56664 104449 56692
rect 104400 56652 104406 56664
rect 104437 56661 104449 56664
rect 104483 56661 104495 56695
rect 104437 56655 104495 56661
rect 104526 56652 104532 56704
rect 104584 56652 104590 56704
rect 1104 56602 7912 56624
rect 1104 56550 4874 56602
rect 4926 56550 4938 56602
rect 4990 56550 5002 56602
rect 5054 56550 5066 56602
rect 5118 56550 5130 56602
rect 5182 56550 7912 56602
rect 1104 56528 7912 56550
rect 104052 56602 108836 56624
rect 104052 56550 106658 56602
rect 106710 56550 106722 56602
rect 106774 56550 106786 56602
rect 106838 56550 106850 56602
rect 106902 56550 106914 56602
rect 106966 56550 108836 56602
rect 104052 56528 108836 56550
rect 104158 56448 104164 56500
rect 104216 56488 104222 56500
rect 104710 56488 104716 56500
rect 104216 56460 104716 56488
rect 104216 56448 104222 56460
rect 104710 56448 104716 56460
rect 104768 56448 104774 56500
rect 104618 56380 104624 56432
rect 104676 56420 104682 56432
rect 104897 56423 104955 56429
rect 104897 56420 104909 56423
rect 104676 56392 104909 56420
rect 104676 56380 104682 56392
rect 104897 56389 104909 56392
rect 104943 56389 104955 56423
rect 104897 56383 104955 56389
rect 104342 56312 104348 56364
rect 104400 56352 104406 56364
rect 104437 56355 104495 56361
rect 104437 56352 104449 56355
rect 104400 56324 104449 56352
rect 104400 56312 104406 56324
rect 104437 56321 104449 56324
rect 104483 56321 104495 56355
rect 104437 56315 104495 56321
rect 1104 56058 7912 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 7912 56058
rect 1104 55984 7912 56006
rect 104052 56058 108836 56080
rect 104052 56006 105922 56058
rect 105974 56006 105986 56058
rect 106038 56006 106050 56058
rect 106102 56006 106114 56058
rect 106166 56006 106178 56058
rect 106230 56006 108836 56058
rect 104052 55984 108836 56006
rect 1104 55514 7912 55536
rect 1104 55462 4874 55514
rect 4926 55462 4938 55514
rect 4990 55462 5002 55514
rect 5054 55462 5066 55514
rect 5118 55462 5130 55514
rect 5182 55462 7912 55514
rect 1104 55440 7912 55462
rect 104052 55514 108836 55536
rect 104052 55462 106658 55514
rect 106710 55462 106722 55514
rect 106774 55462 106786 55514
rect 106838 55462 106850 55514
rect 106902 55462 106914 55514
rect 106966 55462 108836 55514
rect 104052 55440 108836 55462
rect 103790 55360 103796 55412
rect 103848 55400 103854 55412
rect 104437 55403 104495 55409
rect 104437 55400 104449 55403
rect 103848 55372 104449 55400
rect 103848 55360 103854 55372
rect 104437 55369 104449 55372
rect 104483 55400 104495 55403
rect 104897 55403 104955 55409
rect 104897 55400 104909 55403
rect 104483 55372 104909 55400
rect 104483 55369 104495 55372
rect 104437 55363 104495 55369
rect 104897 55369 104909 55372
rect 104943 55369 104955 55403
rect 104897 55363 104955 55369
rect 104526 55292 104532 55344
rect 104584 55332 104590 55344
rect 104713 55335 104771 55341
rect 104713 55332 104725 55335
rect 104584 55304 104725 55332
rect 104584 55292 104590 55304
rect 104636 55273 104664 55304
rect 104713 55301 104725 55304
rect 104759 55301 104771 55335
rect 104713 55295 104771 55301
rect 104621 55267 104679 55273
rect 104621 55233 104633 55267
rect 104667 55264 104679 55267
rect 104667 55236 104701 55264
rect 104667 55233 104679 55236
rect 104621 55227 104679 55233
rect 1104 54970 7912 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 7912 54970
rect 1104 54896 7912 54918
rect 104052 54970 108836 54992
rect 104052 54918 105922 54970
rect 105974 54918 105986 54970
rect 106038 54918 106050 54970
rect 106102 54918 106114 54970
rect 106166 54918 106178 54970
rect 106230 54918 108836 54970
rect 104052 54896 108836 54918
rect 103882 54816 103888 54868
rect 103940 54856 103946 54868
rect 104897 54859 104955 54865
rect 104897 54856 104909 54859
rect 103940 54828 104909 54856
rect 103940 54816 103946 54828
rect 104897 54825 104909 54828
rect 104943 54856 104955 54859
rect 105265 54859 105323 54865
rect 105265 54856 105277 54859
rect 104943 54828 105277 54856
rect 104943 54825 104955 54828
rect 104897 54819 104955 54825
rect 105265 54825 105277 54828
rect 105311 54825 105323 54859
rect 105265 54819 105323 54825
rect 104345 54791 104403 54797
rect 104345 54757 104357 54791
rect 104391 54788 104403 54791
rect 104434 54788 104440 54800
rect 104391 54760 104440 54788
rect 104391 54757 104403 54760
rect 104345 54751 104403 54757
rect 104434 54748 104440 54760
rect 104492 54748 104498 54800
rect 104526 54612 104532 54664
rect 104584 54612 104590 54664
rect 105081 54587 105139 54593
rect 105081 54584 105093 54587
rect 104636 54556 105093 54584
rect 104636 54528 104664 54556
rect 105081 54553 105093 54556
rect 105127 54553 105139 54587
rect 105081 54547 105139 54553
rect 104618 54476 104624 54528
rect 104676 54476 104682 54528
rect 104710 54476 104716 54528
rect 104768 54476 104774 54528
rect 1104 54426 7912 54448
rect 1104 54374 4874 54426
rect 4926 54374 4938 54426
rect 4990 54374 5002 54426
rect 5054 54374 5066 54426
rect 5118 54374 5130 54426
rect 5182 54374 7912 54426
rect 1104 54352 7912 54374
rect 104052 54426 108836 54448
rect 104052 54374 106658 54426
rect 106710 54374 106722 54426
rect 106774 54374 106786 54426
rect 106838 54374 106850 54426
rect 106902 54374 106914 54426
rect 106966 54374 108836 54426
rect 104052 54352 108836 54374
rect 104434 54272 104440 54324
rect 104492 54272 104498 54324
rect 104526 54272 104532 54324
rect 104584 54272 104590 54324
rect 1104 53882 7912 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 7912 53882
rect 1104 53808 7912 53830
rect 104052 53882 108836 53904
rect 104052 53830 105922 53882
rect 105974 53830 105986 53882
rect 106038 53830 106050 53882
rect 106102 53830 106114 53882
rect 106166 53830 106178 53882
rect 106230 53830 108836 53882
rect 104052 53808 108836 53830
rect 1104 53338 7912 53360
rect 1104 53286 4874 53338
rect 4926 53286 4938 53338
rect 4990 53286 5002 53338
rect 5054 53286 5066 53338
rect 5118 53286 5130 53338
rect 5182 53286 7912 53338
rect 1104 53264 7912 53286
rect 104052 53338 108836 53360
rect 104052 53286 106658 53338
rect 106710 53286 106722 53338
rect 106774 53286 106786 53338
rect 106838 53286 106850 53338
rect 106902 53286 106914 53338
rect 106966 53286 108836 53338
rect 104052 53264 108836 53286
rect 1104 52794 7912 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 7912 52794
rect 1104 52720 7912 52742
rect 104052 52794 108836 52816
rect 104052 52742 105922 52794
rect 105974 52742 105986 52794
rect 106038 52742 106050 52794
rect 106102 52742 106114 52794
rect 106166 52742 106178 52794
rect 106230 52742 108836 52794
rect 104052 52720 108836 52742
rect 1104 52250 7912 52272
rect 1104 52198 4874 52250
rect 4926 52198 4938 52250
rect 4990 52198 5002 52250
rect 5054 52198 5066 52250
rect 5118 52198 5130 52250
rect 5182 52198 7912 52250
rect 1104 52176 7912 52198
rect 104052 52250 108836 52272
rect 104052 52198 106658 52250
rect 106710 52198 106722 52250
rect 106774 52198 106786 52250
rect 106838 52198 106850 52250
rect 106902 52198 106914 52250
rect 106966 52198 108836 52250
rect 104052 52176 108836 52198
rect 104437 52139 104495 52145
rect 104437 52105 104449 52139
rect 104483 52136 104495 52139
rect 104526 52136 104532 52148
rect 104483 52108 104532 52136
rect 104483 52105 104495 52108
rect 104437 52099 104495 52105
rect 104526 52096 104532 52108
rect 104584 52096 104590 52148
rect 1104 51706 7912 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 7912 51706
rect 1104 51632 7912 51654
rect 104052 51706 108836 51728
rect 104052 51654 105922 51706
rect 105974 51654 105986 51706
rect 106038 51654 106050 51706
rect 106102 51654 106114 51706
rect 106166 51654 106178 51706
rect 106230 51654 108836 51706
rect 104052 51632 108836 51654
rect 104526 51552 104532 51604
rect 104584 51552 104590 51604
rect 103974 51484 103980 51536
rect 104032 51524 104038 51536
rect 104713 51527 104771 51533
rect 104713 51524 104725 51527
rect 104032 51496 104725 51524
rect 104032 51484 104038 51496
rect 104636 51400 104664 51496
rect 104713 51493 104725 51496
rect 104759 51493 104771 51527
rect 104713 51487 104771 51493
rect 104618 51348 104624 51400
rect 104676 51348 104682 51400
rect 105173 51391 105231 51397
rect 105173 51388 105185 51391
rect 104912 51360 105185 51388
rect 104345 51323 104403 51329
rect 104345 51289 104357 51323
rect 104391 51320 104403 51323
rect 104434 51320 104440 51332
rect 104391 51292 104440 51320
rect 104391 51289 104403 51292
rect 104345 51283 104403 51289
rect 104434 51280 104440 51292
rect 104492 51320 104498 51332
rect 104912 51329 104940 51360
rect 105173 51357 105185 51360
rect 105219 51357 105231 51391
rect 105173 51351 105231 51357
rect 108209 51391 108267 51397
rect 108209 51357 108221 51391
rect 108255 51388 108267 51391
rect 108482 51388 108488 51400
rect 108255 51360 108488 51388
rect 108255 51357 108267 51360
rect 108209 51351 108267 51357
rect 108482 51348 108488 51360
rect 108540 51348 108546 51400
rect 104897 51323 104955 51329
rect 104897 51320 104909 51323
rect 104492 51292 104909 51320
rect 104492 51280 104498 51292
rect 104897 51289 104909 51292
rect 104943 51289 104955 51323
rect 104897 51283 104955 51289
rect 105081 51323 105139 51329
rect 105081 51289 105093 51323
rect 105127 51320 105139 51323
rect 105127 51292 105400 51320
rect 105127 51289 105139 51292
rect 105081 51283 105139 51289
rect 105372 51264 105400 51292
rect 104526 51212 104532 51264
rect 104584 51261 104590 51264
rect 104584 51255 104603 51261
rect 104591 51221 104603 51255
rect 104584 51215 104603 51221
rect 104584 51212 104590 51215
rect 105354 51212 105360 51264
rect 105412 51212 105418 51264
rect 108298 51212 108304 51264
rect 108356 51212 108362 51264
rect 1104 51162 7912 51184
rect 1104 51110 4874 51162
rect 4926 51110 4938 51162
rect 4990 51110 5002 51162
rect 5054 51110 5066 51162
rect 5118 51110 5130 51162
rect 5182 51110 7912 51162
rect 1104 51088 7912 51110
rect 104052 51162 108836 51184
rect 104052 51110 106658 51162
rect 106710 51110 106722 51162
rect 106774 51110 106786 51162
rect 106838 51110 106850 51162
rect 106902 51110 106914 51162
rect 106966 51110 108836 51162
rect 104052 51088 108836 51110
rect 104434 51008 104440 51060
rect 104492 51008 104498 51060
rect 104526 51008 104532 51060
rect 104584 51008 104590 51060
rect 1104 50618 7912 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 7912 50618
rect 1104 50544 7912 50566
rect 104052 50618 108836 50640
rect 104052 50566 105922 50618
rect 105974 50566 105986 50618
rect 106038 50566 106050 50618
rect 106102 50566 106114 50618
rect 106166 50566 106178 50618
rect 106230 50566 108836 50618
rect 104052 50544 108836 50566
rect 1104 50074 7912 50096
rect 1104 50022 4874 50074
rect 4926 50022 4938 50074
rect 4990 50022 5002 50074
rect 5054 50022 5066 50074
rect 5118 50022 5130 50074
rect 5182 50022 7912 50074
rect 1104 50000 7912 50022
rect 104052 50074 108836 50096
rect 104052 50022 106658 50074
rect 106710 50022 106722 50074
rect 106774 50022 106786 50074
rect 106838 50022 106850 50074
rect 106902 50022 106914 50074
rect 106966 50022 108836 50074
rect 104052 50000 108836 50022
rect 104710 49920 104716 49972
rect 104768 49920 104774 49972
rect 104250 49852 104256 49904
rect 104308 49892 104314 49904
rect 104989 49895 105047 49901
rect 104989 49892 105001 49895
rect 104308 49864 105001 49892
rect 104308 49852 104314 49864
rect 104342 49784 104348 49836
rect 104400 49784 104406 49836
rect 104544 49833 104572 49864
rect 104989 49861 105001 49864
rect 105035 49892 105047 49895
rect 105173 49895 105231 49901
rect 105173 49892 105185 49895
rect 105035 49864 105185 49892
rect 105035 49861 105047 49864
rect 104989 49855 105047 49861
rect 105173 49861 105185 49864
rect 105219 49861 105231 49895
rect 105173 49855 105231 49861
rect 104529 49827 104587 49833
rect 104529 49793 104541 49827
rect 104575 49793 104587 49827
rect 104529 49787 104587 49793
rect 104802 49716 104808 49768
rect 104860 49756 104866 49768
rect 105357 49759 105415 49765
rect 105357 49756 105369 49759
rect 104860 49728 105369 49756
rect 104860 49716 104866 49728
rect 105357 49725 105369 49728
rect 105403 49725 105415 49759
rect 105357 49719 105415 49725
rect 1104 49530 7912 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 7912 49530
rect 1104 49456 7912 49478
rect 104052 49530 108836 49552
rect 104052 49478 105922 49530
rect 105974 49478 105986 49530
rect 106038 49478 106050 49530
rect 106102 49478 106114 49530
rect 106166 49478 106178 49530
rect 106230 49478 108836 49530
rect 104052 49456 108836 49478
rect 104250 49376 104256 49428
rect 104308 49416 104314 49428
rect 104345 49419 104403 49425
rect 104345 49416 104357 49419
rect 104308 49388 104357 49416
rect 104308 49376 104314 49388
rect 104345 49385 104357 49388
rect 104391 49385 104403 49419
rect 104345 49379 104403 49385
rect 1104 48986 7912 49008
rect 1104 48934 4874 48986
rect 4926 48934 4938 48986
rect 4990 48934 5002 48986
rect 5054 48934 5066 48986
rect 5118 48934 5130 48986
rect 5182 48934 7912 48986
rect 1104 48912 7912 48934
rect 104052 48986 108836 49008
rect 104052 48934 106658 48986
rect 106710 48934 106722 48986
rect 106774 48934 106786 48986
rect 106838 48934 106850 48986
rect 106902 48934 106914 48986
rect 106966 48934 108836 48986
rect 104052 48912 108836 48934
rect 1104 48442 7912 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 7912 48442
rect 1104 48368 7912 48390
rect 104052 48442 108836 48464
rect 104052 48390 105922 48442
rect 105974 48390 105986 48442
rect 106038 48390 106050 48442
rect 106102 48390 106114 48442
rect 106166 48390 106178 48442
rect 106230 48390 108836 48442
rect 104052 48368 108836 48390
rect 1104 47898 7912 47920
rect 1104 47846 4874 47898
rect 4926 47846 4938 47898
rect 4990 47846 5002 47898
rect 5054 47846 5066 47898
rect 5118 47846 5130 47898
rect 5182 47846 7912 47898
rect 1104 47824 7912 47846
rect 104052 47898 108836 47920
rect 104052 47846 106658 47898
rect 106710 47846 106722 47898
rect 106774 47846 106786 47898
rect 106838 47846 106850 47898
rect 106902 47846 106914 47898
rect 106966 47846 108836 47898
rect 104052 47824 108836 47846
rect 1104 47354 7912 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 7912 47354
rect 1104 47280 7912 47302
rect 104052 47354 108836 47376
rect 104052 47302 105922 47354
rect 105974 47302 105986 47354
rect 106038 47302 106050 47354
rect 106102 47302 106114 47354
rect 106166 47302 106178 47354
rect 106230 47302 108836 47354
rect 104052 47280 108836 47302
rect 1104 46810 7912 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 7912 46810
rect 1104 46736 7912 46758
rect 104052 46810 108836 46832
rect 104052 46758 106658 46810
rect 106710 46758 106722 46810
rect 106774 46758 106786 46810
rect 106838 46758 106850 46810
rect 106902 46758 106914 46810
rect 106966 46758 108836 46810
rect 104052 46736 108836 46758
rect 1104 46266 7912 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 7912 46266
rect 1104 46192 7912 46214
rect 104052 46266 108836 46288
rect 104052 46214 105922 46266
rect 105974 46214 105986 46266
rect 106038 46214 106050 46266
rect 106102 46214 106114 46266
rect 106166 46214 106178 46266
rect 106230 46214 108836 46266
rect 104052 46192 108836 46214
rect 104342 46112 104348 46164
rect 104400 46112 104406 46164
rect 104250 45908 104256 45960
rect 104308 45948 104314 45960
rect 104529 45951 104587 45957
rect 104529 45948 104541 45951
rect 104308 45920 104541 45948
rect 104308 45908 104314 45920
rect 104529 45917 104541 45920
rect 104575 45917 104587 45951
rect 104529 45911 104587 45917
rect 1104 45722 7912 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 7912 45722
rect 1104 45648 7912 45670
rect 104052 45722 108836 45744
rect 104052 45670 106658 45722
rect 106710 45670 106722 45722
rect 106774 45670 106786 45722
rect 106838 45670 106850 45722
rect 106902 45670 106914 45722
rect 106966 45670 108836 45722
rect 104052 45648 108836 45670
rect 104713 45475 104771 45481
rect 104713 45441 104725 45475
rect 104759 45472 104771 45475
rect 105078 45472 105084 45484
rect 104759 45444 105084 45472
rect 104759 45441 104771 45444
rect 104713 45435 104771 45441
rect 105078 45432 105084 45444
rect 105136 45432 105142 45484
rect 104618 45364 104624 45416
rect 104676 45364 104682 45416
rect 104345 45271 104403 45277
rect 104345 45237 104357 45271
rect 104391 45268 104403 45271
rect 105170 45268 105176 45280
rect 104391 45240 105176 45268
rect 104391 45237 104403 45240
rect 104345 45231 104403 45237
rect 105170 45228 105176 45240
rect 105228 45228 105234 45280
rect 1104 45178 7912 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 7912 45178
rect 1104 45104 7912 45126
rect 104052 45178 108836 45200
rect 104052 45126 105922 45178
rect 105974 45126 105986 45178
rect 106038 45126 106050 45178
rect 106102 45126 106114 45178
rect 106166 45126 106178 45178
rect 106230 45126 108836 45178
rect 104052 45104 108836 45126
rect 102778 44888 102784 44940
rect 102836 44928 102842 44940
rect 104437 44931 104495 44937
rect 104437 44928 104449 44931
rect 102836 44900 104449 44928
rect 102836 44888 102842 44900
rect 1104 44634 7912 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 7912 44634
rect 1104 44560 7912 44582
rect 103992 44384 104020 44900
rect 104437 44897 104449 44900
rect 104483 44928 104495 44931
rect 105173 44931 105231 44937
rect 105173 44928 105185 44931
rect 104483 44900 105185 44928
rect 104483 44897 104495 44900
rect 104437 44891 104495 44897
rect 105173 44897 105185 44900
rect 105219 44897 105231 44931
rect 105173 44891 105231 44897
rect 104989 44863 105047 44869
rect 104989 44829 105001 44863
rect 105035 44860 105047 44863
rect 108298 44860 108304 44872
rect 105035 44832 108304 44860
rect 105035 44829 105047 44832
rect 104989 44823 105047 44829
rect 108298 44820 108304 44832
rect 108356 44820 108362 44872
rect 104052 44634 108836 44656
rect 104052 44582 106658 44634
rect 106710 44582 106722 44634
rect 106774 44582 106786 44634
rect 106838 44582 106850 44634
rect 106902 44582 106914 44634
rect 106966 44582 108836 44634
rect 104052 44560 108836 44582
rect 105541 44455 105599 44461
rect 105541 44452 105553 44455
rect 104360 44424 105553 44452
rect 104360 44393 104388 44424
rect 105541 44421 105553 44424
rect 105587 44421 105599 44455
rect 105541 44415 105599 44421
rect 104345 44387 104403 44393
rect 104345 44384 104357 44387
rect 103992 44356 104357 44384
rect 104345 44353 104357 44356
rect 104391 44353 104403 44387
rect 105081 44387 105139 44393
rect 105081 44384 105093 44387
rect 104345 44347 104403 44353
rect 104544 44356 105093 44384
rect 103698 44276 103704 44328
rect 103756 44316 103762 44328
rect 104544 44325 104572 44356
rect 105081 44353 105093 44356
rect 105127 44384 105139 44387
rect 105173 44387 105231 44393
rect 105173 44384 105185 44387
rect 105127 44356 105185 44384
rect 105127 44353 105139 44356
rect 105081 44347 105139 44353
rect 105173 44353 105185 44356
rect 105219 44384 105231 44387
rect 105357 44387 105415 44393
rect 105357 44384 105369 44387
rect 105219 44356 105369 44384
rect 105219 44353 105231 44356
rect 105173 44347 105231 44353
rect 105357 44353 105369 44356
rect 105403 44353 105415 44387
rect 105357 44347 105415 44353
rect 104529 44319 104587 44325
rect 104529 44316 104541 44319
rect 103756 44288 104541 44316
rect 103756 44276 103762 44288
rect 104529 44285 104541 44288
rect 104575 44285 104587 44319
rect 104529 44279 104587 44285
rect 104710 44140 104716 44192
rect 104768 44180 104774 44192
rect 104989 44183 105047 44189
rect 104989 44180 105001 44183
rect 104768 44152 105001 44180
rect 104768 44140 104774 44152
rect 104989 44149 105001 44152
rect 105035 44149 105047 44183
rect 104989 44143 105047 44149
rect 1104 44090 7912 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 7912 44090
rect 1104 44016 7912 44038
rect 104052 44090 108836 44112
rect 104052 44038 105922 44090
rect 105974 44038 105986 44090
rect 106038 44038 106050 44090
rect 106102 44038 106114 44090
rect 106166 44038 106178 44090
rect 106230 44038 108836 44090
rect 104052 44016 108836 44038
rect 1104 43546 7912 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 7912 43546
rect 1104 43472 7912 43494
rect 104052 43546 108836 43568
rect 104052 43494 106658 43546
rect 106710 43494 106722 43546
rect 106774 43494 106786 43546
rect 106838 43494 106850 43546
rect 106902 43494 106914 43546
rect 106966 43494 108836 43546
rect 104052 43472 108836 43494
rect 1104 43002 7912 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 7912 43002
rect 1104 42928 7912 42950
rect 104052 43002 108836 43024
rect 104052 42950 105922 43002
rect 105974 42950 105986 43002
rect 106038 42950 106050 43002
rect 106102 42950 106114 43002
rect 106166 42950 106178 43002
rect 106230 42950 108836 43002
rect 104052 42928 108836 42950
rect 1104 42458 7912 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 7912 42458
rect 1104 42384 7912 42406
rect 104052 42458 108836 42480
rect 104052 42406 106658 42458
rect 106710 42406 106722 42458
rect 106774 42406 106786 42458
rect 106838 42406 106850 42458
rect 106902 42406 106914 42458
rect 106966 42406 108836 42458
rect 104052 42384 108836 42406
rect 105078 42304 105084 42356
rect 105136 42304 105142 42356
rect 104250 42168 104256 42220
rect 104308 42208 104314 42220
rect 104437 42211 104495 42217
rect 104437 42208 104449 42211
rect 104308 42180 104449 42208
rect 104308 42168 104314 42180
rect 104437 42177 104449 42180
rect 104483 42177 104495 42211
rect 104437 42171 104495 42177
rect 1104 41914 7912 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 7912 41914
rect 1104 41840 7912 41862
rect 104052 41914 108836 41936
rect 104052 41862 105922 41914
rect 105974 41862 105986 41914
rect 106038 41862 106050 41914
rect 106102 41862 106114 41914
rect 106166 41862 106178 41914
rect 106230 41862 108836 41914
rect 104052 41840 108836 41862
rect 1581 41735 1639 41741
rect 1581 41701 1593 41735
rect 1627 41732 1639 41735
rect 5534 41732 5540 41744
rect 1627 41704 5540 41732
rect 1627 41701 1639 41704
rect 1581 41695 1639 41701
rect 5534 41692 5540 41704
rect 5592 41692 5598 41744
rect 1210 41556 1216 41608
rect 1268 41596 1274 41608
rect 1397 41599 1455 41605
rect 1397 41596 1409 41599
rect 1268 41568 1409 41596
rect 1268 41556 1274 41568
rect 1397 41565 1409 41568
rect 1443 41596 1455 41599
rect 1673 41599 1731 41605
rect 1673 41596 1685 41599
rect 1443 41568 1685 41596
rect 1443 41565 1455 41568
rect 1397 41559 1455 41565
rect 1673 41565 1685 41568
rect 1719 41565 1731 41599
rect 1673 41559 1731 41565
rect 1104 41370 7912 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 7912 41370
rect 1104 41296 7912 41318
rect 104052 41370 108836 41392
rect 104052 41318 106658 41370
rect 106710 41318 106722 41370
rect 106774 41318 106786 41370
rect 106838 41318 106850 41370
rect 106902 41318 106914 41370
rect 106966 41318 108836 41370
rect 104052 41296 108836 41318
rect 1104 40826 7912 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 7912 40826
rect 1104 40752 7912 40774
rect 104052 40826 108836 40848
rect 104052 40774 105922 40826
rect 105974 40774 105986 40826
rect 106038 40774 106050 40826
rect 106102 40774 106114 40826
rect 106166 40774 106178 40826
rect 106230 40774 108836 40826
rect 104052 40752 108836 40774
rect 1104 40282 7912 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 7912 40282
rect 1104 40208 7912 40230
rect 104052 40282 108836 40304
rect 104052 40230 106658 40282
rect 106710 40230 106722 40282
rect 106774 40230 106786 40282
rect 106838 40230 106850 40282
rect 106902 40230 106914 40282
rect 106966 40230 108836 40282
rect 104052 40208 108836 40230
rect 1581 40171 1639 40177
rect 1581 40137 1593 40171
rect 1627 40168 1639 40171
rect 5534 40168 5540 40180
rect 1627 40140 5540 40168
rect 1627 40137 1639 40140
rect 1581 40131 1639 40137
rect 5534 40128 5540 40140
rect 5592 40128 5598 40180
rect 1394 39992 1400 40044
rect 1452 40032 1458 40044
rect 1673 40035 1731 40041
rect 1673 40032 1685 40035
rect 1452 40004 1685 40032
rect 1452 39992 1458 40004
rect 1673 40001 1685 40004
rect 1719 40001 1731 40035
rect 1673 39995 1731 40001
rect 1104 39738 7912 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 7912 39738
rect 1104 39664 7912 39686
rect 104052 39738 108836 39760
rect 104052 39686 105922 39738
rect 105974 39686 105986 39738
rect 106038 39686 106050 39738
rect 106102 39686 106114 39738
rect 106166 39686 106178 39738
rect 106230 39686 108836 39738
rect 104052 39664 108836 39686
rect 1104 39194 7912 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 7912 39194
rect 1104 39120 7912 39142
rect 104052 39194 108836 39216
rect 104052 39142 106658 39194
rect 106710 39142 106722 39194
rect 106774 39142 106786 39194
rect 106838 39142 106850 39194
rect 106902 39142 106914 39194
rect 106966 39142 108836 39194
rect 104052 39120 108836 39142
rect 104342 38836 104348 38888
rect 104400 38876 104406 38888
rect 105354 38876 105360 38888
rect 104400 38848 105360 38876
rect 104400 38836 104406 38848
rect 105354 38836 105360 38848
rect 105412 38836 105418 38888
rect 1104 38650 7912 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 7912 38650
rect 1104 38576 7912 38598
rect 104052 38650 108836 38672
rect 104052 38598 105922 38650
rect 105974 38598 105986 38650
rect 106038 38598 106050 38650
rect 106102 38598 106114 38650
rect 106166 38598 106178 38650
rect 106230 38598 108836 38650
rect 104052 38576 108836 38598
rect 1581 38471 1639 38477
rect 1581 38437 1593 38471
rect 1627 38468 1639 38471
rect 8386 38468 8392 38480
rect 1627 38440 8392 38468
rect 1627 38437 1639 38440
rect 1581 38431 1639 38437
rect 8386 38428 8392 38440
rect 8444 38428 8450 38480
rect 1210 38292 1216 38344
rect 1268 38332 1274 38344
rect 1397 38335 1455 38341
rect 1397 38332 1409 38335
rect 1268 38304 1409 38332
rect 1268 38292 1274 38304
rect 1397 38301 1409 38304
rect 1443 38332 1455 38335
rect 1673 38335 1731 38341
rect 1673 38332 1685 38335
rect 1443 38304 1685 38332
rect 1443 38301 1455 38304
rect 1397 38295 1455 38301
rect 1673 38301 1685 38304
rect 1719 38301 1731 38335
rect 1673 38295 1731 38301
rect 1104 38106 7912 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 7912 38106
rect 1104 38032 7912 38054
rect 104052 38106 108836 38128
rect 104052 38054 106658 38106
rect 106710 38054 106722 38106
rect 106774 38054 106786 38106
rect 106838 38054 106850 38106
rect 106902 38054 106914 38106
rect 106966 38054 108836 38106
rect 104052 38032 108836 38054
rect 104250 37952 104256 38004
rect 104308 37992 104314 38004
rect 104345 37995 104403 38001
rect 104345 37992 104357 37995
rect 104308 37964 104357 37992
rect 104308 37952 104314 37964
rect 104345 37961 104357 37964
rect 104391 37961 104403 37995
rect 104345 37955 104403 37961
rect 105814 37952 105820 38004
rect 105872 37992 105878 38004
rect 106185 37995 106243 38001
rect 106185 37992 106197 37995
rect 105872 37964 106197 37992
rect 105872 37952 105878 37964
rect 104710 37816 104716 37868
rect 104768 37816 104774 37868
rect 106108 37865 106136 37964
rect 106185 37961 106197 37964
rect 106231 37961 106243 37995
rect 106185 37955 106243 37961
rect 106093 37859 106151 37865
rect 106093 37825 106105 37859
rect 106139 37825 106151 37859
rect 106093 37819 106151 37825
rect 105170 37748 105176 37800
rect 105228 37788 105234 37800
rect 105817 37791 105875 37797
rect 105817 37788 105829 37791
rect 105228 37760 105829 37788
rect 105228 37748 105234 37760
rect 105817 37757 105829 37760
rect 105863 37757 105875 37791
rect 105817 37751 105875 37757
rect 1104 37562 7912 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 7912 37562
rect 1104 37488 7912 37510
rect 104052 37562 108836 37584
rect 104052 37510 105922 37562
rect 105974 37510 105986 37562
rect 106038 37510 106050 37562
rect 106102 37510 106114 37562
rect 106166 37510 106178 37562
rect 106230 37510 108836 37562
rect 104052 37488 108836 37510
rect 104621 37315 104679 37321
rect 104621 37281 104633 37315
rect 104667 37312 104679 37315
rect 104710 37312 104716 37324
rect 104667 37284 104716 37312
rect 104667 37281 104679 37284
rect 104621 37275 104679 37281
rect 104710 37272 104716 37284
rect 104768 37272 104774 37324
rect 1394 37204 1400 37256
rect 1452 37244 1458 37256
rect 1673 37247 1731 37253
rect 1673 37244 1685 37247
rect 1452 37216 1685 37244
rect 1452 37204 1458 37216
rect 1673 37213 1685 37216
rect 1719 37213 1731 37247
rect 1673 37207 1731 37213
rect 104250 37204 104256 37256
rect 104308 37244 104314 37256
rect 104437 37247 104495 37253
rect 104437 37244 104449 37247
rect 104308 37216 104449 37244
rect 104308 37204 104314 37216
rect 104437 37213 104449 37216
rect 104483 37213 104495 37247
rect 104437 37207 104495 37213
rect 9490 37176 9496 37188
rect 1596 37148 9496 37176
rect 1596 37117 1624 37148
rect 9490 37136 9496 37148
rect 9548 37136 9554 37188
rect 1581 37111 1639 37117
rect 1581 37077 1593 37111
rect 1627 37077 1639 37111
rect 1581 37071 1639 37077
rect 1104 37018 7912 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 7912 37018
rect 1104 36944 7912 36966
rect 104052 37018 108836 37040
rect 104052 36966 106658 37018
rect 106710 36966 106722 37018
rect 106774 36966 106786 37018
rect 106838 36966 106850 37018
rect 106902 36966 106914 37018
rect 106966 36966 108836 37018
rect 104052 36944 108836 36966
rect 1104 36474 7912 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 7912 36474
rect 1104 36400 7912 36422
rect 104052 36474 108836 36496
rect 104052 36422 105922 36474
rect 105974 36422 105986 36474
rect 106038 36422 106050 36474
rect 106102 36422 106114 36474
rect 106166 36422 106178 36474
rect 106230 36422 108836 36474
rect 104052 36400 108836 36422
rect 1104 35930 7912 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 7912 35930
rect 1104 35856 7912 35878
rect 104052 35930 108836 35952
rect 104052 35878 106658 35930
rect 106710 35878 106722 35930
rect 106774 35878 106786 35930
rect 106838 35878 106850 35930
rect 106902 35878 106914 35930
rect 106966 35878 108836 35930
rect 104052 35856 108836 35878
rect 1581 35819 1639 35825
rect 1581 35785 1593 35819
rect 1627 35816 1639 35819
rect 9490 35816 9496 35828
rect 1627 35788 9496 35816
rect 1627 35785 1639 35788
rect 1581 35779 1639 35785
rect 9490 35776 9496 35788
rect 9548 35776 9554 35828
rect 1302 35640 1308 35692
rect 1360 35680 1366 35692
rect 1397 35683 1455 35689
rect 1397 35680 1409 35683
rect 1360 35652 1409 35680
rect 1360 35640 1366 35652
rect 1397 35649 1409 35652
rect 1443 35680 1455 35683
rect 1673 35683 1731 35689
rect 1673 35680 1685 35683
rect 1443 35652 1685 35680
rect 1443 35649 1455 35652
rect 1397 35643 1455 35649
rect 1673 35649 1685 35652
rect 1719 35649 1731 35683
rect 1673 35643 1731 35649
rect 1104 35386 7912 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 7912 35386
rect 1104 35312 7912 35334
rect 104052 35386 108836 35408
rect 104052 35334 105922 35386
rect 105974 35334 105986 35386
rect 106038 35334 106050 35386
rect 106102 35334 106114 35386
rect 106166 35334 106178 35386
rect 106230 35334 108836 35386
rect 104052 35312 108836 35334
rect 1104 34842 7912 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 7912 34842
rect 1104 34768 7912 34790
rect 104052 34842 108836 34864
rect 104052 34790 106658 34842
rect 106710 34790 106722 34842
rect 106774 34790 106786 34842
rect 106838 34790 106850 34842
rect 106902 34790 106914 34842
rect 106966 34790 108836 34842
rect 104052 34768 108836 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34728 1639 34731
rect 5534 34728 5540 34740
rect 1627 34700 5540 34728
rect 1627 34697 1639 34700
rect 1581 34691 1639 34697
rect 5534 34688 5540 34700
rect 5592 34688 5598 34740
rect 1394 34552 1400 34604
rect 1452 34592 1458 34604
rect 1673 34595 1731 34601
rect 1673 34592 1685 34595
rect 1452 34564 1685 34592
rect 1452 34552 1458 34564
rect 1673 34561 1685 34564
rect 1719 34561 1731 34595
rect 1673 34555 1731 34561
rect 1104 34298 7912 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 7912 34298
rect 1104 34224 7912 34246
rect 104052 34298 108836 34320
rect 104052 34246 105922 34298
rect 105974 34246 105986 34298
rect 106038 34246 106050 34298
rect 106102 34246 106114 34298
rect 106166 34246 106178 34298
rect 106230 34246 108836 34298
rect 104052 34224 108836 34246
rect 1104 33754 7912 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 7912 33754
rect 1104 33680 7912 33702
rect 104052 33754 108836 33776
rect 104052 33702 106658 33754
rect 106710 33702 106722 33754
rect 106774 33702 106786 33754
rect 106838 33702 106850 33754
rect 106902 33702 106914 33754
rect 106966 33702 108836 33754
rect 104052 33680 108836 33702
rect 1104 33210 7912 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 7912 33210
rect 1104 33136 7912 33158
rect 104052 33210 108836 33232
rect 104052 33158 105922 33210
rect 105974 33158 105986 33210
rect 106038 33158 106050 33210
rect 106102 33158 106114 33210
rect 106166 33158 106178 33210
rect 106230 33158 108836 33210
rect 104052 33136 108836 33158
rect 1104 32666 7912 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 7912 32666
rect 1104 32592 7912 32614
rect 104052 32666 108836 32688
rect 104052 32614 106658 32666
rect 106710 32614 106722 32666
rect 106774 32614 106786 32666
rect 106838 32614 106850 32666
rect 106902 32614 106914 32666
rect 106966 32614 108836 32666
rect 104052 32592 108836 32614
rect 1104 32122 7912 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 7912 32122
rect 1104 32048 7912 32070
rect 104052 32122 108836 32144
rect 104052 32070 105922 32122
rect 105974 32070 105986 32122
rect 106038 32070 106050 32122
rect 106102 32070 106114 32122
rect 106166 32070 106178 32122
rect 106230 32070 108836 32122
rect 104052 32048 108836 32070
rect 1104 31578 7912 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 7912 31578
rect 1104 31504 7912 31526
rect 104052 31578 108836 31600
rect 104052 31526 106658 31578
rect 106710 31526 106722 31578
rect 106774 31526 106786 31578
rect 106838 31526 106850 31578
rect 106902 31526 106914 31578
rect 106966 31526 108836 31578
rect 104052 31504 108836 31526
rect 1104 31034 7912 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 7912 31034
rect 1104 30960 7912 30982
rect 104052 31034 108836 31056
rect 104052 30982 105922 31034
rect 105974 30982 105986 31034
rect 106038 30982 106050 31034
rect 106102 30982 106114 31034
rect 106166 30982 106178 31034
rect 106230 30982 108836 31034
rect 104052 30960 108836 30982
rect 1104 30490 7912 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 7912 30490
rect 1104 30416 7912 30438
rect 104052 30490 108836 30512
rect 104052 30438 106658 30490
rect 106710 30438 106722 30490
rect 106774 30438 106786 30490
rect 106838 30438 106850 30490
rect 106902 30438 106914 30490
rect 106966 30438 108836 30490
rect 104052 30416 108836 30438
rect 1104 29946 7912 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 7912 29946
rect 1104 29872 7912 29894
rect 104052 29946 108836 29968
rect 104052 29894 105922 29946
rect 105974 29894 105986 29946
rect 106038 29894 106050 29946
rect 106102 29894 106114 29946
rect 106166 29894 106178 29946
rect 106230 29894 108836 29946
rect 104052 29872 108836 29894
rect 1104 29402 7912 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 7912 29402
rect 1104 29328 7912 29350
rect 104052 29402 108836 29424
rect 104052 29350 106658 29402
rect 106710 29350 106722 29402
rect 106774 29350 106786 29402
rect 106838 29350 106850 29402
rect 106902 29350 106914 29402
rect 106966 29350 108836 29402
rect 104052 29328 108836 29350
rect 1104 28858 7912 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 7912 28858
rect 1104 28784 7912 28806
rect 104052 28858 108836 28880
rect 104052 28806 105922 28858
rect 105974 28806 105986 28858
rect 106038 28806 106050 28858
rect 106102 28806 106114 28858
rect 106166 28806 106178 28858
rect 106230 28806 108836 28858
rect 104052 28784 108836 28806
rect 1104 28314 7912 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 7912 28314
rect 1104 28240 7912 28262
rect 104052 28314 108836 28336
rect 104052 28262 106658 28314
rect 106710 28262 106722 28314
rect 106774 28262 106786 28314
rect 106838 28262 106850 28314
rect 106902 28262 106914 28314
rect 106966 28262 108836 28314
rect 104052 28240 108836 28262
rect 1104 27770 7912 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 7912 27770
rect 1104 27696 7912 27718
rect 104052 27770 108836 27792
rect 104052 27718 105922 27770
rect 105974 27718 105986 27770
rect 106038 27718 106050 27770
rect 106102 27718 106114 27770
rect 106166 27718 106178 27770
rect 106230 27718 108836 27770
rect 104052 27696 108836 27718
rect 1104 27226 7912 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 7912 27226
rect 1104 27152 7912 27174
rect 104052 27226 108836 27248
rect 104052 27174 106658 27226
rect 106710 27174 106722 27226
rect 106774 27174 106786 27226
rect 106838 27174 106850 27226
rect 106902 27174 106914 27226
rect 106966 27174 108836 27226
rect 104052 27152 108836 27174
rect 1104 26682 7912 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 7912 26682
rect 1104 26608 7912 26630
rect 104052 26682 108836 26704
rect 104052 26630 105922 26682
rect 105974 26630 105986 26682
rect 106038 26630 106050 26682
rect 106102 26630 106114 26682
rect 106166 26630 106178 26682
rect 106230 26630 108836 26682
rect 104052 26608 108836 26630
rect 1104 26138 7912 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 7912 26138
rect 1104 26064 7912 26086
rect 104052 26138 108836 26160
rect 104052 26086 106658 26138
rect 106710 26086 106722 26138
rect 106774 26086 106786 26138
rect 106838 26086 106850 26138
rect 106902 26086 106914 26138
rect 106966 26086 108836 26138
rect 104052 26064 108836 26086
rect 1104 25594 7912 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 7912 25594
rect 1104 25520 7912 25542
rect 104052 25594 108836 25616
rect 104052 25542 105922 25594
rect 105974 25542 105986 25594
rect 106038 25542 106050 25594
rect 106102 25542 106114 25594
rect 106166 25542 106178 25594
rect 106230 25542 108836 25594
rect 104052 25520 108836 25542
rect 102594 25100 102600 25152
rect 102652 25140 102658 25152
rect 104345 25143 104403 25149
rect 104345 25140 104357 25143
rect 102652 25112 104357 25140
rect 102652 25100 102658 25112
rect 104345 25109 104357 25112
rect 104391 25109 104403 25143
rect 104345 25103 104403 25109
rect 1104 25050 7912 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 7912 25050
rect 1104 24976 7912 24998
rect 104052 25050 108836 25072
rect 104052 24998 106658 25050
rect 106710 24998 106722 25050
rect 106774 24998 106786 25050
rect 106838 24998 106850 25050
rect 106902 24998 106914 25050
rect 106966 24998 108836 25050
rect 104052 24976 108836 24998
rect 1104 24506 7912 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 7912 24506
rect 1104 24432 7912 24454
rect 104052 24506 108836 24528
rect 104052 24454 105922 24506
rect 105974 24454 105986 24506
rect 106038 24454 106050 24506
rect 106102 24454 106114 24506
rect 106166 24454 106178 24506
rect 106230 24454 108836 24506
rect 104052 24432 108836 24454
rect 1104 23962 7912 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 7912 23962
rect 1104 23888 7912 23910
rect 104052 23962 108836 23984
rect 104052 23910 106658 23962
rect 106710 23910 106722 23962
rect 106774 23910 106786 23962
rect 106838 23910 106850 23962
rect 106902 23910 106914 23962
rect 106966 23910 108836 23962
rect 104052 23888 108836 23910
rect 101950 23808 101956 23860
rect 102008 23848 102014 23860
rect 104345 23851 104403 23857
rect 104345 23848 104357 23851
rect 102008 23820 104357 23848
rect 102008 23808 102014 23820
rect 104345 23817 104357 23820
rect 104391 23817 104403 23851
rect 104345 23811 104403 23817
rect 1104 23418 7912 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 7912 23418
rect 1104 23344 7912 23366
rect 104052 23418 108836 23440
rect 104052 23366 105922 23418
rect 105974 23366 105986 23418
rect 106038 23366 106050 23418
rect 106102 23366 106114 23418
rect 106166 23366 106178 23418
rect 106230 23366 108836 23418
rect 104052 23344 108836 23366
rect 1104 22874 7912 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 7912 22874
rect 1104 22800 7912 22822
rect 104052 22874 108836 22896
rect 104052 22822 106658 22874
rect 106710 22822 106722 22874
rect 106774 22822 106786 22874
rect 106838 22822 106850 22874
rect 106902 22822 106914 22874
rect 106966 22822 108836 22874
rect 104052 22800 108836 22822
rect 104342 22720 104348 22772
rect 104400 22720 104406 22772
rect 1104 22330 7912 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 7912 22330
rect 1104 22256 7912 22278
rect 104052 22330 108836 22352
rect 104052 22278 105922 22330
rect 105974 22278 105986 22330
rect 106038 22278 106050 22330
rect 106102 22278 106114 22330
rect 106166 22278 106178 22330
rect 106230 22278 108836 22330
rect 104052 22256 108836 22278
rect 1104 21786 7912 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 7912 21786
rect 1104 21712 7912 21734
rect 104052 21786 108836 21808
rect 104052 21734 106658 21786
rect 106710 21734 106722 21786
rect 106774 21734 106786 21786
rect 106838 21734 106850 21786
rect 106902 21734 106914 21786
rect 106966 21734 108836 21786
rect 104052 21712 108836 21734
rect 1104 21242 7912 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 7912 21242
rect 1104 21168 7912 21190
rect 104052 21242 108836 21264
rect 104052 21190 105922 21242
rect 105974 21190 105986 21242
rect 106038 21190 106050 21242
rect 106102 21190 106114 21242
rect 106166 21190 106178 21242
rect 106230 21190 108836 21242
rect 104052 21168 108836 21190
rect 1104 20698 7912 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 7912 20698
rect 1104 20624 7912 20646
rect 104052 20698 108836 20720
rect 104052 20646 106658 20698
rect 106710 20646 106722 20698
rect 106774 20646 106786 20698
rect 106838 20646 106850 20698
rect 106902 20646 106914 20698
rect 106966 20646 108836 20698
rect 104052 20624 108836 20646
rect 1104 20154 7912 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 7912 20154
rect 1104 20080 7912 20102
rect 104052 20154 108836 20176
rect 104052 20102 105922 20154
rect 105974 20102 105986 20154
rect 106038 20102 106050 20154
rect 106102 20102 106114 20154
rect 106166 20102 106178 20154
rect 106230 20102 108836 20154
rect 104052 20080 108836 20102
rect 1104 19610 7912 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 7912 19610
rect 1104 19536 7912 19558
rect 104052 19610 108836 19632
rect 104052 19558 106658 19610
rect 106710 19558 106722 19610
rect 106774 19558 106786 19610
rect 106838 19558 106850 19610
rect 106902 19558 106914 19610
rect 106966 19558 108836 19610
rect 104052 19536 108836 19558
rect 1104 19066 7912 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 7912 19066
rect 1104 18992 7912 19014
rect 104052 19066 108836 19088
rect 104052 19014 105922 19066
rect 105974 19014 105986 19066
rect 106038 19014 106050 19066
rect 106102 19014 106114 19066
rect 106166 19014 106178 19066
rect 106230 19014 108836 19066
rect 104052 18992 108836 19014
rect 1104 18522 7912 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 7912 18522
rect 1104 18448 7912 18470
rect 104052 18522 108836 18544
rect 104052 18470 106658 18522
rect 106710 18470 106722 18522
rect 106774 18470 106786 18522
rect 106838 18470 106850 18522
rect 106902 18470 106914 18522
rect 106966 18470 108836 18522
rect 104052 18448 108836 18470
rect 1104 17978 7912 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 7912 17978
rect 1104 17904 7912 17926
rect 104052 17978 108836 18000
rect 104052 17926 105922 17978
rect 105974 17926 105986 17978
rect 106038 17926 106050 17978
rect 106102 17926 106114 17978
rect 106166 17926 106178 17978
rect 106230 17926 108836 17978
rect 104052 17904 108836 17926
rect 1104 17434 7912 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 7912 17434
rect 1104 17360 7912 17382
rect 104052 17434 108836 17456
rect 104052 17382 106658 17434
rect 106710 17382 106722 17434
rect 106774 17382 106786 17434
rect 106838 17382 106850 17434
rect 106902 17382 106914 17434
rect 106966 17382 108836 17434
rect 104052 17360 108836 17382
rect 1104 16890 7912 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 7912 16890
rect 1104 16816 7912 16838
rect 104052 16890 108836 16912
rect 104052 16838 105922 16890
rect 105974 16838 105986 16890
rect 106038 16838 106050 16890
rect 106102 16838 106114 16890
rect 106166 16838 106178 16890
rect 106230 16838 108836 16890
rect 104052 16816 108836 16838
rect 1104 16346 7912 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 7912 16346
rect 1104 16272 7912 16294
rect 104052 16346 108836 16368
rect 104052 16294 106658 16346
rect 106710 16294 106722 16346
rect 106774 16294 106786 16346
rect 106838 16294 106850 16346
rect 106902 16294 106914 16346
rect 106966 16294 108836 16346
rect 104052 16272 108836 16294
rect 1302 16056 1308 16108
rect 1360 16096 1366 16108
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 1360 16068 1409 16096
rect 1360 16056 1366 16068
rect 1397 16065 1409 16068
rect 1443 16096 1455 16099
rect 1673 16099 1731 16105
rect 1673 16096 1685 16099
rect 1443 16068 1685 16096
rect 1443 16065 1455 16068
rect 1397 16059 1455 16065
rect 1673 16065 1685 16068
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 9490 15960 9496 15972
rect 1627 15932 9496 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 9490 15920 9496 15932
rect 9548 15920 9554 15972
rect 1104 15802 7912 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 7912 15802
rect 1104 15728 7912 15750
rect 104052 15802 108836 15824
rect 104052 15750 105922 15802
rect 105974 15750 105986 15802
rect 106038 15750 106050 15802
rect 106102 15750 106114 15802
rect 106166 15750 106178 15802
rect 106230 15750 108836 15802
rect 104052 15728 108836 15750
rect 1104 15258 7912 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 7912 15258
rect 1104 15184 7912 15206
rect 104052 15258 108836 15280
rect 104052 15206 106658 15258
rect 106710 15206 106722 15258
rect 106774 15206 106786 15258
rect 106838 15206 106850 15258
rect 106902 15206 106914 15258
rect 106966 15206 108836 15258
rect 104052 15184 108836 15206
rect 1104 14714 7912 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 7912 14714
rect 1104 14640 7912 14662
rect 104052 14714 108836 14736
rect 104052 14662 105922 14714
rect 105974 14662 105986 14714
rect 106038 14662 106050 14714
rect 106102 14662 106114 14714
rect 106166 14662 106178 14714
rect 106230 14662 108836 14714
rect 104052 14640 108836 14662
rect 1104 14170 7912 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 7912 14170
rect 1104 14096 7912 14118
rect 104052 14170 108836 14192
rect 104052 14118 106658 14170
rect 106710 14118 106722 14170
rect 106774 14118 106786 14170
rect 106838 14118 106850 14170
rect 106902 14118 106914 14170
rect 106966 14118 108836 14170
rect 104052 14096 108836 14118
rect 1104 13626 7912 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 7912 13626
rect 1104 13552 7912 13574
rect 104052 13626 108836 13648
rect 104052 13574 105922 13626
rect 105974 13574 105986 13626
rect 106038 13574 106050 13626
rect 106102 13574 106114 13626
rect 106166 13574 106178 13626
rect 106230 13574 108836 13626
rect 104052 13552 108836 13574
rect 1104 13082 7912 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 7912 13082
rect 1104 13008 7912 13030
rect 104052 13082 108836 13104
rect 104052 13030 106658 13082
rect 106710 13030 106722 13082
rect 106774 13030 106786 13082
rect 106838 13030 106850 13082
rect 106902 13030 106914 13082
rect 106966 13030 108836 13082
rect 104052 13008 108836 13030
rect 1104 12538 7912 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 7912 12538
rect 1104 12464 7912 12486
rect 104052 12538 108836 12560
rect 104052 12486 105922 12538
rect 105974 12486 105986 12538
rect 106038 12486 106050 12538
rect 106102 12486 106114 12538
rect 106166 12486 106178 12538
rect 106230 12486 108836 12538
rect 104052 12464 108836 12486
rect 1104 11994 7912 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 7912 11994
rect 1104 11920 7912 11942
rect 104052 11994 108836 12016
rect 104052 11942 106658 11994
rect 106710 11942 106722 11994
rect 106774 11942 106786 11994
rect 106838 11942 106850 11994
rect 106902 11942 106914 11994
rect 106966 11942 108836 11994
rect 104052 11920 108836 11942
rect 1104 11450 7912 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 7912 11450
rect 1104 11376 7912 11398
rect 104052 11450 108836 11472
rect 104052 11398 105922 11450
rect 105974 11398 105986 11450
rect 106038 11398 106050 11450
rect 106102 11398 106114 11450
rect 106166 11398 106178 11450
rect 106230 11398 108836 11450
rect 104052 11376 108836 11398
rect 1104 10906 7912 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 7912 10906
rect 1104 10832 7912 10854
rect 104052 10906 108836 10928
rect 104052 10854 106658 10906
rect 106710 10854 106722 10906
rect 106774 10854 106786 10906
rect 106838 10854 106850 10906
rect 106902 10854 106914 10906
rect 106966 10854 108836 10906
rect 104052 10832 108836 10854
rect 1104 10362 7912 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 7912 10362
rect 1104 10288 7912 10310
rect 104052 10362 108836 10384
rect 104052 10310 105922 10362
rect 105974 10310 105986 10362
rect 106038 10310 106050 10362
rect 106102 10310 106114 10362
rect 106166 10310 106178 10362
rect 106230 10310 108836 10362
rect 104052 10288 108836 10310
rect 90726 10004 90732 10056
rect 90784 10044 90790 10056
rect 104710 10044 104716 10056
rect 90784 10016 104716 10044
rect 90784 10004 90790 10016
rect 104710 10004 104716 10016
rect 104768 10004 104774 10056
rect 90818 9936 90824 9988
rect 90876 9976 90882 9988
rect 103790 9976 103796 9988
rect 90876 9948 103796 9976
rect 90876 9936 90882 9948
rect 103790 9936 103796 9948
rect 103848 9936 103854 9988
rect 1104 9818 7912 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 7912 9818
rect 1104 9744 7912 9766
rect 104052 9818 108836 9840
rect 104052 9766 106658 9818
rect 106710 9766 106722 9818
rect 106774 9766 106786 9818
rect 106838 9766 106850 9818
rect 106902 9766 106914 9818
rect 106966 9766 108836 9818
rect 104052 9744 108836 9766
rect 1104 9274 7912 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 7912 9274
rect 1104 9200 7912 9222
rect 104052 9274 108836 9296
rect 104052 9222 105922 9274
rect 105974 9222 105986 9274
rect 106038 9222 106050 9274
rect 106102 9222 106114 9274
rect 106166 9222 106178 9274
rect 106230 9222 108836 9274
rect 104052 9200 108836 9222
rect 1104 8730 7912 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 7912 8730
rect 1104 8656 7912 8678
rect 104052 8730 108836 8752
rect 104052 8678 106658 8730
rect 106710 8678 106722 8730
rect 106774 8678 106786 8730
rect 106838 8678 106850 8730
rect 106902 8678 106914 8730
rect 106966 8678 108836 8730
rect 104052 8656 108836 8678
rect 1104 8186 7912 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 7912 8186
rect 1104 8112 7912 8134
rect 104052 8186 108836 8208
rect 104052 8134 105922 8186
rect 105974 8134 105986 8186
rect 106038 8134 106050 8186
rect 106102 8134 106114 8186
rect 106166 8134 106178 8186
rect 106230 8134 108836 8186
rect 104052 8112 108836 8134
rect 1104 7642 108836 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 66314 7642
rect 66366 7590 66378 7642
rect 66430 7590 66442 7642
rect 66494 7590 66506 7642
rect 66558 7590 66570 7642
rect 66622 7590 97034 7642
rect 97086 7590 97098 7642
rect 97150 7590 97162 7642
rect 97214 7590 97226 7642
rect 97278 7590 97290 7642
rect 97342 7590 106658 7642
rect 106710 7590 106722 7642
rect 106774 7590 106786 7642
rect 106838 7590 106850 7642
rect 106902 7590 106914 7642
rect 106966 7590 108836 7642
rect 1104 7568 108836 7590
rect 16114 7488 16120 7540
rect 16172 7488 16178 7540
rect 90634 7488 90640 7540
rect 90692 7488 90698 7540
rect 90726 7488 90732 7540
rect 90784 7488 90790 7540
rect 91002 7488 91008 7540
rect 91060 7488 91066 7540
rect 1104 7098 108836 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 96374 7098
rect 96426 7046 96438 7098
rect 96490 7046 96502 7098
rect 96554 7046 96566 7098
rect 96618 7046 96630 7098
rect 96682 7046 105922 7098
rect 105974 7046 105986 7098
rect 106038 7046 106050 7098
rect 106102 7046 106114 7098
rect 106166 7046 106178 7098
rect 106230 7046 108836 7098
rect 1104 7024 108836 7046
rect 1104 6554 108836 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 66314 6554
rect 66366 6502 66378 6554
rect 66430 6502 66442 6554
rect 66494 6502 66506 6554
rect 66558 6502 66570 6554
rect 66622 6502 97034 6554
rect 97086 6502 97098 6554
rect 97150 6502 97162 6554
rect 97214 6502 97226 6554
rect 97278 6502 97290 6554
rect 97342 6502 108836 6554
rect 1104 6480 108836 6502
rect 1104 6010 108836 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 96374 6010
rect 96426 5958 96438 6010
rect 96490 5958 96502 6010
rect 96554 5958 96566 6010
rect 96618 5958 96630 6010
rect 96682 5958 108836 6010
rect 1104 5936 108836 5958
rect 1104 5466 108836 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 66314 5466
rect 66366 5414 66378 5466
rect 66430 5414 66442 5466
rect 66494 5414 66506 5466
rect 66558 5414 66570 5466
rect 66622 5414 97034 5466
rect 97086 5414 97098 5466
rect 97150 5414 97162 5466
rect 97214 5414 97226 5466
rect 97278 5414 97290 5466
rect 97342 5414 108836 5466
rect 1104 5392 108836 5414
rect 1104 4922 108836 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 96374 4922
rect 96426 4870 96438 4922
rect 96490 4870 96502 4922
rect 96554 4870 96566 4922
rect 96618 4870 96630 4922
rect 96682 4870 108836 4922
rect 1104 4848 108836 4870
rect 1104 4378 108836 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 66314 4378
rect 66366 4326 66378 4378
rect 66430 4326 66442 4378
rect 66494 4326 66506 4378
rect 66558 4326 66570 4378
rect 66622 4326 97034 4378
rect 97086 4326 97098 4378
rect 97150 4326 97162 4378
rect 97214 4326 97226 4378
rect 97278 4326 97290 4378
rect 97342 4326 108836 4378
rect 1104 4304 108836 4326
rect 1104 3834 108836 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 96374 3834
rect 96426 3782 96438 3834
rect 96490 3782 96502 3834
rect 96554 3782 96566 3834
rect 96618 3782 96630 3834
rect 96682 3782 108836 3834
rect 1104 3760 108836 3782
rect 1104 3290 108836 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 66314 3290
rect 66366 3238 66378 3290
rect 66430 3238 66442 3290
rect 66494 3238 66506 3290
rect 66558 3238 66570 3290
rect 66622 3238 97034 3290
rect 97086 3238 97098 3290
rect 97150 3238 97162 3290
rect 97214 3238 97226 3290
rect 97278 3238 97290 3290
rect 97342 3238 108836 3290
rect 1104 3216 108836 3238
rect 1104 2746 108836 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 96374 2746
rect 96426 2694 96438 2746
rect 96490 2694 96502 2746
rect 96554 2694 96566 2746
rect 96618 2694 96630 2746
rect 96682 2694 108836 2746
rect 1104 2672 108836 2694
rect 23474 2592 23480 2644
rect 23532 2592 23538 2644
rect 24762 2592 24768 2644
rect 24820 2592 24826 2644
rect 25866 2592 25872 2644
rect 25924 2592 25930 2644
rect 27154 2592 27160 2644
rect 27212 2592 27218 2644
rect 28442 2592 28448 2644
rect 28500 2592 28506 2644
rect 29270 2592 29276 2644
rect 29328 2592 29334 2644
rect 30558 2592 30564 2644
rect 30616 2592 30622 2644
rect 31662 2592 31668 2644
rect 31720 2592 31726 2644
rect 32950 2592 32956 2644
rect 33008 2592 33014 2644
rect 34238 2592 34244 2644
rect 34296 2592 34302 2644
rect 35434 2592 35440 2644
rect 35492 2632 35498 2644
rect 35529 2635 35587 2641
rect 35529 2632 35541 2635
rect 35492 2604 35541 2632
rect 35492 2592 35498 2604
rect 35529 2601 35541 2604
rect 35575 2601 35587 2635
rect 35529 2595 35587 2601
rect 36354 2592 36360 2644
rect 36412 2592 36418 2644
rect 37458 2592 37464 2644
rect 37516 2592 37522 2644
rect 38746 2592 38752 2644
rect 38804 2592 38810 2644
rect 39942 2592 39948 2644
rect 40000 2632 40006 2644
rect 40037 2635 40095 2641
rect 40037 2632 40049 2635
rect 40000 2604 40049 2632
rect 40000 2592 40006 2604
rect 40037 2601 40049 2604
rect 40083 2601 40095 2635
rect 40037 2595 40095 2601
rect 41322 2592 41328 2644
rect 41380 2592 41386 2644
rect 42150 2592 42156 2644
rect 42208 2592 42214 2644
rect 43438 2592 43444 2644
rect 43496 2592 43502 2644
rect 23293 2431 23351 2437
rect 23293 2428 23305 2431
rect 23216 2400 23305 2428
rect 23216 2304 23244 2400
rect 23293 2397 23305 2400
rect 23339 2397 23351 2431
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23293 2391 23351 2397
rect 24504 2400 24593 2428
rect 24504 2304 24532 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 24581 2391 24639 2397
rect 25792 2400 26065 2428
rect 25792 2304 25820 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 26053 2391 26111 2397
rect 27080 2400 27353 2428
rect 27080 2304 27108 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 28629 2431 28687 2437
rect 28629 2428 28641 2431
rect 27341 2391 27399 2397
rect 28368 2400 28641 2428
rect 28368 2304 28396 2400
rect 28629 2397 28641 2400
rect 28675 2397 28687 2431
rect 29089 2431 29147 2437
rect 29089 2428 29101 2431
rect 28629 2391 28687 2397
rect 29012 2400 29101 2428
rect 29012 2304 29040 2400
rect 29089 2397 29101 2400
rect 29135 2397 29147 2431
rect 30377 2431 30435 2437
rect 30377 2428 30389 2431
rect 29089 2391 29147 2397
rect 30300 2400 30389 2428
rect 30300 2304 30328 2400
rect 30377 2397 30389 2400
rect 30423 2397 30435 2431
rect 31849 2431 31907 2437
rect 31849 2428 31861 2431
rect 30377 2391 30435 2397
rect 31588 2400 31861 2428
rect 31588 2304 31616 2400
rect 31849 2397 31861 2400
rect 31895 2397 31907 2431
rect 33137 2431 33195 2437
rect 33137 2428 33149 2431
rect 31849 2391 31907 2397
rect 32876 2400 33149 2428
rect 32876 2304 32904 2400
rect 33137 2397 33149 2400
rect 33183 2397 33195 2431
rect 34425 2431 34483 2437
rect 34425 2428 34437 2431
rect 33137 2391 33195 2397
rect 34164 2400 34437 2428
rect 34164 2304 34192 2400
rect 34425 2397 34437 2400
rect 34471 2397 34483 2431
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 34425 2391 34483 2397
rect 35452 2400 35725 2428
rect 35452 2304 35480 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 35713 2391 35771 2397
rect 36096 2400 36185 2428
rect 36096 2304 36124 2400
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 37645 2431 37703 2437
rect 37645 2428 37657 2431
rect 36173 2391 36231 2397
rect 37384 2400 37657 2428
rect 37384 2304 37412 2400
rect 37645 2397 37657 2400
rect 37691 2397 37703 2431
rect 38933 2431 38991 2437
rect 38933 2428 38945 2431
rect 37645 2391 37703 2397
rect 38672 2400 38945 2428
rect 38672 2304 38700 2400
rect 38933 2397 38945 2400
rect 38979 2397 38991 2431
rect 40221 2431 40279 2437
rect 40221 2428 40233 2431
rect 38933 2391 38991 2397
rect 39960 2400 40233 2428
rect 39960 2304 39988 2400
rect 40221 2397 40233 2400
rect 40267 2397 40279 2431
rect 41509 2431 41567 2437
rect 41509 2428 41521 2431
rect 40221 2391 40279 2397
rect 41248 2400 41521 2428
rect 41248 2304 41276 2400
rect 41509 2397 41521 2400
rect 41555 2397 41567 2431
rect 41969 2431 42027 2437
rect 41969 2428 41981 2431
rect 41509 2391 41567 2397
rect 41892 2400 41981 2428
rect 41892 2304 41920 2400
rect 41969 2397 41981 2400
rect 42015 2397 42027 2431
rect 43257 2431 43315 2437
rect 43257 2428 43269 2431
rect 41969 2391 42027 2397
rect 43180 2400 43269 2428
rect 43180 2304 43208 2400
rect 43257 2397 43269 2400
rect 43303 2397 43315 2431
rect 43257 2391 43315 2397
rect 23198 2252 23204 2304
rect 23256 2252 23262 2304
rect 24486 2252 24492 2304
rect 24544 2252 24550 2304
rect 25774 2252 25780 2304
rect 25832 2252 25838 2304
rect 27062 2252 27068 2304
rect 27120 2252 27126 2304
rect 28350 2252 28356 2304
rect 28408 2252 28414 2304
rect 28994 2252 29000 2304
rect 29052 2252 29058 2304
rect 30282 2252 30288 2304
rect 30340 2252 30346 2304
rect 31570 2252 31576 2304
rect 31628 2252 31634 2304
rect 32858 2252 32864 2304
rect 32916 2252 32922 2304
rect 34146 2252 34152 2304
rect 34204 2252 34210 2304
rect 35434 2252 35440 2304
rect 35492 2252 35498 2304
rect 36078 2252 36084 2304
rect 36136 2252 36142 2304
rect 37366 2252 37372 2304
rect 37424 2252 37430 2304
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 39942 2252 39948 2304
rect 40000 2252 40006 2304
rect 41230 2252 41236 2304
rect 41288 2252 41294 2304
rect 41874 2252 41880 2304
rect 41932 2252 41938 2304
rect 43162 2252 43168 2304
rect 43220 2252 43226 2304
rect 1104 2202 108836 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 66314 2202
rect 66366 2150 66378 2202
rect 66430 2150 66442 2202
rect 66494 2150 66506 2202
rect 66558 2150 66570 2202
rect 66622 2150 97034 2202
rect 97086 2150 97098 2202
rect 97150 2150 97162 2202
rect 97214 2150 97226 2202
rect 97278 2150 97290 2202
rect 97342 2150 108836 2202
rect 1104 2128 108836 2150
<< via1 >>
rect 98552 128324 98604 128376
rect 102140 128324 102192 128376
rect 4874 127270 4926 127322
rect 4938 127270 4990 127322
rect 5002 127270 5054 127322
rect 5066 127270 5118 127322
rect 5130 127270 5182 127322
rect 35594 127270 35646 127322
rect 35658 127270 35710 127322
rect 35722 127270 35774 127322
rect 35786 127270 35838 127322
rect 35850 127270 35902 127322
rect 66314 127270 66366 127322
rect 66378 127270 66430 127322
rect 66442 127270 66494 127322
rect 66506 127270 66558 127322
rect 66570 127270 66622 127322
rect 97034 127270 97086 127322
rect 97098 127270 97150 127322
rect 97162 127270 97214 127322
rect 97226 127270 97278 127322
rect 97290 127270 97342 127322
rect 4214 126726 4266 126778
rect 4278 126726 4330 126778
rect 4342 126726 4394 126778
rect 4406 126726 4458 126778
rect 4470 126726 4522 126778
rect 34934 126726 34986 126778
rect 34998 126726 35050 126778
rect 35062 126726 35114 126778
rect 35126 126726 35178 126778
rect 35190 126726 35242 126778
rect 65654 126726 65706 126778
rect 65718 126726 65770 126778
rect 65782 126726 65834 126778
rect 65846 126726 65898 126778
rect 65910 126726 65962 126778
rect 96374 126726 96426 126778
rect 96438 126726 96490 126778
rect 96502 126726 96554 126778
rect 96566 126726 96618 126778
rect 96630 126726 96682 126778
rect 105922 126726 105974 126778
rect 105986 126726 106038 126778
rect 106050 126726 106102 126778
rect 106114 126726 106166 126778
rect 106178 126726 106230 126778
rect 36084 126395 36136 126404
rect 36084 126361 36093 126395
rect 36093 126361 36127 126395
rect 36127 126361 36136 126395
rect 36084 126352 36136 126361
rect 36268 126395 36320 126404
rect 36268 126361 36277 126395
rect 36277 126361 36311 126395
rect 36311 126361 36320 126395
rect 36268 126352 36320 126361
rect 37740 126395 37792 126404
rect 37740 126361 37749 126395
rect 37749 126361 37783 126395
rect 37783 126361 37792 126395
rect 37740 126352 37792 126361
rect 42340 126420 42392 126472
rect 102600 126420 102652 126472
rect 41328 126395 41380 126404
rect 41328 126361 41337 126395
rect 41337 126361 41371 126395
rect 41371 126361 41380 126395
rect 41328 126352 41380 126361
rect 45192 126395 45244 126404
rect 45192 126361 45201 126395
rect 45201 126361 45235 126395
rect 45235 126361 45244 126395
rect 45192 126352 45244 126361
rect 48504 126395 48556 126404
rect 48504 126361 48513 126395
rect 48513 126361 48547 126395
rect 48547 126361 48556 126395
rect 48504 126352 48556 126361
rect 49700 126395 49752 126404
rect 49700 126361 49709 126395
rect 49709 126361 49743 126395
rect 49743 126361 49752 126395
rect 49700 126352 49752 126361
rect 56784 126352 56836 126404
rect 59360 126395 59412 126404
rect 59360 126361 59369 126395
rect 59369 126361 59403 126395
rect 59403 126361 59412 126395
rect 59360 126352 59412 126361
rect 61844 126395 61896 126404
rect 61844 126361 61853 126395
rect 61853 126361 61887 126395
rect 61887 126361 61896 126395
rect 61844 126352 61896 126361
rect 63960 126395 64012 126404
rect 63960 126361 63969 126395
rect 63969 126361 64003 126395
rect 64003 126361 64012 126395
rect 63960 126352 64012 126361
rect 64420 126352 64472 126404
rect 66076 126352 66128 126404
rect 68560 126352 68612 126404
rect 71412 126395 71464 126404
rect 71412 126361 71421 126395
rect 71421 126361 71455 126395
rect 71455 126361 71464 126395
rect 71412 126352 71464 126361
rect 77300 126395 77352 126404
rect 77300 126361 77309 126395
rect 77309 126361 77343 126395
rect 77343 126361 77352 126395
rect 77300 126352 77352 126361
rect 102324 126352 102376 126404
rect 37648 126327 37700 126336
rect 37648 126293 37657 126327
rect 37657 126293 37691 126327
rect 37691 126293 37700 126327
rect 37648 126284 37700 126293
rect 40960 126327 41012 126336
rect 40960 126293 40969 126327
rect 40969 126293 41003 126327
rect 41003 126293 41012 126327
rect 40960 126284 41012 126293
rect 41420 126327 41472 126336
rect 41420 126293 41429 126327
rect 41429 126293 41463 126327
rect 41463 126293 41472 126327
rect 41420 126284 41472 126293
rect 45100 126327 45152 126336
rect 45100 126293 45109 126327
rect 45109 126293 45143 126327
rect 45143 126293 45152 126327
rect 45100 126284 45152 126293
rect 48412 126327 48464 126336
rect 48412 126293 48421 126327
rect 48421 126293 48455 126327
rect 48455 126293 48464 126327
rect 48412 126284 48464 126293
rect 49608 126327 49660 126336
rect 49608 126293 49617 126327
rect 49617 126293 49651 126327
rect 49651 126293 49660 126327
rect 49608 126284 49660 126293
rect 59728 126327 59780 126336
rect 59728 126293 59737 126327
rect 59737 126293 59771 126327
rect 59771 126293 59780 126327
rect 59728 126284 59780 126293
rect 62212 126327 62264 126336
rect 62212 126293 62221 126327
rect 62221 126293 62255 126327
rect 62255 126293 62264 126327
rect 62212 126284 62264 126293
rect 64328 126327 64380 126336
rect 64328 126293 64337 126327
rect 64337 126293 64371 126327
rect 64371 126293 64380 126327
rect 64328 126284 64380 126293
rect 65984 126327 66036 126336
rect 65984 126293 65993 126327
rect 65993 126293 66027 126327
rect 66027 126293 66036 126327
rect 65984 126284 66036 126293
rect 67088 126327 67140 126336
rect 67088 126293 67097 126327
rect 67097 126293 67131 126327
rect 67131 126293 67140 126327
rect 67088 126284 67140 126293
rect 70860 126327 70912 126336
rect 70860 126293 70869 126327
rect 70869 126293 70903 126327
rect 70903 126293 70912 126327
rect 70860 126284 70912 126293
rect 71780 126327 71832 126336
rect 71780 126293 71789 126327
rect 71789 126293 71823 126327
rect 71823 126293 71832 126327
rect 71780 126284 71832 126293
rect 86316 126327 86368 126336
rect 86316 126293 86325 126327
rect 86325 126293 86359 126327
rect 86359 126293 86368 126327
rect 86316 126284 86368 126293
rect 87328 126327 87380 126336
rect 87328 126293 87337 126327
rect 87337 126293 87371 126327
rect 87371 126293 87380 126327
rect 87328 126284 87380 126293
rect 96068 126284 96120 126336
rect 4874 126182 4926 126234
rect 4938 126182 4990 126234
rect 5002 126182 5054 126234
rect 5066 126182 5118 126234
rect 5130 126182 5182 126234
rect 35594 126182 35646 126234
rect 35658 126182 35710 126234
rect 35722 126182 35774 126234
rect 35786 126182 35838 126234
rect 35850 126182 35902 126234
rect 66314 126182 66366 126234
rect 66378 126182 66430 126234
rect 66442 126182 66494 126234
rect 66506 126182 66558 126234
rect 66570 126182 66622 126234
rect 97034 126182 97086 126234
rect 97098 126182 97150 126234
rect 97162 126182 97214 126234
rect 97226 126182 97278 126234
rect 97290 126182 97342 126234
rect 106658 126182 106710 126234
rect 106722 126182 106774 126234
rect 106786 126182 106838 126234
rect 106850 126182 106902 126234
rect 106914 126182 106966 126234
rect 9588 126080 9640 126132
rect 49608 126080 49660 126132
rect 59728 126080 59780 126132
rect 103520 126080 103572 126132
rect 8208 126012 8260 126064
rect 45100 126012 45152 126064
rect 62212 126012 62264 126064
rect 102416 126012 102468 126064
rect 8116 125944 8168 125996
rect 41420 125944 41472 125996
rect 64328 125944 64380 125996
rect 102692 125944 102744 125996
rect 7932 125876 7984 125928
rect 40960 125876 41012 125928
rect 65984 125876 66036 125928
rect 103612 125876 103664 125928
rect 7840 125808 7892 125860
rect 37648 125808 37700 125860
rect 67088 125808 67140 125860
rect 102508 125808 102560 125860
rect 9496 125740 9548 125792
rect 36268 125740 36320 125792
rect 71780 125740 71832 125792
rect 103704 125740 103756 125792
rect 4214 125638 4266 125690
rect 4278 125638 4330 125690
rect 4342 125638 4394 125690
rect 4406 125638 4458 125690
rect 4470 125638 4522 125690
rect 8024 125672 8076 125724
rect 48412 125672 48464 125724
rect 70860 125672 70912 125724
rect 102232 125672 102284 125724
rect 105922 125638 105974 125690
rect 105986 125638 106038 125690
rect 106050 125638 106102 125690
rect 106114 125638 106166 125690
rect 106178 125638 106230 125690
rect 4874 125094 4926 125146
rect 4938 125094 4990 125146
rect 5002 125094 5054 125146
rect 5066 125094 5118 125146
rect 5130 125094 5182 125146
rect 106658 125094 106710 125146
rect 106722 125094 106774 125146
rect 106786 125094 106838 125146
rect 106850 125094 106902 125146
rect 106914 125094 106966 125146
rect 4214 124550 4266 124602
rect 4278 124550 4330 124602
rect 4342 124550 4394 124602
rect 4406 124550 4458 124602
rect 4470 124550 4522 124602
rect 105922 124550 105974 124602
rect 105986 124550 106038 124602
rect 106050 124550 106102 124602
rect 106114 124550 106166 124602
rect 106178 124550 106230 124602
rect 4874 124006 4926 124058
rect 4938 124006 4990 124058
rect 5002 124006 5054 124058
rect 5066 124006 5118 124058
rect 5130 124006 5182 124058
rect 106658 124006 106710 124058
rect 106722 124006 106774 124058
rect 106786 124006 106838 124058
rect 106850 124006 106902 124058
rect 106914 124006 106966 124058
rect 87328 123700 87380 123752
rect 104440 123700 104492 123752
rect 4214 123462 4266 123514
rect 4278 123462 4330 123514
rect 4342 123462 4394 123514
rect 4406 123462 4458 123514
rect 4470 123462 4522 123514
rect 105922 123462 105974 123514
rect 105986 123462 106038 123514
rect 106050 123462 106102 123514
rect 106114 123462 106166 123514
rect 106178 123462 106230 123514
rect 4874 122918 4926 122970
rect 4938 122918 4990 122970
rect 5002 122918 5054 122970
rect 5066 122918 5118 122970
rect 5130 122918 5182 122970
rect 106658 122918 106710 122970
rect 106722 122918 106774 122970
rect 106786 122918 106838 122970
rect 106850 122918 106902 122970
rect 106914 122918 106966 122970
rect 4214 122374 4266 122426
rect 4278 122374 4330 122426
rect 4342 122374 4394 122426
rect 4406 122374 4458 122426
rect 4470 122374 4522 122426
rect 105922 122374 105974 122426
rect 105986 122374 106038 122426
rect 106050 122374 106102 122426
rect 106114 122374 106166 122426
rect 106178 122374 106230 122426
rect 4874 121830 4926 121882
rect 4938 121830 4990 121882
rect 5002 121830 5054 121882
rect 5066 121830 5118 121882
rect 5130 121830 5182 121882
rect 106658 121830 106710 121882
rect 106722 121830 106774 121882
rect 106786 121830 106838 121882
rect 106850 121830 106902 121882
rect 106914 121830 106966 121882
rect 4214 121286 4266 121338
rect 4278 121286 4330 121338
rect 4342 121286 4394 121338
rect 4406 121286 4458 121338
rect 4470 121286 4522 121338
rect 105922 121286 105974 121338
rect 105986 121286 106038 121338
rect 106050 121286 106102 121338
rect 106114 121286 106166 121338
rect 106178 121286 106230 121338
rect 4874 120742 4926 120794
rect 4938 120742 4990 120794
rect 5002 120742 5054 120794
rect 5066 120742 5118 120794
rect 5130 120742 5182 120794
rect 106658 120742 106710 120794
rect 106722 120742 106774 120794
rect 106786 120742 106838 120794
rect 106850 120742 106902 120794
rect 106914 120742 106966 120794
rect 4214 120198 4266 120250
rect 4278 120198 4330 120250
rect 4342 120198 4394 120250
rect 4406 120198 4458 120250
rect 4470 120198 4522 120250
rect 105922 120198 105974 120250
rect 105986 120198 106038 120250
rect 106050 120198 106102 120250
rect 106114 120198 106166 120250
rect 106178 120198 106230 120250
rect 104348 119935 104400 119944
rect 104348 119901 104357 119935
rect 104357 119901 104391 119935
rect 104391 119901 104400 119935
rect 104348 119892 104400 119901
rect 4874 119654 4926 119706
rect 4938 119654 4990 119706
rect 5002 119654 5054 119706
rect 5066 119654 5118 119706
rect 5130 119654 5182 119706
rect 106658 119654 106710 119706
rect 106722 119654 106774 119706
rect 106786 119654 106838 119706
rect 106850 119654 106902 119706
rect 106914 119654 106966 119706
rect 4214 119110 4266 119162
rect 4278 119110 4330 119162
rect 4342 119110 4394 119162
rect 4406 119110 4458 119162
rect 4470 119110 4522 119162
rect 105922 119110 105974 119162
rect 105986 119110 106038 119162
rect 106050 119110 106102 119162
rect 106114 119110 106166 119162
rect 106178 119110 106230 119162
rect 4874 118566 4926 118618
rect 4938 118566 4990 118618
rect 5002 118566 5054 118618
rect 5066 118566 5118 118618
rect 5130 118566 5182 118618
rect 106658 118566 106710 118618
rect 106722 118566 106774 118618
rect 106786 118566 106838 118618
rect 106850 118566 106902 118618
rect 106914 118566 106966 118618
rect 4214 118022 4266 118074
rect 4278 118022 4330 118074
rect 4342 118022 4394 118074
rect 4406 118022 4458 118074
rect 4470 118022 4522 118074
rect 105922 118022 105974 118074
rect 105986 118022 106038 118074
rect 106050 118022 106102 118074
rect 106114 118022 106166 118074
rect 106178 118022 106230 118074
rect 4874 117478 4926 117530
rect 4938 117478 4990 117530
rect 5002 117478 5054 117530
rect 5066 117478 5118 117530
rect 5130 117478 5182 117530
rect 106658 117478 106710 117530
rect 106722 117478 106774 117530
rect 106786 117478 106838 117530
rect 106850 117478 106902 117530
rect 106914 117478 106966 117530
rect 4214 116934 4266 116986
rect 4278 116934 4330 116986
rect 4342 116934 4394 116986
rect 4406 116934 4458 116986
rect 4470 116934 4522 116986
rect 105922 116934 105974 116986
rect 105986 116934 106038 116986
rect 106050 116934 106102 116986
rect 106114 116934 106166 116986
rect 106178 116934 106230 116986
rect 4874 116390 4926 116442
rect 4938 116390 4990 116442
rect 5002 116390 5054 116442
rect 5066 116390 5118 116442
rect 5130 116390 5182 116442
rect 106658 116390 106710 116442
rect 106722 116390 106774 116442
rect 106786 116390 106838 116442
rect 106850 116390 106902 116442
rect 106914 116390 106966 116442
rect 4214 115846 4266 115898
rect 4278 115846 4330 115898
rect 4342 115846 4394 115898
rect 4406 115846 4458 115898
rect 4470 115846 4522 115898
rect 105922 115846 105974 115898
rect 105986 115846 106038 115898
rect 106050 115846 106102 115898
rect 106114 115846 106166 115898
rect 106178 115846 106230 115898
rect 4874 115302 4926 115354
rect 4938 115302 4990 115354
rect 5002 115302 5054 115354
rect 5066 115302 5118 115354
rect 5130 115302 5182 115354
rect 106658 115302 106710 115354
rect 106722 115302 106774 115354
rect 106786 115302 106838 115354
rect 106850 115302 106902 115354
rect 106914 115302 106966 115354
rect 4214 114758 4266 114810
rect 4278 114758 4330 114810
rect 4342 114758 4394 114810
rect 4406 114758 4458 114810
rect 4470 114758 4522 114810
rect 105922 114758 105974 114810
rect 105986 114758 106038 114810
rect 106050 114758 106102 114810
rect 106114 114758 106166 114810
rect 106178 114758 106230 114810
rect 4874 114214 4926 114266
rect 4938 114214 4990 114266
rect 5002 114214 5054 114266
rect 5066 114214 5118 114266
rect 5130 114214 5182 114266
rect 106658 114214 106710 114266
rect 106722 114214 106774 114266
rect 106786 114214 106838 114266
rect 106850 114214 106902 114266
rect 106914 114214 106966 114266
rect 4214 113670 4266 113722
rect 4278 113670 4330 113722
rect 4342 113670 4394 113722
rect 4406 113670 4458 113722
rect 4470 113670 4522 113722
rect 105922 113670 105974 113722
rect 105986 113670 106038 113722
rect 106050 113670 106102 113722
rect 106114 113670 106166 113722
rect 106178 113670 106230 113722
rect 4874 113126 4926 113178
rect 4938 113126 4990 113178
rect 5002 113126 5054 113178
rect 5066 113126 5118 113178
rect 5130 113126 5182 113178
rect 106658 113126 106710 113178
rect 106722 113126 106774 113178
rect 106786 113126 106838 113178
rect 106850 113126 106902 113178
rect 106914 113126 106966 113178
rect 4214 112582 4266 112634
rect 4278 112582 4330 112634
rect 4342 112582 4394 112634
rect 4406 112582 4458 112634
rect 4470 112582 4522 112634
rect 105922 112582 105974 112634
rect 105986 112582 106038 112634
rect 106050 112582 106102 112634
rect 106114 112582 106166 112634
rect 106178 112582 106230 112634
rect 4874 112038 4926 112090
rect 4938 112038 4990 112090
rect 5002 112038 5054 112090
rect 5066 112038 5118 112090
rect 5130 112038 5182 112090
rect 106658 112038 106710 112090
rect 106722 112038 106774 112090
rect 106786 112038 106838 112090
rect 106850 112038 106902 112090
rect 106914 112038 106966 112090
rect 4214 111494 4266 111546
rect 4278 111494 4330 111546
rect 4342 111494 4394 111546
rect 4406 111494 4458 111546
rect 4470 111494 4522 111546
rect 105922 111494 105974 111546
rect 105986 111494 106038 111546
rect 106050 111494 106102 111546
rect 106114 111494 106166 111546
rect 106178 111494 106230 111546
rect 4874 110950 4926 111002
rect 4938 110950 4990 111002
rect 5002 110950 5054 111002
rect 5066 110950 5118 111002
rect 5130 110950 5182 111002
rect 106658 110950 106710 111002
rect 106722 110950 106774 111002
rect 106786 110950 106838 111002
rect 106850 110950 106902 111002
rect 106914 110950 106966 111002
rect 4214 110406 4266 110458
rect 4278 110406 4330 110458
rect 4342 110406 4394 110458
rect 4406 110406 4458 110458
rect 4470 110406 4522 110458
rect 105922 110406 105974 110458
rect 105986 110406 106038 110458
rect 106050 110406 106102 110458
rect 106114 110406 106166 110458
rect 106178 110406 106230 110458
rect 4874 109862 4926 109914
rect 4938 109862 4990 109914
rect 5002 109862 5054 109914
rect 5066 109862 5118 109914
rect 5130 109862 5182 109914
rect 106658 109862 106710 109914
rect 106722 109862 106774 109914
rect 106786 109862 106838 109914
rect 106850 109862 106902 109914
rect 106914 109862 106966 109914
rect 4214 109318 4266 109370
rect 4278 109318 4330 109370
rect 4342 109318 4394 109370
rect 4406 109318 4458 109370
rect 4470 109318 4522 109370
rect 105922 109318 105974 109370
rect 105986 109318 106038 109370
rect 106050 109318 106102 109370
rect 106114 109318 106166 109370
rect 106178 109318 106230 109370
rect 4874 108774 4926 108826
rect 4938 108774 4990 108826
rect 5002 108774 5054 108826
rect 5066 108774 5118 108826
rect 5130 108774 5182 108826
rect 106658 108774 106710 108826
rect 106722 108774 106774 108826
rect 106786 108774 106838 108826
rect 106850 108774 106902 108826
rect 106914 108774 106966 108826
rect 4214 108230 4266 108282
rect 4278 108230 4330 108282
rect 4342 108230 4394 108282
rect 4406 108230 4458 108282
rect 4470 108230 4522 108282
rect 105922 108230 105974 108282
rect 105986 108230 106038 108282
rect 106050 108230 106102 108282
rect 106114 108230 106166 108282
rect 106178 108230 106230 108282
rect 4874 107686 4926 107738
rect 4938 107686 4990 107738
rect 5002 107686 5054 107738
rect 5066 107686 5118 107738
rect 5130 107686 5182 107738
rect 106658 107686 106710 107738
rect 106722 107686 106774 107738
rect 106786 107686 106838 107738
rect 106850 107686 106902 107738
rect 106914 107686 106966 107738
rect 4214 107142 4266 107194
rect 4278 107142 4330 107194
rect 4342 107142 4394 107194
rect 4406 107142 4458 107194
rect 4470 107142 4522 107194
rect 105922 107142 105974 107194
rect 105986 107142 106038 107194
rect 106050 107142 106102 107194
rect 106114 107142 106166 107194
rect 106178 107142 106230 107194
rect 4874 106598 4926 106650
rect 4938 106598 4990 106650
rect 5002 106598 5054 106650
rect 5066 106598 5118 106650
rect 5130 106598 5182 106650
rect 106658 106598 106710 106650
rect 106722 106598 106774 106650
rect 106786 106598 106838 106650
rect 106850 106598 106902 106650
rect 106914 106598 106966 106650
rect 4214 106054 4266 106106
rect 4278 106054 4330 106106
rect 4342 106054 4394 106106
rect 4406 106054 4458 106106
rect 4470 106054 4522 106106
rect 105922 106054 105974 106106
rect 105986 106054 106038 106106
rect 106050 106054 106102 106106
rect 106114 106054 106166 106106
rect 106178 106054 106230 106106
rect 4874 105510 4926 105562
rect 4938 105510 4990 105562
rect 5002 105510 5054 105562
rect 5066 105510 5118 105562
rect 5130 105510 5182 105562
rect 106658 105510 106710 105562
rect 106722 105510 106774 105562
rect 106786 105510 106838 105562
rect 106850 105510 106902 105562
rect 106914 105510 106966 105562
rect 4214 104966 4266 105018
rect 4278 104966 4330 105018
rect 4342 104966 4394 105018
rect 4406 104966 4458 105018
rect 4470 104966 4522 105018
rect 105922 104966 105974 105018
rect 105986 104966 106038 105018
rect 106050 104966 106102 105018
rect 106114 104966 106166 105018
rect 106178 104966 106230 105018
rect 4874 104422 4926 104474
rect 4938 104422 4990 104474
rect 5002 104422 5054 104474
rect 5066 104422 5118 104474
rect 5130 104422 5182 104474
rect 106658 104422 106710 104474
rect 106722 104422 106774 104474
rect 106786 104422 106838 104474
rect 106850 104422 106902 104474
rect 106914 104422 106966 104474
rect 4214 103878 4266 103930
rect 4278 103878 4330 103930
rect 4342 103878 4394 103930
rect 4406 103878 4458 103930
rect 4470 103878 4522 103930
rect 105922 103878 105974 103930
rect 105986 103878 106038 103930
rect 106050 103878 106102 103930
rect 106114 103878 106166 103930
rect 106178 103878 106230 103930
rect 4874 103334 4926 103386
rect 4938 103334 4990 103386
rect 5002 103334 5054 103386
rect 5066 103334 5118 103386
rect 5130 103334 5182 103386
rect 106658 103334 106710 103386
rect 106722 103334 106774 103386
rect 106786 103334 106838 103386
rect 106850 103334 106902 103386
rect 106914 103334 106966 103386
rect 4214 102790 4266 102842
rect 4278 102790 4330 102842
rect 4342 102790 4394 102842
rect 4406 102790 4458 102842
rect 4470 102790 4522 102842
rect 105922 102790 105974 102842
rect 105986 102790 106038 102842
rect 106050 102790 106102 102842
rect 106114 102790 106166 102842
rect 106178 102790 106230 102842
rect 4874 102246 4926 102298
rect 4938 102246 4990 102298
rect 5002 102246 5054 102298
rect 5066 102246 5118 102298
rect 5130 102246 5182 102298
rect 106658 102246 106710 102298
rect 106722 102246 106774 102298
rect 106786 102246 106838 102298
rect 106850 102246 106902 102298
rect 106914 102246 106966 102298
rect 4214 101702 4266 101754
rect 4278 101702 4330 101754
rect 4342 101702 4394 101754
rect 4406 101702 4458 101754
rect 4470 101702 4522 101754
rect 105922 101702 105974 101754
rect 105986 101702 106038 101754
rect 106050 101702 106102 101754
rect 106114 101702 106166 101754
rect 106178 101702 106230 101754
rect 8392 101532 8444 101584
rect 1216 101396 1268 101448
rect 4874 101158 4926 101210
rect 4938 101158 4990 101210
rect 5002 101158 5054 101210
rect 5066 101158 5118 101210
rect 5130 101158 5182 101210
rect 106658 101158 106710 101210
rect 106722 101158 106774 101210
rect 106786 101158 106838 101210
rect 106850 101158 106902 101210
rect 106914 101158 106966 101210
rect 4214 100614 4266 100666
rect 4278 100614 4330 100666
rect 4342 100614 4394 100666
rect 4406 100614 4458 100666
rect 4470 100614 4522 100666
rect 105922 100614 105974 100666
rect 105986 100614 106038 100666
rect 106050 100614 106102 100666
rect 106114 100614 106166 100666
rect 106178 100614 106230 100666
rect 4874 100070 4926 100122
rect 4938 100070 4990 100122
rect 5002 100070 5054 100122
rect 5066 100070 5118 100122
rect 5130 100070 5182 100122
rect 106658 100070 106710 100122
rect 106722 100070 106774 100122
rect 106786 100070 106838 100122
rect 106850 100070 106902 100122
rect 106914 100070 106966 100122
rect 1400 99875 1452 99884
rect 1400 99841 1409 99875
rect 1409 99841 1443 99875
rect 1443 99841 1452 99875
rect 1400 99832 1452 99841
rect 8392 99696 8444 99748
rect 4214 99526 4266 99578
rect 4278 99526 4330 99578
rect 4342 99526 4394 99578
rect 4406 99526 4458 99578
rect 4470 99526 4522 99578
rect 105922 99526 105974 99578
rect 105986 99526 106038 99578
rect 106050 99526 106102 99578
rect 106114 99526 106166 99578
rect 106178 99526 106230 99578
rect 4874 98982 4926 99034
rect 4938 98982 4990 99034
rect 5002 98982 5054 99034
rect 5066 98982 5118 99034
rect 5130 98982 5182 99034
rect 106658 98982 106710 99034
rect 106722 98982 106774 99034
rect 106786 98982 106838 99034
rect 106850 98982 106902 99034
rect 106914 98982 106966 99034
rect 1308 98744 1360 98796
rect 8392 98608 8444 98660
rect 4214 98438 4266 98490
rect 4278 98438 4330 98490
rect 4342 98438 4394 98490
rect 4406 98438 4458 98490
rect 4470 98438 4522 98490
rect 105922 98438 105974 98490
rect 105986 98438 106038 98490
rect 106050 98438 106102 98490
rect 106114 98438 106166 98490
rect 106178 98438 106230 98490
rect 4874 97894 4926 97946
rect 4938 97894 4990 97946
rect 5002 97894 5054 97946
rect 5066 97894 5118 97946
rect 5130 97894 5182 97946
rect 106658 97894 106710 97946
rect 106722 97894 106774 97946
rect 106786 97894 106838 97946
rect 106850 97894 106902 97946
rect 106914 97894 106966 97946
rect 4214 97350 4266 97402
rect 4278 97350 4330 97402
rect 4342 97350 4394 97402
rect 4406 97350 4458 97402
rect 4470 97350 4522 97402
rect 105922 97350 105974 97402
rect 105986 97350 106038 97402
rect 106050 97350 106102 97402
rect 106114 97350 106166 97402
rect 106178 97350 106230 97402
rect 8392 97180 8444 97232
rect 1308 97044 1360 97096
rect 4874 96806 4926 96858
rect 4938 96806 4990 96858
rect 5002 96806 5054 96858
rect 5066 96806 5118 96858
rect 5130 96806 5182 96858
rect 106658 96806 106710 96858
rect 106722 96806 106774 96858
rect 106786 96806 106838 96858
rect 106850 96806 106902 96858
rect 106914 96806 106966 96858
rect 4214 96262 4266 96314
rect 4278 96262 4330 96314
rect 4342 96262 4394 96314
rect 4406 96262 4458 96314
rect 4470 96262 4522 96314
rect 105922 96262 105974 96314
rect 105986 96262 106038 96314
rect 106050 96262 106102 96314
rect 106114 96262 106166 96314
rect 106178 96262 106230 96314
rect 8392 96092 8444 96144
rect 1216 95956 1268 96008
rect 4874 95718 4926 95770
rect 4938 95718 4990 95770
rect 5002 95718 5054 95770
rect 5066 95718 5118 95770
rect 5130 95718 5182 95770
rect 106658 95718 106710 95770
rect 106722 95718 106774 95770
rect 106786 95718 106838 95770
rect 106850 95718 106902 95770
rect 106914 95718 106966 95770
rect 4214 95174 4266 95226
rect 4278 95174 4330 95226
rect 4342 95174 4394 95226
rect 4406 95174 4458 95226
rect 4470 95174 4522 95226
rect 105922 95174 105974 95226
rect 105986 95174 106038 95226
rect 106050 95174 106102 95226
rect 106114 95174 106166 95226
rect 106178 95174 106230 95226
rect 4874 94630 4926 94682
rect 4938 94630 4990 94682
rect 5002 94630 5054 94682
rect 5066 94630 5118 94682
rect 5130 94630 5182 94682
rect 106658 94630 106710 94682
rect 106722 94630 106774 94682
rect 106786 94630 106838 94682
rect 106850 94630 106902 94682
rect 106914 94630 106966 94682
rect 1308 94392 1360 94444
rect 8392 94256 8444 94308
rect 4214 94086 4266 94138
rect 4278 94086 4330 94138
rect 4342 94086 4394 94138
rect 4406 94086 4458 94138
rect 4470 94086 4522 94138
rect 105922 94086 105974 94138
rect 105986 94086 106038 94138
rect 106050 94086 106102 94138
rect 106114 94086 106166 94138
rect 106178 94086 106230 94138
rect 4874 93542 4926 93594
rect 4938 93542 4990 93594
rect 5002 93542 5054 93594
rect 5066 93542 5118 93594
rect 5130 93542 5182 93594
rect 106658 93542 106710 93594
rect 106722 93542 106774 93594
rect 106786 93542 106838 93594
rect 106850 93542 106902 93594
rect 106914 93542 106966 93594
rect 4214 92998 4266 93050
rect 4278 92998 4330 93050
rect 4342 92998 4394 93050
rect 4406 92998 4458 93050
rect 4470 92998 4522 93050
rect 105922 92998 105974 93050
rect 105986 92998 106038 93050
rect 106050 92998 106102 93050
rect 106114 92998 106166 93050
rect 106178 92998 106230 93050
rect 4874 92454 4926 92506
rect 4938 92454 4990 92506
rect 5002 92454 5054 92506
rect 5066 92454 5118 92506
rect 5130 92454 5182 92506
rect 106658 92454 106710 92506
rect 106722 92454 106774 92506
rect 106786 92454 106838 92506
rect 106850 92454 106902 92506
rect 106914 92454 106966 92506
rect 4214 91910 4266 91962
rect 4278 91910 4330 91962
rect 4342 91910 4394 91962
rect 4406 91910 4458 91962
rect 4470 91910 4522 91962
rect 105922 91910 105974 91962
rect 105986 91910 106038 91962
rect 106050 91910 106102 91962
rect 106114 91910 106166 91962
rect 106178 91910 106230 91962
rect 4874 91366 4926 91418
rect 4938 91366 4990 91418
rect 5002 91366 5054 91418
rect 5066 91366 5118 91418
rect 5130 91366 5182 91418
rect 106658 91366 106710 91418
rect 106722 91366 106774 91418
rect 106786 91366 106838 91418
rect 106850 91366 106902 91418
rect 106914 91366 106966 91418
rect 4214 90822 4266 90874
rect 4278 90822 4330 90874
rect 4342 90822 4394 90874
rect 4406 90822 4458 90874
rect 4470 90822 4522 90874
rect 105922 90822 105974 90874
rect 105986 90822 106038 90874
rect 106050 90822 106102 90874
rect 106114 90822 106166 90874
rect 106178 90822 106230 90874
rect 4874 90278 4926 90330
rect 4938 90278 4990 90330
rect 5002 90278 5054 90330
rect 5066 90278 5118 90330
rect 5130 90278 5182 90330
rect 106658 90278 106710 90330
rect 106722 90278 106774 90330
rect 106786 90278 106838 90330
rect 106850 90278 106902 90330
rect 106914 90278 106966 90330
rect 4214 89734 4266 89786
rect 4278 89734 4330 89786
rect 4342 89734 4394 89786
rect 4406 89734 4458 89786
rect 4470 89734 4522 89786
rect 105922 89734 105974 89786
rect 105986 89734 106038 89786
rect 106050 89734 106102 89786
rect 106114 89734 106166 89786
rect 106178 89734 106230 89786
rect 4874 89190 4926 89242
rect 4938 89190 4990 89242
rect 5002 89190 5054 89242
rect 5066 89190 5118 89242
rect 5130 89190 5182 89242
rect 106658 89190 106710 89242
rect 106722 89190 106774 89242
rect 106786 89190 106838 89242
rect 106850 89190 106902 89242
rect 106914 89190 106966 89242
rect 4214 88646 4266 88698
rect 4278 88646 4330 88698
rect 4342 88646 4394 88698
rect 4406 88646 4458 88698
rect 4470 88646 4522 88698
rect 105922 88646 105974 88698
rect 105986 88646 106038 88698
rect 106050 88646 106102 88698
rect 106114 88646 106166 88698
rect 106178 88646 106230 88698
rect 4874 88102 4926 88154
rect 4938 88102 4990 88154
rect 5002 88102 5054 88154
rect 5066 88102 5118 88154
rect 5130 88102 5182 88154
rect 106658 88102 106710 88154
rect 106722 88102 106774 88154
rect 106786 88102 106838 88154
rect 106850 88102 106902 88154
rect 106914 88102 106966 88154
rect 4214 87558 4266 87610
rect 4278 87558 4330 87610
rect 4342 87558 4394 87610
rect 4406 87558 4458 87610
rect 4470 87558 4522 87610
rect 105922 87558 105974 87610
rect 105986 87558 106038 87610
rect 106050 87558 106102 87610
rect 106114 87558 106166 87610
rect 106178 87558 106230 87610
rect 4874 87014 4926 87066
rect 4938 87014 4990 87066
rect 5002 87014 5054 87066
rect 5066 87014 5118 87066
rect 5130 87014 5182 87066
rect 106658 87014 106710 87066
rect 106722 87014 106774 87066
rect 106786 87014 106838 87066
rect 106850 87014 106902 87066
rect 106914 87014 106966 87066
rect 4214 86470 4266 86522
rect 4278 86470 4330 86522
rect 4342 86470 4394 86522
rect 4406 86470 4458 86522
rect 4470 86470 4522 86522
rect 105922 86470 105974 86522
rect 105986 86470 106038 86522
rect 106050 86470 106102 86522
rect 106114 86470 106166 86522
rect 106178 86470 106230 86522
rect 104716 86411 104768 86420
rect 104716 86377 104725 86411
rect 104725 86377 104759 86411
rect 104759 86377 104768 86411
rect 104716 86368 104768 86377
rect 104808 86096 104860 86148
rect 4874 85926 4926 85978
rect 4938 85926 4990 85978
rect 5002 85926 5054 85978
rect 5066 85926 5118 85978
rect 5130 85926 5182 85978
rect 106658 85926 106710 85978
rect 106722 85926 106774 85978
rect 106786 85926 106838 85978
rect 106850 85926 106902 85978
rect 106914 85926 106966 85978
rect 104716 85688 104768 85740
rect 104808 85620 104860 85672
rect 105820 85552 105872 85604
rect 4214 85382 4266 85434
rect 4278 85382 4330 85434
rect 4342 85382 4394 85434
rect 4406 85382 4458 85434
rect 4470 85382 4522 85434
rect 105922 85382 105974 85434
rect 105986 85382 106038 85434
rect 106050 85382 106102 85434
rect 106114 85382 106166 85434
rect 106178 85382 106230 85434
rect 104440 85323 104492 85332
rect 104440 85289 104449 85323
rect 104449 85289 104483 85323
rect 104483 85289 104492 85323
rect 104440 85280 104492 85289
rect 104716 85076 104768 85128
rect 4874 84838 4926 84890
rect 4938 84838 4990 84890
rect 5002 84838 5054 84890
rect 5066 84838 5118 84890
rect 5130 84838 5182 84890
rect 106658 84838 106710 84890
rect 106722 84838 106774 84890
rect 106786 84838 106838 84890
rect 106850 84838 106902 84890
rect 106914 84838 106966 84890
rect 4214 84294 4266 84346
rect 4278 84294 4330 84346
rect 4342 84294 4394 84346
rect 4406 84294 4458 84346
rect 4470 84294 4522 84346
rect 105922 84294 105974 84346
rect 105986 84294 106038 84346
rect 106050 84294 106102 84346
rect 106114 84294 106166 84346
rect 106178 84294 106230 84346
rect 4874 83750 4926 83802
rect 4938 83750 4990 83802
rect 5002 83750 5054 83802
rect 5066 83750 5118 83802
rect 5130 83750 5182 83802
rect 106658 83750 106710 83802
rect 106722 83750 106774 83802
rect 106786 83750 106838 83802
rect 106850 83750 106902 83802
rect 106914 83750 106966 83802
rect 4214 83206 4266 83258
rect 4278 83206 4330 83258
rect 4342 83206 4394 83258
rect 4406 83206 4458 83258
rect 4470 83206 4522 83258
rect 105922 83206 105974 83258
rect 105986 83206 106038 83258
rect 106050 83206 106102 83258
rect 106114 83206 106166 83258
rect 106178 83206 106230 83258
rect 4874 82662 4926 82714
rect 4938 82662 4990 82714
rect 5002 82662 5054 82714
rect 5066 82662 5118 82714
rect 5130 82662 5182 82714
rect 106658 82662 106710 82714
rect 106722 82662 106774 82714
rect 106786 82662 106838 82714
rect 106850 82662 106902 82714
rect 106914 82662 106966 82714
rect 4214 82118 4266 82170
rect 4278 82118 4330 82170
rect 4342 82118 4394 82170
rect 4406 82118 4458 82170
rect 4470 82118 4522 82170
rect 105922 82118 105974 82170
rect 105986 82118 106038 82170
rect 106050 82118 106102 82170
rect 106114 82118 106166 82170
rect 106178 82118 106230 82170
rect 4874 81574 4926 81626
rect 4938 81574 4990 81626
rect 5002 81574 5054 81626
rect 5066 81574 5118 81626
rect 5130 81574 5182 81626
rect 106658 81574 106710 81626
rect 106722 81574 106774 81626
rect 106786 81574 106838 81626
rect 106850 81574 106902 81626
rect 106914 81574 106966 81626
rect 4214 81030 4266 81082
rect 4278 81030 4330 81082
rect 4342 81030 4394 81082
rect 4406 81030 4458 81082
rect 4470 81030 4522 81082
rect 105922 81030 105974 81082
rect 105986 81030 106038 81082
rect 106050 81030 106102 81082
rect 106114 81030 106166 81082
rect 106178 81030 106230 81082
rect 4874 80486 4926 80538
rect 4938 80486 4990 80538
rect 5002 80486 5054 80538
rect 5066 80486 5118 80538
rect 5130 80486 5182 80538
rect 106658 80486 106710 80538
rect 106722 80486 106774 80538
rect 106786 80486 106838 80538
rect 106850 80486 106902 80538
rect 106914 80486 106966 80538
rect 104164 80248 104216 80300
rect 104532 80044 104584 80096
rect 4214 79942 4266 79994
rect 4278 79942 4330 79994
rect 4342 79942 4394 79994
rect 4406 79942 4458 79994
rect 4470 79942 4522 79994
rect 105922 79942 105974 79994
rect 105986 79942 106038 79994
rect 106050 79942 106102 79994
rect 106114 79942 106166 79994
rect 106178 79942 106230 79994
rect 4874 79398 4926 79450
rect 4938 79398 4990 79450
rect 5002 79398 5054 79450
rect 5066 79398 5118 79450
rect 5130 79398 5182 79450
rect 106658 79398 106710 79450
rect 106722 79398 106774 79450
rect 106786 79398 106838 79450
rect 106850 79398 106902 79450
rect 106914 79398 106966 79450
rect 104072 79092 104124 79144
rect 105176 79092 105228 79144
rect 103888 78956 103940 79008
rect 4214 78854 4266 78906
rect 4278 78854 4330 78906
rect 4342 78854 4394 78906
rect 4406 78854 4458 78906
rect 4470 78854 4522 78906
rect 105922 78854 105974 78906
rect 105986 78854 106038 78906
rect 106050 78854 106102 78906
rect 106114 78854 106166 78906
rect 106178 78854 106230 78906
rect 104624 78752 104676 78804
rect 104440 78659 104492 78668
rect 104440 78625 104463 78659
rect 104463 78625 104492 78659
rect 104440 78616 104492 78625
rect 104256 78548 104308 78600
rect 1308 78480 1360 78532
rect 7564 78480 7616 78532
rect 104072 78480 104124 78532
rect 105176 78591 105228 78600
rect 105176 78557 105185 78591
rect 105185 78557 105219 78591
rect 105219 78557 105228 78591
rect 105176 78548 105228 78557
rect 103888 78412 103940 78464
rect 104808 78480 104860 78532
rect 104716 78455 104768 78464
rect 104716 78421 104725 78455
rect 104725 78421 104759 78455
rect 104759 78421 104768 78455
rect 104716 78412 104768 78421
rect 105544 78455 105596 78464
rect 105544 78421 105553 78455
rect 105553 78421 105587 78455
rect 105587 78421 105596 78455
rect 105544 78412 105596 78421
rect 4874 78310 4926 78362
rect 4938 78310 4990 78362
rect 5002 78310 5054 78362
rect 5066 78310 5118 78362
rect 5130 78310 5182 78362
rect 106658 78310 106710 78362
rect 106722 78310 106774 78362
rect 106786 78310 106838 78362
rect 106850 78310 106902 78362
rect 106914 78310 106966 78362
rect 104440 78208 104492 78260
rect 104624 78208 104676 78260
rect 105544 78208 105596 78260
rect 1308 78072 1360 78124
rect 104440 78072 104492 78124
rect 7656 77936 7708 77988
rect 105636 77911 105688 77920
rect 105636 77877 105645 77911
rect 105645 77877 105679 77911
rect 105679 77877 105688 77911
rect 105636 77868 105688 77877
rect 106280 77868 106332 77920
rect 4214 77766 4266 77818
rect 4278 77766 4330 77818
rect 4342 77766 4394 77818
rect 4406 77766 4458 77818
rect 4470 77766 4522 77818
rect 105922 77766 105974 77818
rect 105986 77766 106038 77818
rect 106050 77766 106102 77818
rect 106114 77766 106166 77818
rect 106178 77766 106230 77818
rect 102784 77460 102836 77512
rect 105636 77460 105688 77512
rect 104440 77324 104492 77376
rect 4874 77222 4926 77274
rect 4938 77222 4990 77274
rect 5002 77222 5054 77274
rect 5066 77222 5118 77274
rect 5130 77222 5182 77274
rect 106658 77222 106710 77274
rect 106722 77222 106774 77274
rect 106786 77222 106838 77274
rect 106850 77222 106902 77274
rect 106914 77222 106966 77274
rect 1216 76984 1268 77036
rect 8944 76848 8996 76900
rect 4214 76678 4266 76730
rect 4278 76678 4330 76730
rect 4342 76678 4394 76730
rect 4406 76678 4458 76730
rect 4470 76678 4522 76730
rect 105922 76678 105974 76730
rect 105986 76678 106038 76730
rect 106050 76678 106102 76730
rect 106114 76678 106166 76730
rect 106178 76678 106230 76730
rect 1216 76304 1268 76356
rect 8852 76304 8904 76356
rect 4874 76134 4926 76186
rect 4938 76134 4990 76186
rect 5002 76134 5054 76186
rect 5066 76134 5118 76186
rect 5130 76134 5182 76186
rect 106658 76134 106710 76186
rect 106722 76134 106774 76186
rect 106786 76134 106838 76186
rect 106850 76134 106902 76186
rect 106914 76134 106966 76186
rect 5540 76032 5592 76084
rect 104256 76032 104308 76084
rect 104532 75964 104584 76016
rect 1400 75939 1452 75948
rect 1400 75905 1409 75939
rect 1409 75905 1443 75939
rect 1443 75905 1452 75939
rect 1400 75896 1452 75905
rect 106280 76032 106332 76084
rect 105820 75871 105872 75880
rect 105820 75837 105829 75871
rect 105829 75837 105863 75871
rect 105863 75837 105872 75871
rect 105820 75828 105872 75837
rect 4214 75590 4266 75642
rect 4278 75590 4330 75642
rect 4342 75590 4394 75642
rect 4406 75590 4458 75642
rect 4470 75590 4522 75642
rect 105922 75590 105974 75642
rect 105986 75590 106038 75642
rect 106050 75590 106102 75642
rect 106114 75590 106166 75642
rect 106178 75590 106230 75642
rect 104256 75284 104308 75336
rect 1308 75216 1360 75268
rect 6920 75216 6972 75268
rect 102048 75148 102100 75200
rect 4874 75046 4926 75098
rect 4938 75046 4990 75098
rect 5002 75046 5054 75098
rect 5066 75046 5118 75098
rect 5130 75046 5182 75098
rect 106658 75046 106710 75098
rect 106722 75046 106774 75098
rect 106786 75046 106838 75098
rect 106850 75046 106902 75098
rect 106914 75046 106966 75098
rect 4214 74502 4266 74554
rect 4278 74502 4330 74554
rect 4342 74502 4394 74554
rect 4406 74502 4458 74554
rect 4470 74502 4522 74554
rect 105922 74502 105974 74554
rect 105986 74502 106038 74554
rect 106050 74502 106102 74554
rect 106114 74502 106166 74554
rect 106178 74502 106230 74554
rect 1216 74128 1268 74180
rect 1860 74103 1912 74112
rect 1860 74069 1869 74103
rect 1869 74069 1903 74103
rect 1903 74069 1912 74103
rect 1860 74060 1912 74069
rect 4874 73958 4926 74010
rect 4938 73958 4990 74010
rect 5002 73958 5054 74010
rect 5066 73958 5118 74010
rect 5130 73958 5182 74010
rect 106658 73958 106710 74010
rect 106722 73958 106774 74010
rect 106786 73958 106838 74010
rect 106850 73958 106902 74010
rect 106914 73958 106966 74010
rect 1308 73720 1360 73772
rect 9128 73720 9180 73772
rect 9588 73720 9640 73772
rect 9588 73584 9640 73636
rect 4214 73414 4266 73466
rect 4278 73414 4330 73466
rect 4342 73414 4394 73466
rect 4406 73414 4458 73466
rect 4470 73414 4522 73466
rect 105922 73414 105974 73466
rect 105986 73414 106038 73466
rect 106050 73414 106102 73466
rect 106114 73414 106166 73466
rect 106178 73414 106230 73466
rect 9036 73176 9088 73228
rect 1492 73083 1544 73092
rect 1492 73049 1501 73083
rect 1501 73049 1535 73083
rect 1535 73049 1544 73083
rect 1492 73040 1544 73049
rect 4874 72870 4926 72922
rect 4938 72870 4990 72922
rect 5002 72870 5054 72922
rect 5066 72870 5118 72922
rect 5130 72870 5182 72922
rect 106658 72870 106710 72922
rect 106722 72870 106774 72922
rect 106786 72870 106838 72922
rect 106850 72870 106902 72922
rect 106914 72870 106966 72922
rect 1308 72632 1360 72684
rect 9496 72496 9548 72548
rect 4214 72326 4266 72378
rect 4278 72326 4330 72378
rect 4342 72326 4394 72378
rect 4406 72326 4458 72378
rect 4470 72326 4522 72378
rect 105922 72326 105974 72378
rect 105986 72326 106038 72378
rect 106050 72326 106102 72378
rect 106114 72326 106166 72378
rect 106178 72326 106230 72378
rect 4874 71782 4926 71834
rect 4938 71782 4990 71834
rect 5002 71782 5054 71834
rect 5066 71782 5118 71834
rect 5130 71782 5182 71834
rect 106658 71782 106710 71834
rect 106722 71782 106774 71834
rect 106786 71782 106838 71834
rect 106850 71782 106902 71834
rect 106914 71782 106966 71834
rect 1860 71680 1912 71732
rect 9404 71680 9456 71732
rect 1216 71544 1268 71596
rect 1860 71383 1912 71392
rect 1860 71349 1869 71383
rect 1869 71349 1903 71383
rect 1903 71349 1912 71383
rect 1860 71340 1912 71349
rect 4214 71238 4266 71290
rect 4278 71238 4330 71290
rect 4342 71238 4394 71290
rect 4406 71238 4458 71290
rect 4470 71238 4522 71290
rect 105922 71238 105974 71290
rect 105986 71238 106038 71290
rect 106050 71238 106102 71290
rect 106114 71238 106166 71290
rect 106178 71238 106230 71290
rect 9220 70932 9272 70984
rect 1308 70864 1360 70916
rect 2228 70796 2280 70848
rect 4874 70694 4926 70746
rect 4938 70694 4990 70746
rect 5002 70694 5054 70746
rect 5066 70694 5118 70746
rect 5130 70694 5182 70746
rect 106658 70694 106710 70746
rect 106722 70694 106774 70746
rect 106786 70694 106838 70746
rect 106850 70694 106902 70746
rect 106914 70694 106966 70746
rect 2228 70431 2280 70440
rect 2228 70397 2237 70431
rect 2237 70397 2271 70431
rect 2271 70397 2280 70431
rect 2228 70388 2280 70397
rect 8392 70388 8444 70440
rect 4214 70150 4266 70202
rect 4278 70150 4330 70202
rect 4342 70150 4394 70202
rect 4406 70150 4458 70202
rect 4470 70150 4522 70202
rect 105922 70150 105974 70202
rect 105986 70150 106038 70202
rect 106050 70150 106102 70202
rect 106114 70150 106166 70202
rect 106178 70150 106230 70202
rect 1860 69980 1912 70032
rect 38660 69980 38712 70032
rect 73620 69980 73672 70032
rect 103704 69980 103756 70032
rect 9588 69912 9640 69964
rect 43260 69912 43312 69964
rect 71780 69912 71832 69964
rect 102692 69912 102744 69964
rect 9036 69844 9088 69896
rect 40960 69844 41012 69896
rect 70952 69844 71004 69896
rect 103612 69844 103664 69896
rect 1308 69776 1360 69828
rect 9496 69776 9548 69828
rect 39764 69776 39816 69828
rect 69296 69776 69348 69828
rect 102508 69776 102560 69828
rect 37464 69708 37516 69760
rect 68468 69708 68520 69760
rect 102600 69708 102652 69760
rect 107568 69708 107620 69760
rect 108488 69751 108540 69760
rect 108488 69717 108497 69751
rect 108497 69717 108531 69751
rect 108531 69717 108540 69751
rect 108488 69708 108540 69717
rect 4874 69606 4926 69658
rect 4938 69606 4990 69658
rect 5002 69606 5054 69658
rect 5066 69606 5118 69658
rect 5130 69606 5182 69658
rect 66996 69640 67048 69692
rect 103520 69640 103572 69692
rect 106658 69606 106710 69658
rect 106722 69606 106774 69658
rect 106786 69606 106838 69658
rect 106850 69606 106902 69658
rect 106914 69606 106966 69658
rect 7656 69504 7708 69556
rect 32864 69504 32916 69556
rect 7564 69436 7616 69488
rect 36360 69436 36412 69488
rect 6920 69368 6972 69420
rect 35164 69368 35216 69420
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 105922 69062 105974 69114
rect 105986 69062 106038 69114
rect 106050 69062 106102 69114
rect 106114 69062 106166 69114
rect 106178 69062 106230 69114
rect 88616 68756 88668 68808
rect 1216 68688 1268 68740
rect 95884 68688 95936 68740
rect 42156 68620 42208 68672
rect 97172 68620 97224 68672
rect 103704 68620 103756 68672
rect 4874 68518 4926 68570
rect 4938 68518 4990 68570
rect 5002 68518 5054 68570
rect 5066 68518 5118 68570
rect 5130 68518 5182 68570
rect 7840 68416 7892 68468
rect 33600 68416 33652 68468
rect 108488 68663 108540 68672
rect 108488 68629 108497 68663
rect 108497 68629 108531 68663
rect 108531 68629 108540 68663
rect 108488 68620 108540 68629
rect 106658 68518 106710 68570
rect 106722 68518 106774 68570
rect 106786 68518 106838 68570
rect 106850 68518 106902 68570
rect 106914 68518 106966 68570
rect 7932 68348 7984 68400
rect 33692 68348 33744 68400
rect 88340 68348 88392 68400
rect 93584 68348 93636 68400
rect 1308 68280 1360 68332
rect 9312 68280 9364 68332
rect 35992 68280 36044 68332
rect 90640 68280 90692 68332
rect 95700 68280 95752 68332
rect 2044 68212 2096 68264
rect 89168 68212 89220 68264
rect 30472 68144 30524 68196
rect 90732 68144 90784 68196
rect 91560 68144 91612 68196
rect 94044 68212 94096 68264
rect 103796 68212 103848 68264
rect 25780 68076 25832 68128
rect 88892 68076 88944 68128
rect 93492 68076 93544 68128
rect 96068 68144 96120 68196
rect 102600 68144 102652 68196
rect 95608 68076 95660 68128
rect 96160 68076 96212 68128
rect 103704 68076 103756 68128
rect 104164 68076 104216 68128
rect 108488 68119 108540 68128
rect 108488 68085 108497 68119
rect 108497 68085 108531 68119
rect 108531 68085 108540 68119
rect 108488 68076 108540 68085
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 65654 67974 65706 68026
rect 65718 67974 65770 68026
rect 65782 67974 65834 68026
rect 65846 67974 65898 68026
rect 65910 67974 65962 68026
rect 96374 67974 96426 68026
rect 96438 67974 96490 68026
rect 96502 67974 96554 68026
rect 96566 67974 96618 68026
rect 96630 67974 96682 68026
rect 105922 67974 105974 68026
rect 105986 67974 106038 68026
rect 106050 67974 106102 68026
rect 106114 67974 106166 68026
rect 106178 67974 106230 68026
rect 2044 67872 2096 67924
rect 23480 67915 23532 67924
rect 1676 67804 1728 67856
rect 23480 67881 23489 67915
rect 23489 67881 23523 67915
rect 23523 67881 23532 67915
rect 23480 67872 23532 67881
rect 24676 67915 24728 67924
rect 24676 67881 24685 67915
rect 24685 67881 24719 67915
rect 24719 67881 24728 67915
rect 24676 67872 24728 67881
rect 25780 67872 25832 67924
rect 26976 67915 27028 67924
rect 26976 67881 26985 67915
rect 26985 67881 27019 67915
rect 27019 67881 27028 67915
rect 26976 67872 27028 67881
rect 29552 67915 29604 67924
rect 29552 67881 29561 67915
rect 29561 67881 29595 67915
rect 29595 67881 29604 67915
rect 29552 67872 29604 67881
rect 30472 67915 30524 67924
rect 30472 67881 30481 67915
rect 30481 67881 30515 67915
rect 30515 67881 30524 67915
rect 30472 67872 30524 67881
rect 31760 67915 31812 67924
rect 31760 67881 31769 67915
rect 31769 67881 31803 67915
rect 31803 67881 31812 67915
rect 31760 67872 31812 67881
rect 32864 67915 32916 67924
rect 32864 67881 32873 67915
rect 32873 67881 32907 67915
rect 32907 67881 32916 67915
rect 32864 67872 32916 67881
rect 33968 67915 34020 67924
rect 33968 67881 33977 67915
rect 33977 67881 34011 67915
rect 34011 67881 34020 67915
rect 33968 67872 34020 67881
rect 35164 67915 35216 67924
rect 35164 67881 35173 67915
rect 35173 67881 35207 67915
rect 35207 67881 35216 67915
rect 35164 67872 35216 67881
rect 36360 67915 36412 67924
rect 36360 67881 36369 67915
rect 36369 67881 36403 67915
rect 36403 67881 36412 67915
rect 36360 67872 36412 67881
rect 37464 67915 37516 67924
rect 37464 67881 37473 67915
rect 37473 67881 37507 67915
rect 37507 67881 37516 67915
rect 37464 67872 37516 67881
rect 38660 67915 38712 67924
rect 38660 67881 38669 67915
rect 38669 67881 38703 67915
rect 38703 67881 38712 67915
rect 38660 67872 38712 67881
rect 39764 67872 39816 67924
rect 40960 67872 41012 67924
rect 42156 67915 42208 67924
rect 42156 67881 42165 67915
rect 42165 67881 42199 67915
rect 42199 67881 42208 67915
rect 42156 67872 42208 67881
rect 43260 67872 43312 67924
rect 69756 67915 69808 67924
rect 69756 67881 69765 67915
rect 69765 67881 69799 67915
rect 69799 67881 69808 67915
rect 69756 67872 69808 67881
rect 88340 67915 88392 67924
rect 88340 67881 88349 67915
rect 88349 67881 88383 67915
rect 88383 67881 88392 67915
rect 88340 67872 88392 67881
rect 88892 67915 88944 67924
rect 88892 67881 88901 67915
rect 88901 67881 88935 67915
rect 88935 67881 88944 67915
rect 88892 67872 88944 67881
rect 89168 67915 89220 67924
rect 89168 67881 89177 67915
rect 89177 67881 89211 67915
rect 89211 67881 89220 67915
rect 89168 67872 89220 67881
rect 90732 67872 90784 67924
rect 90824 67872 90876 67924
rect 94136 67872 94188 67924
rect 95056 67872 95108 67924
rect 97172 67915 97224 67924
rect 97172 67881 97181 67915
rect 97181 67881 97215 67915
rect 97215 67881 97224 67915
rect 97172 67872 97224 67881
rect 8392 67804 8444 67856
rect 90916 67847 90968 67856
rect 90916 67813 90925 67847
rect 90925 67813 90959 67847
rect 90959 67813 90968 67847
rect 90916 67804 90968 67813
rect 91008 67804 91060 67856
rect 10324 67736 10376 67788
rect 28080 67736 28132 67788
rect 90364 67779 90416 67788
rect 90364 67745 90373 67779
rect 90373 67745 90407 67779
rect 90407 67745 90416 67779
rect 90364 67736 90416 67745
rect 94964 67804 95016 67856
rect 29000 67711 29052 67720
rect 29000 67677 29009 67711
rect 29009 67677 29043 67711
rect 29043 67677 29052 67711
rect 29000 67668 29052 67677
rect 85672 67668 85724 67720
rect 87512 67711 87564 67720
rect 87512 67677 87521 67711
rect 87521 67677 87555 67711
rect 87555 67677 87564 67711
rect 87512 67668 87564 67677
rect 89076 67711 89128 67720
rect 89076 67677 89085 67711
rect 89085 67677 89119 67711
rect 89119 67677 89128 67711
rect 89076 67668 89128 67677
rect 1124 67600 1176 67652
rect 16396 67600 16448 67652
rect 22100 67600 22152 67652
rect 22376 67532 22428 67584
rect 86224 67600 86276 67652
rect 89812 67600 89864 67652
rect 91468 67668 91520 67720
rect 99196 67804 99248 67856
rect 108488 67847 108540 67856
rect 108488 67813 108497 67847
rect 108497 67813 108531 67847
rect 108531 67813 108540 67847
rect 108488 67804 108540 67813
rect 96988 67779 97040 67788
rect 96988 67745 96997 67779
rect 96997 67745 97031 67779
rect 97031 67745 97040 67779
rect 96988 67736 97040 67745
rect 102048 67736 102100 67788
rect 91744 67643 91796 67652
rect 91744 67609 91753 67643
rect 91753 67609 91787 67643
rect 91787 67609 91796 67643
rect 91744 67600 91796 67609
rect 31024 67532 31076 67584
rect 32864 67532 32916 67584
rect 38660 67532 38712 67584
rect 68284 67532 68336 67584
rect 69664 67532 69716 67584
rect 69848 67575 69900 67584
rect 69848 67541 69857 67575
rect 69857 67541 69891 67575
rect 69891 67541 69900 67575
rect 69848 67532 69900 67541
rect 89260 67532 89312 67584
rect 90640 67575 90692 67584
rect 90640 67541 90665 67575
rect 90665 67541 90692 67575
rect 90640 67532 90692 67541
rect 90824 67575 90876 67584
rect 90824 67541 90833 67575
rect 90833 67541 90867 67575
rect 90867 67541 90876 67575
rect 90824 67532 90876 67541
rect 90916 67532 90968 67584
rect 93400 67668 93452 67720
rect 92664 67643 92716 67652
rect 92664 67609 92673 67643
rect 92673 67609 92707 67643
rect 92707 67609 92716 67643
rect 92664 67600 92716 67609
rect 94136 67668 94188 67720
rect 93952 67600 94004 67652
rect 93676 67575 93728 67584
rect 93676 67541 93685 67575
rect 93685 67541 93719 67575
rect 93719 67541 93728 67575
rect 93676 67532 93728 67541
rect 93768 67532 93820 67584
rect 95056 67668 95108 67720
rect 95332 67711 95384 67720
rect 95332 67677 95341 67711
rect 95341 67677 95375 67711
rect 95375 67677 95384 67711
rect 95332 67668 95384 67677
rect 95608 67711 95660 67720
rect 95608 67677 95617 67711
rect 95617 67677 95651 67711
rect 95651 67677 95660 67711
rect 95608 67668 95660 67677
rect 96620 67711 96672 67720
rect 96620 67677 96629 67711
rect 96629 67677 96663 67711
rect 96663 67677 96672 67711
rect 96620 67668 96672 67677
rect 103612 67668 103664 67720
rect 103796 67668 103848 67720
rect 95700 67575 95752 67584
rect 95700 67541 95709 67575
rect 95709 67541 95743 67575
rect 95743 67541 95752 67575
rect 95700 67532 95752 67541
rect 95792 67575 95844 67584
rect 95792 67541 95801 67575
rect 95801 67541 95835 67575
rect 95835 67541 95844 67575
rect 95792 67532 95844 67541
rect 95976 67575 96028 67584
rect 95976 67541 95985 67575
rect 95985 67541 96019 67575
rect 96019 67541 96028 67575
rect 95976 67532 96028 67541
rect 98184 67532 98236 67584
rect 102600 67532 102652 67584
rect 4874 67430 4926 67482
rect 4938 67430 4990 67482
rect 5002 67430 5054 67482
rect 5066 67430 5118 67482
rect 5130 67430 5182 67482
rect 35594 67430 35646 67482
rect 35658 67430 35710 67482
rect 35722 67430 35774 67482
rect 35786 67430 35838 67482
rect 35850 67430 35902 67482
rect 66314 67430 66366 67482
rect 66378 67430 66430 67482
rect 66442 67430 66494 67482
rect 66506 67430 66558 67482
rect 66570 67430 66622 67482
rect 97034 67430 97086 67482
rect 97098 67430 97150 67482
rect 97162 67430 97214 67482
rect 97226 67430 97278 67482
rect 97290 67430 97342 67482
rect 106658 67430 106710 67482
rect 106722 67430 106774 67482
rect 106786 67430 106838 67482
rect 106850 67430 106902 67482
rect 106914 67430 106966 67482
rect 18880 67371 18932 67380
rect 18880 67337 18889 67371
rect 18889 67337 18923 67371
rect 18923 67337 18932 67371
rect 18880 67328 18932 67337
rect 24308 67260 24360 67312
rect 24676 67328 24728 67380
rect 35348 67371 35400 67380
rect 35348 67337 35357 67371
rect 35357 67337 35391 67371
rect 35391 67337 35400 67371
rect 35348 67328 35400 67337
rect 35992 67328 36044 67380
rect 38660 67371 38712 67380
rect 38660 67337 38669 67371
rect 38669 67337 38703 67371
rect 38703 67337 38712 67371
rect 38660 67328 38712 67337
rect 39948 67328 40000 67380
rect 47860 67328 47912 67380
rect 66996 67371 67048 67380
rect 66996 67337 67005 67371
rect 67005 67337 67039 67371
rect 67039 67337 67048 67371
rect 66996 67328 67048 67337
rect 69020 67328 69072 67380
rect 69756 67328 69808 67380
rect 70952 67371 71004 67380
rect 70952 67337 70961 67371
rect 70961 67337 70995 67371
rect 70995 67337 71004 67371
rect 70952 67328 71004 67337
rect 73988 67328 74040 67380
rect 75368 67371 75420 67380
rect 45744 67260 45796 67312
rect 46664 67303 46716 67312
rect 46664 67269 46673 67303
rect 46673 67269 46707 67303
rect 46707 67269 46716 67303
rect 46664 67260 46716 67269
rect 17316 67192 17368 67244
rect 29000 67192 29052 67244
rect 31208 67192 31260 67244
rect 32772 67192 32824 67244
rect 33508 67192 33560 67244
rect 33692 67235 33744 67244
rect 33692 67201 33701 67235
rect 33701 67201 33735 67235
rect 33735 67201 33744 67235
rect 33692 67192 33744 67201
rect 39028 67235 39080 67244
rect 39028 67201 39037 67235
rect 39037 67201 39071 67235
rect 39071 67201 39080 67235
rect 39028 67192 39080 67201
rect 20352 67124 20404 67176
rect 848 66988 900 67040
rect 20260 66988 20312 67040
rect 25044 67167 25096 67176
rect 25044 67133 25053 67167
rect 25053 67133 25087 67167
rect 25087 67133 25096 67167
rect 25044 67124 25096 67133
rect 29092 67124 29144 67176
rect 32956 67124 33008 67176
rect 34244 67124 34296 67176
rect 32864 67056 32916 67108
rect 39120 67167 39172 67176
rect 39120 67133 39129 67167
rect 39129 67133 39163 67167
rect 39163 67133 39172 67167
rect 39120 67124 39172 67133
rect 21272 67031 21324 67040
rect 21272 66997 21281 67031
rect 21281 66997 21315 67031
rect 21315 66997 21324 67031
rect 21272 66988 21324 66997
rect 22008 66988 22060 67040
rect 23296 67031 23348 67040
rect 23296 66997 23305 67031
rect 23305 66997 23339 67031
rect 23339 66997 23348 67031
rect 23296 66988 23348 66997
rect 25780 66988 25832 67040
rect 30564 67031 30616 67040
rect 30564 66997 30573 67031
rect 30573 66997 30607 67031
rect 30607 66997 30616 67031
rect 30564 66988 30616 66997
rect 31024 66988 31076 67040
rect 33508 66988 33560 67040
rect 40408 67167 40460 67176
rect 40408 67133 40417 67167
rect 40417 67133 40451 67167
rect 40451 67133 40460 67167
rect 40408 67124 40460 67133
rect 44456 67167 44508 67176
rect 44456 67133 44465 67167
rect 44465 67133 44499 67167
rect 44499 67133 44508 67167
rect 44456 67124 44508 67133
rect 47492 67192 47544 67244
rect 62396 67235 62448 67244
rect 62396 67201 62405 67235
rect 62405 67201 62439 67235
rect 62439 67201 62448 67235
rect 62396 67192 62448 67201
rect 68468 67303 68520 67312
rect 39396 67056 39448 67108
rect 39948 67031 40000 67040
rect 39948 66997 39957 67031
rect 39957 66997 39991 67031
rect 39991 66997 40000 67031
rect 39948 66988 40000 66997
rect 40408 66988 40460 67040
rect 43996 67031 44048 67040
rect 43996 66997 44005 67031
rect 44005 66997 44039 67031
rect 44039 66997 44048 67031
rect 43996 66988 44048 66997
rect 60740 67099 60792 67108
rect 60740 67065 60749 67099
rect 60749 67065 60783 67099
rect 60783 67065 60792 67099
rect 62212 67099 62264 67108
rect 60740 67056 60792 67065
rect 62212 67065 62221 67099
rect 62221 67065 62255 67099
rect 62255 67065 62264 67099
rect 62212 67056 62264 67065
rect 63408 67056 63460 67108
rect 68468 67269 68477 67303
rect 68477 67269 68511 67303
rect 68511 67269 68520 67303
rect 68468 67260 68520 67269
rect 68560 67235 68612 67244
rect 68560 67201 68569 67235
rect 68569 67201 68603 67235
rect 68603 67201 68612 67235
rect 68560 67192 68612 67201
rect 68284 67167 68336 67176
rect 68284 67133 68293 67167
rect 68293 67133 68327 67167
rect 68327 67133 68336 67167
rect 68284 67124 68336 67133
rect 75368 67337 75377 67371
rect 75377 67337 75411 67371
rect 75411 67337 75420 67371
rect 75368 67328 75420 67337
rect 75460 67371 75512 67380
rect 75460 67337 75469 67371
rect 75469 67337 75503 67371
rect 75503 67337 75512 67371
rect 75460 67328 75512 67337
rect 75828 67371 75880 67380
rect 75828 67337 75837 67371
rect 75837 67337 75871 67371
rect 75871 67337 75880 67371
rect 75828 67328 75880 67337
rect 89352 67328 89404 67380
rect 69480 67192 69532 67244
rect 71780 67235 71832 67244
rect 71780 67201 71789 67235
rect 71789 67201 71823 67235
rect 71823 67201 71832 67235
rect 71780 67192 71832 67201
rect 71872 67235 71924 67244
rect 71872 67201 71881 67235
rect 71881 67201 71915 67235
rect 71915 67201 71924 67235
rect 71872 67192 71924 67201
rect 73620 67235 73672 67244
rect 73620 67201 73629 67235
rect 73629 67201 73663 67235
rect 73663 67201 73672 67235
rect 73620 67192 73672 67201
rect 73712 67235 73764 67244
rect 73712 67201 73721 67235
rect 73721 67201 73755 67235
rect 73755 67201 73764 67235
rect 73712 67192 73764 67201
rect 67548 67056 67600 67108
rect 69756 67124 69808 67176
rect 69940 67167 69992 67176
rect 69940 67133 69949 67167
rect 69949 67133 69983 67167
rect 69983 67133 69992 67167
rect 69940 67124 69992 67133
rect 70032 67124 70084 67176
rect 75644 67192 75696 67244
rect 76196 67235 76248 67244
rect 76196 67201 76205 67235
rect 76205 67201 76239 67235
rect 76239 67201 76248 67235
rect 76196 67192 76248 67201
rect 77392 67192 77444 67244
rect 77576 67192 77628 67244
rect 86960 67192 87012 67244
rect 87512 67192 87564 67244
rect 88524 67192 88576 67244
rect 88616 67235 88668 67244
rect 88616 67201 88625 67235
rect 88625 67201 88659 67235
rect 88659 67201 88668 67235
rect 88616 67192 88668 67201
rect 89260 67235 89312 67244
rect 89260 67201 89269 67235
rect 89269 67201 89303 67235
rect 89303 67201 89312 67235
rect 89260 67192 89312 67201
rect 89536 67192 89588 67244
rect 70400 67056 70452 67108
rect 70584 67099 70636 67108
rect 70584 67065 70593 67099
rect 70593 67065 70627 67099
rect 70627 67065 70636 67099
rect 70584 67056 70636 67065
rect 85212 67124 85264 67176
rect 77944 67056 77996 67108
rect 66168 66988 66220 67040
rect 69480 67031 69532 67040
rect 69480 66997 69489 67031
rect 69489 66997 69523 67031
rect 69523 66997 69532 67031
rect 69480 66988 69532 66997
rect 75644 66988 75696 67040
rect 79784 66988 79836 67040
rect 79876 66988 79928 67040
rect 83096 66988 83148 67040
rect 85580 67167 85632 67176
rect 85580 67133 85589 67167
rect 85589 67133 85623 67167
rect 85623 67133 85632 67167
rect 85580 67124 85632 67133
rect 91560 67303 91612 67312
rect 91560 67269 91569 67303
rect 91569 67269 91603 67303
rect 91603 67269 91612 67303
rect 91560 67260 91612 67269
rect 92112 67328 92164 67380
rect 93308 67328 93360 67380
rect 95792 67328 95844 67380
rect 95884 67371 95936 67380
rect 95884 67337 95893 67371
rect 95893 67337 95927 67371
rect 95927 67337 95936 67371
rect 95884 67328 95936 67337
rect 96712 67328 96764 67380
rect 93584 67260 93636 67312
rect 92020 67235 92072 67244
rect 92020 67201 92029 67235
rect 92029 67201 92063 67235
rect 92063 67201 92072 67235
rect 92020 67192 92072 67201
rect 86224 66988 86276 67040
rect 88432 67056 88484 67108
rect 89812 67056 89864 67108
rect 87604 66988 87656 67040
rect 87788 66988 87840 67040
rect 89352 66988 89404 67040
rect 92020 66988 92072 67040
rect 92296 67167 92348 67176
rect 92296 67133 92305 67167
rect 92305 67133 92339 67167
rect 92339 67133 92348 67167
rect 92296 67124 92348 67133
rect 93768 67167 93820 67176
rect 93768 67133 93777 67167
rect 93777 67133 93811 67167
rect 93811 67133 93820 67167
rect 93768 67124 93820 67133
rect 93400 67056 93452 67108
rect 93676 66988 93728 67040
rect 94504 67124 94556 67176
rect 94780 67124 94832 67176
rect 96712 67192 96764 67244
rect 96804 67124 96856 67176
rect 96252 67031 96304 67040
rect 96252 66997 96261 67031
rect 96261 66997 96295 67031
rect 96295 66997 96304 67031
rect 96252 66988 96304 66997
rect 96712 66988 96764 67040
rect 98184 67260 98236 67312
rect 99380 67260 99432 67312
rect 99196 67235 99248 67244
rect 99196 67201 99205 67235
rect 99205 67201 99239 67235
rect 99239 67201 99248 67235
rect 99196 67192 99248 67201
rect 99748 67328 99800 67380
rect 102784 67328 102836 67380
rect 101772 67303 101824 67312
rect 101772 67269 101781 67303
rect 101781 67269 101815 67303
rect 101815 67269 101824 67303
rect 101772 67260 101824 67269
rect 101956 67303 102008 67312
rect 101956 67269 101965 67303
rect 101965 67269 101999 67303
rect 101999 67269 102008 67303
rect 101956 67260 102008 67269
rect 99564 67124 99616 67176
rect 103060 67056 103112 67108
rect 101864 66988 101916 67040
rect 106188 66988 106240 67040
rect 108488 67031 108540 67040
rect 108488 66997 108497 67031
rect 108497 66997 108531 67031
rect 108531 66997 108540 67031
rect 108488 66988 108540 66997
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 96374 66886 96426 66938
rect 96438 66886 96490 66938
rect 96502 66886 96554 66938
rect 96566 66886 96618 66938
rect 96630 66886 96682 66938
rect 2780 66784 2832 66836
rect 23296 66784 23348 66836
rect 24308 66784 24360 66836
rect 29736 66827 29788 66836
rect 29736 66793 29745 66827
rect 29745 66793 29779 66827
rect 29779 66793 29788 66827
rect 29736 66784 29788 66793
rect 43996 66784 44048 66836
rect 3424 66716 3476 66768
rect 18880 66716 18932 66768
rect 17316 66691 17368 66700
rect 17316 66657 17325 66691
rect 17325 66657 17359 66691
rect 17359 66657 17368 66691
rect 17316 66648 17368 66657
rect 19340 66648 19392 66700
rect 27068 66759 27120 66768
rect 27068 66725 27077 66759
rect 27077 66725 27111 66759
rect 27111 66725 27120 66759
rect 27068 66716 27120 66725
rect 21824 66512 21876 66564
rect 20260 66487 20312 66496
rect 20260 66453 20269 66487
rect 20269 66453 20303 66487
rect 20303 66453 20312 66487
rect 20260 66444 20312 66453
rect 20444 66487 20496 66496
rect 20444 66453 20453 66487
rect 20453 66453 20487 66487
rect 20487 66453 20496 66487
rect 20444 66444 20496 66453
rect 22008 66512 22060 66564
rect 25044 66648 25096 66700
rect 29092 66716 29144 66768
rect 32772 66759 32824 66768
rect 32772 66725 32781 66759
rect 32781 66725 32815 66759
rect 32815 66725 32824 66759
rect 32772 66716 32824 66725
rect 33048 66716 33100 66768
rect 34244 66759 34296 66768
rect 22376 66623 22428 66632
rect 22376 66589 22385 66623
rect 22385 66589 22419 66623
rect 22419 66589 22428 66623
rect 22376 66580 22428 66589
rect 25780 66580 25832 66632
rect 29000 66580 29052 66632
rect 24676 66555 24728 66564
rect 24676 66521 24685 66555
rect 24685 66521 24719 66555
rect 24719 66521 24728 66555
rect 24676 66512 24728 66521
rect 26148 66487 26200 66496
rect 26148 66453 26157 66487
rect 26157 66453 26191 66487
rect 26191 66453 26200 66487
rect 26148 66444 26200 66453
rect 30104 66487 30156 66496
rect 30104 66453 30113 66487
rect 30113 66453 30147 66487
rect 30147 66453 30156 66487
rect 30104 66444 30156 66453
rect 31024 66512 31076 66564
rect 33048 66623 33100 66632
rect 33048 66589 33057 66623
rect 33057 66589 33091 66623
rect 33091 66589 33100 66623
rect 33048 66580 33100 66589
rect 33600 66691 33652 66700
rect 33600 66657 33609 66691
rect 33609 66657 33643 66691
rect 33643 66657 33652 66691
rect 33600 66648 33652 66657
rect 34244 66725 34253 66759
rect 34253 66725 34287 66759
rect 34287 66725 34296 66759
rect 34244 66716 34296 66725
rect 53656 66716 53708 66768
rect 68560 66784 68612 66836
rect 75828 66784 75880 66836
rect 79876 66784 79928 66836
rect 80152 66784 80204 66836
rect 83096 66784 83148 66836
rect 33876 66648 33928 66700
rect 68284 66648 68336 66700
rect 70032 66648 70084 66700
rect 70952 66716 71004 66768
rect 71780 66716 71832 66768
rect 76196 66648 76248 66700
rect 35992 66580 36044 66632
rect 31944 66487 31996 66496
rect 31944 66453 31953 66487
rect 31953 66453 31987 66487
rect 31987 66453 31996 66487
rect 31944 66444 31996 66453
rect 32772 66444 32824 66496
rect 33600 66444 33652 66496
rect 57888 66444 57940 66496
rect 67640 66512 67692 66564
rect 69940 66512 69992 66564
rect 70308 66623 70360 66632
rect 70308 66589 70317 66623
rect 70317 66589 70351 66623
rect 70351 66589 70360 66623
rect 70308 66580 70360 66589
rect 70584 66580 70636 66632
rect 75920 66580 75972 66632
rect 77944 66580 77996 66632
rect 79968 66648 80020 66700
rect 83372 66648 83424 66700
rect 79784 66623 79836 66632
rect 79784 66589 79793 66623
rect 79793 66589 79827 66623
rect 79827 66589 79836 66623
rect 85672 66716 85724 66768
rect 84844 66691 84896 66700
rect 84844 66657 84853 66691
rect 84853 66657 84887 66691
rect 84887 66657 84896 66691
rect 84844 66648 84896 66657
rect 84660 66623 84712 66632
rect 79784 66580 79836 66589
rect 69296 66487 69348 66496
rect 69296 66453 69305 66487
rect 69305 66453 69339 66487
rect 69339 66453 69348 66487
rect 69296 66444 69348 66453
rect 69848 66444 69900 66496
rect 77576 66487 77628 66496
rect 77576 66453 77585 66487
rect 77585 66453 77619 66487
rect 77619 66453 77628 66487
rect 77576 66444 77628 66453
rect 80152 66487 80204 66496
rect 80152 66453 80161 66487
rect 80161 66453 80195 66487
rect 80195 66453 80204 66487
rect 80152 66444 80204 66453
rect 84660 66589 84669 66623
rect 84669 66589 84703 66623
rect 84703 66589 84712 66623
rect 84660 66580 84712 66589
rect 85396 66691 85448 66700
rect 85396 66657 85405 66691
rect 85405 66657 85439 66691
rect 85439 66657 85448 66691
rect 85396 66648 85448 66657
rect 86224 66691 86276 66700
rect 86224 66657 86233 66691
rect 86233 66657 86267 66691
rect 86267 66657 86276 66691
rect 88340 66784 88392 66836
rect 92020 66784 92072 66836
rect 94504 66784 94556 66836
rect 94964 66827 95016 66836
rect 94964 66793 94973 66827
rect 94973 66793 95007 66827
rect 95007 66793 95016 66827
rect 94964 66784 95016 66793
rect 96160 66827 96212 66836
rect 96160 66793 96169 66827
rect 96169 66793 96203 66827
rect 96203 66793 96212 66827
rect 96160 66784 96212 66793
rect 96252 66784 96304 66836
rect 99380 66784 99432 66836
rect 99472 66784 99524 66836
rect 104256 66784 104308 66836
rect 86224 66648 86276 66657
rect 88432 66648 88484 66700
rect 96068 66716 96120 66768
rect 96436 66716 96488 66768
rect 96712 66716 96764 66768
rect 104624 66716 104676 66768
rect 94044 66648 94096 66700
rect 89628 66580 89680 66632
rect 93216 66623 93268 66632
rect 93216 66589 93225 66623
rect 93225 66589 93259 66623
rect 93259 66589 93268 66623
rect 93216 66580 93268 66589
rect 85304 66512 85356 66564
rect 84936 66487 84988 66496
rect 84936 66453 84945 66487
rect 84945 66453 84979 66487
rect 84979 66453 84988 66487
rect 84936 66444 84988 66453
rect 87880 66444 87932 66496
rect 87972 66487 88024 66496
rect 87972 66453 87981 66487
rect 87981 66453 88015 66487
rect 88015 66453 88024 66487
rect 87972 66444 88024 66453
rect 88340 66512 88392 66564
rect 90272 66487 90324 66496
rect 90272 66453 90281 66487
rect 90281 66453 90315 66487
rect 90315 66453 90324 66487
rect 90272 66444 90324 66453
rect 90916 66444 90968 66496
rect 93032 66444 93084 66496
rect 93492 66555 93544 66564
rect 93492 66521 93501 66555
rect 93501 66521 93535 66555
rect 93535 66521 93544 66555
rect 93492 66512 93544 66521
rect 93584 66512 93636 66564
rect 94964 66512 95016 66564
rect 94872 66444 94924 66496
rect 96160 66580 96212 66632
rect 96620 66580 96672 66632
rect 98368 66580 98420 66632
rect 99472 66580 99524 66632
rect 95700 66512 95752 66564
rect 98276 66512 98328 66564
rect 95792 66487 95844 66496
rect 95792 66453 95801 66487
rect 95801 66453 95835 66487
rect 95835 66453 95844 66487
rect 95792 66444 95844 66453
rect 96160 66444 96212 66496
rect 96896 66444 96948 66496
rect 99748 66487 99800 66496
rect 99748 66453 99757 66487
rect 99757 66453 99791 66487
rect 99791 66453 99800 66487
rect 99748 66444 99800 66453
rect 101772 66623 101824 66632
rect 101772 66589 101781 66623
rect 101781 66589 101815 66623
rect 101815 66589 101824 66623
rect 101772 66580 101824 66589
rect 101864 66580 101916 66632
rect 102140 66623 102192 66632
rect 102140 66589 102149 66623
rect 102149 66589 102183 66623
rect 102183 66589 102192 66623
rect 102140 66580 102192 66589
rect 101956 66555 102008 66564
rect 101956 66521 101965 66555
rect 101965 66521 101999 66555
rect 101999 66521 102008 66555
rect 101956 66512 102008 66521
rect 104808 66444 104860 66496
rect 4874 66342 4926 66394
rect 4938 66342 4990 66394
rect 5002 66342 5054 66394
rect 5066 66342 5118 66394
rect 5130 66342 5182 66394
rect 35594 66342 35646 66394
rect 35658 66342 35710 66394
rect 35722 66342 35774 66394
rect 35786 66342 35838 66394
rect 35850 66342 35902 66394
rect 66314 66342 66366 66394
rect 66378 66342 66430 66394
rect 66442 66342 66494 66394
rect 66506 66342 66558 66394
rect 66570 66342 66622 66394
rect 97034 66342 97086 66394
rect 97098 66342 97150 66394
rect 97162 66342 97214 66394
rect 97226 66342 97278 66394
rect 97290 66342 97342 66394
rect 106658 66342 106710 66394
rect 106722 66342 106774 66394
rect 106786 66342 106838 66394
rect 106850 66342 106902 66394
rect 106914 66342 106966 66394
rect 9588 66240 9640 66292
rect 16396 66240 16448 66292
rect 20444 66240 20496 66292
rect 22008 66172 22060 66224
rect 16580 66104 16632 66156
rect 20260 66104 20312 66156
rect 21272 66104 21324 66156
rect 848 65900 900 65952
rect 23572 66104 23624 66156
rect 29092 66240 29144 66292
rect 30104 66240 30156 66292
rect 31944 66240 31996 66292
rect 32956 66240 33008 66292
rect 39396 66240 39448 66292
rect 70308 66240 70360 66292
rect 77576 66240 77628 66292
rect 80152 66240 80204 66292
rect 86960 66240 87012 66292
rect 23756 66172 23808 66224
rect 30564 66172 30616 66224
rect 31024 66215 31076 66224
rect 31024 66181 31033 66215
rect 31033 66181 31067 66215
rect 31067 66181 31076 66215
rect 31024 66172 31076 66181
rect 31208 66215 31260 66224
rect 31208 66181 31217 66215
rect 31217 66181 31251 66215
rect 31251 66181 31260 66215
rect 31208 66172 31260 66181
rect 57888 66172 57940 66224
rect 83372 66215 83424 66224
rect 83372 66181 83381 66215
rect 83381 66181 83415 66215
rect 83415 66181 83424 66215
rect 83372 66172 83424 66181
rect 88340 66240 88392 66292
rect 88432 66240 88484 66292
rect 89628 66240 89680 66292
rect 93308 66283 93360 66292
rect 93308 66249 93317 66283
rect 93317 66249 93351 66283
rect 93351 66249 93360 66283
rect 93308 66240 93360 66249
rect 22376 66036 22428 66088
rect 32772 66036 32824 66088
rect 60740 66104 60792 66156
rect 73988 66036 74040 66088
rect 86500 66104 86552 66156
rect 86224 66036 86276 66088
rect 88064 66104 88116 66156
rect 88432 66104 88484 66156
rect 88616 66104 88668 66156
rect 89076 66147 89128 66156
rect 89076 66113 89085 66147
rect 89085 66113 89119 66147
rect 89119 66113 89128 66147
rect 89076 66104 89128 66113
rect 89812 66172 89864 66224
rect 92940 66172 92992 66224
rect 93032 66172 93084 66224
rect 96712 66240 96764 66292
rect 98276 66283 98328 66292
rect 98276 66249 98285 66283
rect 98285 66249 98319 66283
rect 98319 66249 98328 66283
rect 98276 66240 98328 66249
rect 96068 66215 96120 66224
rect 96068 66181 96077 66215
rect 96077 66181 96111 66215
rect 96111 66181 96120 66215
rect 96068 66172 96120 66181
rect 96436 66172 96488 66224
rect 98368 66215 98420 66224
rect 98368 66181 98377 66215
rect 98377 66181 98411 66215
rect 98411 66181 98420 66215
rect 98368 66172 98420 66181
rect 86592 65968 86644 66020
rect 92664 66104 92716 66156
rect 90916 66036 90968 66088
rect 92296 66036 92348 66088
rect 53656 65943 53708 65952
rect 53656 65909 53665 65943
rect 53665 65909 53699 65943
rect 53699 65909 53708 65943
rect 53656 65900 53708 65909
rect 85580 65943 85632 65952
rect 85580 65909 85589 65943
rect 85589 65909 85623 65943
rect 85623 65909 85632 65943
rect 85580 65900 85632 65909
rect 86500 65943 86552 65952
rect 86500 65909 86509 65943
rect 86509 65909 86543 65943
rect 86543 65909 86552 65943
rect 86500 65900 86552 65909
rect 86776 65900 86828 65952
rect 88432 65943 88484 65952
rect 88432 65909 88441 65943
rect 88441 65909 88475 65943
rect 88475 65909 88484 65943
rect 88432 65900 88484 65909
rect 93492 66036 93544 66088
rect 93952 66147 94004 66156
rect 93952 66113 93961 66147
rect 93961 66113 93995 66147
rect 93995 66113 94004 66147
rect 93952 66104 94004 66113
rect 94504 66104 94556 66156
rect 96344 66147 96396 66156
rect 96344 66113 96353 66147
rect 96353 66113 96387 66147
rect 96387 66113 96396 66147
rect 99196 66240 99248 66292
rect 99380 66240 99432 66292
rect 99748 66172 99800 66224
rect 102140 66172 102192 66224
rect 96344 66104 96396 66113
rect 95976 66036 96028 66088
rect 100208 66147 100260 66156
rect 100208 66113 100217 66147
rect 100217 66113 100251 66147
rect 100251 66113 100260 66147
rect 100208 66104 100260 66113
rect 102048 66104 102100 66156
rect 108304 66147 108356 66156
rect 108304 66113 108313 66147
rect 108313 66113 108347 66147
rect 108347 66113 108356 66147
rect 108304 66104 108356 66113
rect 93952 65968 94004 66020
rect 94872 65968 94924 66020
rect 90272 65900 90324 65952
rect 91192 65943 91244 65952
rect 91192 65909 91201 65943
rect 91201 65909 91235 65943
rect 91235 65909 91244 65943
rect 91192 65900 91244 65909
rect 93032 65943 93084 65952
rect 93032 65909 93041 65943
rect 93041 65909 93075 65943
rect 93075 65909 93084 65943
rect 93032 65900 93084 65909
rect 93492 65943 93544 65952
rect 93492 65909 93501 65943
rect 93501 65909 93535 65943
rect 93535 65909 93544 65943
rect 93492 65900 93544 65909
rect 96620 65900 96672 65952
rect 96804 65943 96856 65952
rect 96804 65909 96834 65943
rect 96834 65909 96856 65943
rect 96804 65900 96856 65909
rect 98368 65943 98420 65952
rect 98368 65909 98377 65943
rect 98377 65909 98411 65943
rect 98411 65909 98420 65943
rect 98368 65900 98420 65909
rect 99564 65968 99616 66020
rect 100208 65900 100260 65952
rect 100576 65943 100628 65952
rect 100576 65909 100585 65943
rect 100585 65909 100619 65943
rect 100619 65909 100628 65943
rect 100576 65900 100628 65909
rect 108488 66011 108540 66020
rect 108488 65977 108497 66011
rect 108497 65977 108531 66011
rect 108531 65977 108540 66011
rect 108488 65968 108540 65977
rect 103796 65900 103848 65952
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 96374 65798 96426 65850
rect 96438 65798 96490 65850
rect 96502 65798 96554 65850
rect 96566 65798 96618 65850
rect 96630 65798 96682 65850
rect 105922 65798 105974 65850
rect 105986 65798 106038 65850
rect 106050 65798 106102 65850
rect 106114 65798 106166 65850
rect 106178 65798 106230 65850
rect 86960 65696 87012 65748
rect 93032 65696 93084 65748
rect 103888 65696 103940 65748
rect 87788 65628 87840 65680
rect 89628 65628 89680 65680
rect 91192 65628 91244 65680
rect 108304 65628 108356 65680
rect 75920 65560 75972 65612
rect 86500 65560 86552 65612
rect 88064 65560 88116 65612
rect 91744 65560 91796 65612
rect 100576 65560 100628 65612
rect 104164 65560 104216 65612
rect 30104 65492 30156 65544
rect 96712 65492 96764 65544
rect 85580 65424 85632 65476
rect 107568 65424 107620 65476
rect 848 65356 900 65408
rect 93492 65356 93544 65408
rect 104992 65356 105044 65408
rect 108488 65399 108540 65408
rect 108488 65365 108497 65399
rect 108497 65365 108531 65399
rect 108531 65365 108540 65399
rect 108488 65356 108540 65365
rect 4874 65254 4926 65306
rect 4938 65254 4990 65306
rect 5002 65254 5054 65306
rect 5066 65254 5118 65306
rect 5130 65254 5182 65306
rect 98368 65288 98420 65340
rect 103428 65288 103480 65340
rect 106658 65254 106710 65306
rect 106722 65254 106774 65306
rect 106786 65254 106838 65306
rect 106850 65254 106902 65306
rect 106914 65254 106966 65306
rect 96068 65152 96120 65204
rect 104440 65152 104492 65204
rect 1400 64923 1452 64932
rect 1400 64889 1409 64923
rect 1409 64889 1443 64923
rect 1443 64889 1452 64923
rect 1400 64880 1452 64889
rect 87604 65016 87656 65068
rect 26148 64880 26200 64932
rect 108488 64923 108540 64932
rect 108488 64889 108497 64923
rect 108497 64889 108531 64923
rect 108531 64889 108540 64923
rect 108488 64880 108540 64889
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 105922 64710 105974 64762
rect 105986 64710 106038 64762
rect 106050 64710 106102 64762
rect 106114 64710 106166 64762
rect 106178 64710 106230 64762
rect 22008 64404 22060 64456
rect 88524 64404 88576 64456
rect 848 64268 900 64320
rect 1860 64268 1912 64320
rect 10324 64268 10376 64320
rect 108488 64311 108540 64320
rect 108488 64277 108497 64311
rect 108497 64277 108531 64311
rect 108531 64277 108540 64311
rect 108488 64268 108540 64277
rect 4874 64166 4926 64218
rect 4938 64166 4990 64218
rect 5002 64166 5054 64218
rect 5066 64166 5118 64218
rect 5130 64166 5182 64218
rect 77392 64132 77444 64184
rect 102784 64132 102836 64184
rect 106658 64166 106710 64218
rect 106722 64166 106774 64218
rect 106786 64166 106838 64218
rect 106850 64166 106902 64218
rect 106914 64166 106966 64218
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 105922 63622 105974 63674
rect 105986 63622 106038 63674
rect 106050 63622 106102 63674
rect 106114 63622 106166 63674
rect 106178 63622 106230 63674
rect 848 63452 900 63504
rect 2780 63452 2832 63504
rect 4874 63078 4926 63130
rect 4938 63078 4990 63130
rect 5002 63078 5054 63130
rect 5066 63078 5118 63130
rect 5130 63078 5182 63130
rect 106658 63078 106710 63130
rect 106722 63078 106774 63130
rect 106786 63078 106838 63130
rect 106850 63078 106902 63130
rect 106914 63078 106966 63130
rect 3424 62976 3476 63028
rect 848 62704 900 62756
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 105922 62534 105974 62586
rect 105986 62534 106038 62586
rect 106050 62534 106102 62586
rect 106114 62534 106166 62586
rect 106178 62534 106230 62586
rect 1860 62475 1912 62484
rect 1860 62441 1869 62475
rect 1869 62441 1903 62475
rect 1903 62441 1912 62475
rect 1860 62432 1912 62441
rect 1492 62203 1544 62212
rect 1492 62169 1501 62203
rect 1501 62169 1535 62203
rect 1535 62169 1544 62203
rect 1492 62160 1544 62169
rect 4874 61990 4926 62042
rect 4938 61990 4990 62042
rect 5002 61990 5054 62042
rect 5066 61990 5118 62042
rect 5130 61990 5182 62042
rect 106658 61990 106710 62042
rect 106722 61990 106774 62042
rect 106786 61990 106838 62042
rect 106850 61990 106902 62042
rect 106914 61990 106966 62042
rect 1676 61863 1728 61872
rect 1676 61829 1685 61863
rect 1685 61829 1719 61863
rect 1719 61829 1728 61863
rect 1676 61820 1728 61829
rect 1308 61752 1360 61804
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 105922 61446 105974 61498
rect 105986 61446 106038 61498
rect 106050 61446 106102 61498
rect 106114 61446 106166 61498
rect 106178 61446 106230 61498
rect 4874 60902 4926 60954
rect 4938 60902 4990 60954
rect 5002 60902 5054 60954
rect 5066 60902 5118 60954
rect 5130 60902 5182 60954
rect 106658 60902 106710 60954
rect 106722 60902 106774 60954
rect 106786 60902 106838 60954
rect 106850 60902 106902 60954
rect 106914 60902 106966 60954
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 105922 60358 105974 60410
rect 105986 60358 106038 60410
rect 106050 60358 106102 60410
rect 106114 60358 106166 60410
rect 106178 60358 106230 60410
rect 103980 60052 104032 60104
rect 4874 59814 4926 59866
rect 4938 59814 4990 59866
rect 5002 59814 5054 59866
rect 5066 59814 5118 59866
rect 5130 59814 5182 59866
rect 106658 59814 106710 59866
rect 106722 59814 106774 59866
rect 106786 59814 106838 59866
rect 106850 59814 106902 59866
rect 106914 59814 106966 59866
rect 104440 59755 104492 59764
rect 104440 59721 104449 59755
rect 104449 59721 104483 59755
rect 104483 59721 104492 59755
rect 104440 59712 104492 59721
rect 103428 59576 103480 59628
rect 103980 59508 104032 59560
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 105922 59270 105974 59322
rect 105986 59270 106038 59322
rect 106050 59270 106102 59322
rect 106114 59270 106166 59322
rect 106178 59270 106230 59322
rect 4874 58726 4926 58778
rect 4938 58726 4990 58778
rect 5002 58726 5054 58778
rect 5066 58726 5118 58778
rect 5130 58726 5182 58778
rect 106658 58726 106710 58778
rect 106722 58726 106774 58778
rect 106786 58726 106838 58778
rect 106850 58726 106902 58778
rect 106914 58726 106966 58778
rect 105636 58667 105688 58676
rect 105636 58633 105645 58667
rect 105645 58633 105679 58667
rect 105679 58633 105688 58667
rect 105636 58624 105688 58633
rect 105820 58624 105872 58676
rect 104348 58599 104400 58608
rect 104348 58565 104357 58599
rect 104357 58565 104391 58599
rect 104391 58565 104400 58599
rect 104348 58556 104400 58565
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 105922 58182 105974 58234
rect 105986 58182 106038 58234
rect 106050 58182 106102 58234
rect 106114 58182 106166 58234
rect 106178 58182 106230 58234
rect 104348 58123 104400 58132
rect 104348 58089 104357 58123
rect 104357 58089 104391 58123
rect 104391 58089 104400 58123
rect 104348 58080 104400 58089
rect 4874 57638 4926 57690
rect 4938 57638 4990 57690
rect 5002 57638 5054 57690
rect 5066 57638 5118 57690
rect 5130 57638 5182 57690
rect 106658 57638 106710 57690
rect 106722 57638 106774 57690
rect 106786 57638 106838 57690
rect 106850 57638 106902 57690
rect 106914 57638 106966 57690
rect 104256 57536 104308 57588
rect 104532 57579 104584 57588
rect 104532 57545 104541 57579
rect 104541 57545 104575 57579
rect 104575 57545 104584 57579
rect 104532 57536 104584 57545
rect 103796 57468 103848 57520
rect 104716 57468 104768 57520
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 105922 57094 105974 57146
rect 105986 57094 106038 57146
rect 106050 57094 106102 57146
rect 106114 57094 106166 57146
rect 106178 57094 106230 57146
rect 104992 57035 105044 57044
rect 104992 57001 105001 57035
rect 105001 57001 105035 57035
rect 105035 57001 105044 57035
rect 104992 56992 105044 57001
rect 104164 56856 104216 56908
rect 104440 56856 104492 56908
rect 104716 56899 104768 56908
rect 104716 56865 104725 56899
rect 104725 56865 104759 56899
rect 104759 56865 104768 56899
rect 104716 56856 104768 56865
rect 104808 56899 104860 56908
rect 104808 56865 104817 56899
rect 104817 56865 104851 56899
rect 104851 56865 104860 56899
rect 104808 56856 104860 56865
rect 104256 56788 104308 56840
rect 104348 56652 104400 56704
rect 104532 56695 104584 56704
rect 104532 56661 104541 56695
rect 104541 56661 104575 56695
rect 104575 56661 104584 56695
rect 104532 56652 104584 56661
rect 4874 56550 4926 56602
rect 4938 56550 4990 56602
rect 5002 56550 5054 56602
rect 5066 56550 5118 56602
rect 5130 56550 5182 56602
rect 106658 56550 106710 56602
rect 106722 56550 106774 56602
rect 106786 56550 106838 56602
rect 106850 56550 106902 56602
rect 106914 56550 106966 56602
rect 104164 56448 104216 56500
rect 104716 56491 104768 56500
rect 104716 56457 104725 56491
rect 104725 56457 104759 56491
rect 104759 56457 104768 56491
rect 104716 56448 104768 56457
rect 104624 56423 104676 56432
rect 104624 56389 104633 56423
rect 104633 56389 104667 56423
rect 104667 56389 104676 56423
rect 104624 56380 104676 56389
rect 104348 56312 104400 56364
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 105922 56006 105974 56058
rect 105986 56006 106038 56058
rect 106050 56006 106102 56058
rect 106114 56006 106166 56058
rect 106178 56006 106230 56058
rect 4874 55462 4926 55514
rect 4938 55462 4990 55514
rect 5002 55462 5054 55514
rect 5066 55462 5118 55514
rect 5130 55462 5182 55514
rect 106658 55462 106710 55514
rect 106722 55462 106774 55514
rect 106786 55462 106838 55514
rect 106850 55462 106902 55514
rect 106914 55462 106966 55514
rect 103796 55360 103848 55412
rect 104532 55292 104584 55344
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 105922 54918 105974 54970
rect 105986 54918 106038 54970
rect 106050 54918 106102 54970
rect 106114 54918 106166 54970
rect 106178 54918 106230 54970
rect 103888 54816 103940 54868
rect 104440 54748 104492 54800
rect 104532 54655 104584 54664
rect 104532 54621 104541 54655
rect 104541 54621 104575 54655
rect 104575 54621 104584 54655
rect 104532 54612 104584 54621
rect 104624 54519 104676 54528
rect 104624 54485 104633 54519
rect 104633 54485 104667 54519
rect 104667 54485 104676 54519
rect 104624 54476 104676 54485
rect 104716 54519 104768 54528
rect 104716 54485 104725 54519
rect 104725 54485 104759 54519
rect 104759 54485 104768 54519
rect 104716 54476 104768 54485
rect 4874 54374 4926 54426
rect 4938 54374 4990 54426
rect 5002 54374 5054 54426
rect 5066 54374 5118 54426
rect 5130 54374 5182 54426
rect 106658 54374 106710 54426
rect 106722 54374 106774 54426
rect 106786 54374 106838 54426
rect 106850 54374 106902 54426
rect 106914 54374 106966 54426
rect 104440 54315 104492 54324
rect 104440 54281 104449 54315
rect 104449 54281 104483 54315
rect 104483 54281 104492 54315
rect 104440 54272 104492 54281
rect 104532 54315 104584 54324
rect 104532 54281 104541 54315
rect 104541 54281 104575 54315
rect 104575 54281 104584 54315
rect 104532 54272 104584 54281
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 105922 53830 105974 53882
rect 105986 53830 106038 53882
rect 106050 53830 106102 53882
rect 106114 53830 106166 53882
rect 106178 53830 106230 53882
rect 4874 53286 4926 53338
rect 4938 53286 4990 53338
rect 5002 53286 5054 53338
rect 5066 53286 5118 53338
rect 5130 53286 5182 53338
rect 106658 53286 106710 53338
rect 106722 53286 106774 53338
rect 106786 53286 106838 53338
rect 106850 53286 106902 53338
rect 106914 53286 106966 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 105922 52742 105974 52794
rect 105986 52742 106038 52794
rect 106050 52742 106102 52794
rect 106114 52742 106166 52794
rect 106178 52742 106230 52794
rect 4874 52198 4926 52250
rect 4938 52198 4990 52250
rect 5002 52198 5054 52250
rect 5066 52198 5118 52250
rect 5130 52198 5182 52250
rect 106658 52198 106710 52250
rect 106722 52198 106774 52250
rect 106786 52198 106838 52250
rect 106850 52198 106902 52250
rect 106914 52198 106966 52250
rect 104532 52096 104584 52148
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 105922 51654 105974 51706
rect 105986 51654 106038 51706
rect 106050 51654 106102 51706
rect 106114 51654 106166 51706
rect 106178 51654 106230 51706
rect 104532 51595 104584 51604
rect 104532 51561 104541 51595
rect 104541 51561 104575 51595
rect 104575 51561 104584 51595
rect 104532 51552 104584 51561
rect 103980 51484 104032 51536
rect 104624 51348 104676 51400
rect 104440 51280 104492 51332
rect 108488 51391 108540 51400
rect 108488 51357 108497 51391
rect 108497 51357 108531 51391
rect 108531 51357 108540 51391
rect 108488 51348 108540 51357
rect 104532 51255 104584 51264
rect 104532 51221 104557 51255
rect 104557 51221 104584 51255
rect 104532 51212 104584 51221
rect 105360 51255 105412 51264
rect 105360 51221 105369 51255
rect 105369 51221 105403 51255
rect 105403 51221 105412 51255
rect 105360 51212 105412 51221
rect 108304 51255 108356 51264
rect 108304 51221 108313 51255
rect 108313 51221 108347 51255
rect 108347 51221 108356 51255
rect 108304 51212 108356 51221
rect 4874 51110 4926 51162
rect 4938 51110 4990 51162
rect 5002 51110 5054 51162
rect 5066 51110 5118 51162
rect 5130 51110 5182 51162
rect 106658 51110 106710 51162
rect 106722 51110 106774 51162
rect 106786 51110 106838 51162
rect 106850 51110 106902 51162
rect 106914 51110 106966 51162
rect 104440 51051 104492 51060
rect 104440 51017 104449 51051
rect 104449 51017 104483 51051
rect 104483 51017 104492 51051
rect 104440 51008 104492 51017
rect 104532 51051 104584 51060
rect 104532 51017 104541 51051
rect 104541 51017 104575 51051
rect 104575 51017 104584 51051
rect 104532 51008 104584 51017
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 105922 50566 105974 50618
rect 105986 50566 106038 50618
rect 106050 50566 106102 50618
rect 106114 50566 106166 50618
rect 106178 50566 106230 50618
rect 4874 50022 4926 50074
rect 4938 50022 4990 50074
rect 5002 50022 5054 50074
rect 5066 50022 5118 50074
rect 5130 50022 5182 50074
rect 106658 50022 106710 50074
rect 106722 50022 106774 50074
rect 106786 50022 106838 50074
rect 106850 50022 106902 50074
rect 106914 50022 106966 50074
rect 104716 49963 104768 49972
rect 104716 49929 104725 49963
rect 104725 49929 104759 49963
rect 104759 49929 104768 49963
rect 104716 49920 104768 49929
rect 104256 49852 104308 49904
rect 104348 49827 104400 49836
rect 104348 49793 104357 49827
rect 104357 49793 104391 49827
rect 104391 49793 104400 49827
rect 104348 49784 104400 49793
rect 104808 49759 104860 49768
rect 104808 49725 104817 49759
rect 104817 49725 104851 49759
rect 104851 49725 104860 49759
rect 104808 49716 104860 49725
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 105922 49478 105974 49530
rect 105986 49478 106038 49530
rect 106050 49478 106102 49530
rect 106114 49478 106166 49530
rect 106178 49478 106230 49530
rect 104256 49376 104308 49428
rect 4874 48934 4926 48986
rect 4938 48934 4990 48986
rect 5002 48934 5054 48986
rect 5066 48934 5118 48986
rect 5130 48934 5182 48986
rect 106658 48934 106710 48986
rect 106722 48934 106774 48986
rect 106786 48934 106838 48986
rect 106850 48934 106902 48986
rect 106914 48934 106966 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 105922 48390 105974 48442
rect 105986 48390 106038 48442
rect 106050 48390 106102 48442
rect 106114 48390 106166 48442
rect 106178 48390 106230 48442
rect 4874 47846 4926 47898
rect 4938 47846 4990 47898
rect 5002 47846 5054 47898
rect 5066 47846 5118 47898
rect 5130 47846 5182 47898
rect 106658 47846 106710 47898
rect 106722 47846 106774 47898
rect 106786 47846 106838 47898
rect 106850 47846 106902 47898
rect 106914 47846 106966 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 105922 47302 105974 47354
rect 105986 47302 106038 47354
rect 106050 47302 106102 47354
rect 106114 47302 106166 47354
rect 106178 47302 106230 47354
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 106658 46758 106710 46810
rect 106722 46758 106774 46810
rect 106786 46758 106838 46810
rect 106850 46758 106902 46810
rect 106914 46758 106966 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 105922 46214 105974 46266
rect 105986 46214 106038 46266
rect 106050 46214 106102 46266
rect 106114 46214 106166 46266
rect 106178 46214 106230 46266
rect 104348 46155 104400 46164
rect 104348 46121 104357 46155
rect 104357 46121 104391 46155
rect 104391 46121 104400 46155
rect 104348 46112 104400 46121
rect 104256 45908 104308 45960
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 106658 45670 106710 45722
rect 106722 45670 106774 45722
rect 106786 45670 106838 45722
rect 106850 45670 106902 45722
rect 106914 45670 106966 45722
rect 105084 45432 105136 45484
rect 104624 45407 104676 45416
rect 104624 45373 104633 45407
rect 104633 45373 104667 45407
rect 104667 45373 104676 45407
rect 104624 45364 104676 45373
rect 105176 45228 105228 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 105922 45126 105974 45178
rect 105986 45126 106038 45178
rect 106050 45126 106102 45178
rect 106114 45126 106166 45178
rect 106178 45126 106230 45178
rect 102784 44888 102836 44940
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 108304 44820 108356 44872
rect 106658 44582 106710 44634
rect 106722 44582 106774 44634
rect 106786 44582 106838 44634
rect 106850 44582 106902 44634
rect 106914 44582 106966 44634
rect 103704 44276 103756 44328
rect 104716 44140 104768 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 105922 44038 105974 44090
rect 105986 44038 106038 44090
rect 106050 44038 106102 44090
rect 106114 44038 106166 44090
rect 106178 44038 106230 44090
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 106658 43494 106710 43546
rect 106722 43494 106774 43546
rect 106786 43494 106838 43546
rect 106850 43494 106902 43546
rect 106914 43494 106966 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 105922 42950 105974 43002
rect 105986 42950 106038 43002
rect 106050 42950 106102 43002
rect 106114 42950 106166 43002
rect 106178 42950 106230 43002
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 106658 42406 106710 42458
rect 106722 42406 106774 42458
rect 106786 42406 106838 42458
rect 106850 42406 106902 42458
rect 106914 42406 106966 42458
rect 105084 42347 105136 42356
rect 105084 42313 105093 42347
rect 105093 42313 105127 42347
rect 105127 42313 105136 42347
rect 105084 42304 105136 42313
rect 104256 42168 104308 42220
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 105922 41862 105974 41914
rect 105986 41862 106038 41914
rect 106050 41862 106102 41914
rect 106114 41862 106166 41914
rect 106178 41862 106230 41914
rect 5540 41692 5592 41744
rect 1216 41556 1268 41608
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 106658 41318 106710 41370
rect 106722 41318 106774 41370
rect 106786 41318 106838 41370
rect 106850 41318 106902 41370
rect 106914 41318 106966 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 105922 40774 105974 40826
rect 105986 40774 106038 40826
rect 106050 40774 106102 40826
rect 106114 40774 106166 40826
rect 106178 40774 106230 40826
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 106658 40230 106710 40282
rect 106722 40230 106774 40282
rect 106786 40230 106838 40282
rect 106850 40230 106902 40282
rect 106914 40230 106966 40282
rect 5540 40128 5592 40180
rect 1400 40035 1452 40044
rect 1400 40001 1409 40035
rect 1409 40001 1443 40035
rect 1443 40001 1452 40035
rect 1400 39992 1452 40001
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 105922 39686 105974 39738
rect 105986 39686 106038 39738
rect 106050 39686 106102 39738
rect 106114 39686 106166 39738
rect 106178 39686 106230 39738
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 106658 39142 106710 39194
rect 106722 39142 106774 39194
rect 106786 39142 106838 39194
rect 106850 39142 106902 39194
rect 106914 39142 106966 39194
rect 104348 38836 104400 38888
rect 105360 38836 105412 38888
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 105922 38598 105974 38650
rect 105986 38598 106038 38650
rect 106050 38598 106102 38650
rect 106114 38598 106166 38650
rect 106178 38598 106230 38650
rect 8392 38428 8444 38480
rect 1216 38292 1268 38344
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 106658 38054 106710 38106
rect 106722 38054 106774 38106
rect 106786 38054 106838 38106
rect 106850 38054 106902 38106
rect 106914 38054 106966 38106
rect 104256 37952 104308 38004
rect 105820 37952 105872 38004
rect 104716 37816 104768 37868
rect 105176 37748 105228 37800
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 105922 37510 105974 37562
rect 105986 37510 106038 37562
rect 106050 37510 106102 37562
rect 106114 37510 106166 37562
rect 106178 37510 106230 37562
rect 104716 37315 104768 37324
rect 104716 37281 104725 37315
rect 104725 37281 104759 37315
rect 104759 37281 104768 37315
rect 104716 37272 104768 37281
rect 1400 37247 1452 37256
rect 1400 37213 1409 37247
rect 1409 37213 1443 37247
rect 1443 37213 1452 37247
rect 1400 37204 1452 37213
rect 104256 37204 104308 37256
rect 9496 37136 9548 37188
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 106658 36966 106710 37018
rect 106722 36966 106774 37018
rect 106786 36966 106838 37018
rect 106850 36966 106902 37018
rect 106914 36966 106966 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 105922 36422 105974 36474
rect 105986 36422 106038 36474
rect 106050 36422 106102 36474
rect 106114 36422 106166 36474
rect 106178 36422 106230 36474
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 106658 35878 106710 35930
rect 106722 35878 106774 35930
rect 106786 35878 106838 35930
rect 106850 35878 106902 35930
rect 106914 35878 106966 35930
rect 9496 35776 9548 35828
rect 1308 35640 1360 35692
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 105922 35334 105974 35386
rect 105986 35334 106038 35386
rect 106050 35334 106102 35386
rect 106114 35334 106166 35386
rect 106178 35334 106230 35386
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 106658 34790 106710 34842
rect 106722 34790 106774 34842
rect 106786 34790 106838 34842
rect 106850 34790 106902 34842
rect 106914 34790 106966 34842
rect 5540 34688 5592 34740
rect 1400 34595 1452 34604
rect 1400 34561 1409 34595
rect 1409 34561 1443 34595
rect 1443 34561 1452 34595
rect 1400 34552 1452 34561
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 105922 34246 105974 34298
rect 105986 34246 106038 34298
rect 106050 34246 106102 34298
rect 106114 34246 106166 34298
rect 106178 34246 106230 34298
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 106658 33702 106710 33754
rect 106722 33702 106774 33754
rect 106786 33702 106838 33754
rect 106850 33702 106902 33754
rect 106914 33702 106966 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 105922 33158 105974 33210
rect 105986 33158 106038 33210
rect 106050 33158 106102 33210
rect 106114 33158 106166 33210
rect 106178 33158 106230 33210
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 106658 32614 106710 32666
rect 106722 32614 106774 32666
rect 106786 32614 106838 32666
rect 106850 32614 106902 32666
rect 106914 32614 106966 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 105922 32070 105974 32122
rect 105986 32070 106038 32122
rect 106050 32070 106102 32122
rect 106114 32070 106166 32122
rect 106178 32070 106230 32122
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 106658 31526 106710 31578
rect 106722 31526 106774 31578
rect 106786 31526 106838 31578
rect 106850 31526 106902 31578
rect 106914 31526 106966 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 105922 30982 105974 31034
rect 105986 30982 106038 31034
rect 106050 30982 106102 31034
rect 106114 30982 106166 31034
rect 106178 30982 106230 31034
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 106658 30438 106710 30490
rect 106722 30438 106774 30490
rect 106786 30438 106838 30490
rect 106850 30438 106902 30490
rect 106914 30438 106966 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 105922 29894 105974 29946
rect 105986 29894 106038 29946
rect 106050 29894 106102 29946
rect 106114 29894 106166 29946
rect 106178 29894 106230 29946
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 106658 29350 106710 29402
rect 106722 29350 106774 29402
rect 106786 29350 106838 29402
rect 106850 29350 106902 29402
rect 106914 29350 106966 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 105922 28806 105974 28858
rect 105986 28806 106038 28858
rect 106050 28806 106102 28858
rect 106114 28806 106166 28858
rect 106178 28806 106230 28858
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 106658 28262 106710 28314
rect 106722 28262 106774 28314
rect 106786 28262 106838 28314
rect 106850 28262 106902 28314
rect 106914 28262 106966 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 105922 27718 105974 27770
rect 105986 27718 106038 27770
rect 106050 27718 106102 27770
rect 106114 27718 106166 27770
rect 106178 27718 106230 27770
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 106658 27174 106710 27226
rect 106722 27174 106774 27226
rect 106786 27174 106838 27226
rect 106850 27174 106902 27226
rect 106914 27174 106966 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 105922 26630 105974 26682
rect 105986 26630 106038 26682
rect 106050 26630 106102 26682
rect 106114 26630 106166 26682
rect 106178 26630 106230 26682
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 106658 26086 106710 26138
rect 106722 26086 106774 26138
rect 106786 26086 106838 26138
rect 106850 26086 106902 26138
rect 106914 26086 106966 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 105922 25542 105974 25594
rect 105986 25542 106038 25594
rect 106050 25542 106102 25594
rect 106114 25542 106166 25594
rect 106178 25542 106230 25594
rect 102600 25100 102652 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 106658 24998 106710 25050
rect 106722 24998 106774 25050
rect 106786 24998 106838 25050
rect 106850 24998 106902 25050
rect 106914 24998 106966 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 105922 24454 105974 24506
rect 105986 24454 106038 24506
rect 106050 24454 106102 24506
rect 106114 24454 106166 24506
rect 106178 24454 106230 24506
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 106658 23910 106710 23962
rect 106722 23910 106774 23962
rect 106786 23910 106838 23962
rect 106850 23910 106902 23962
rect 106914 23910 106966 23962
rect 101956 23808 102008 23860
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 105922 23366 105974 23418
rect 105986 23366 106038 23418
rect 106050 23366 106102 23418
rect 106114 23366 106166 23418
rect 106178 23366 106230 23418
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 106658 22822 106710 22874
rect 106722 22822 106774 22874
rect 106786 22822 106838 22874
rect 106850 22822 106902 22874
rect 106914 22822 106966 22874
rect 104348 22763 104400 22772
rect 104348 22729 104357 22763
rect 104357 22729 104391 22763
rect 104391 22729 104400 22763
rect 104348 22720 104400 22729
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 105922 22278 105974 22330
rect 105986 22278 106038 22330
rect 106050 22278 106102 22330
rect 106114 22278 106166 22330
rect 106178 22278 106230 22330
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 106658 21734 106710 21786
rect 106722 21734 106774 21786
rect 106786 21734 106838 21786
rect 106850 21734 106902 21786
rect 106914 21734 106966 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 105922 21190 105974 21242
rect 105986 21190 106038 21242
rect 106050 21190 106102 21242
rect 106114 21190 106166 21242
rect 106178 21190 106230 21242
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 106658 20646 106710 20698
rect 106722 20646 106774 20698
rect 106786 20646 106838 20698
rect 106850 20646 106902 20698
rect 106914 20646 106966 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 105922 20102 105974 20154
rect 105986 20102 106038 20154
rect 106050 20102 106102 20154
rect 106114 20102 106166 20154
rect 106178 20102 106230 20154
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 106658 19558 106710 19610
rect 106722 19558 106774 19610
rect 106786 19558 106838 19610
rect 106850 19558 106902 19610
rect 106914 19558 106966 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 105922 19014 105974 19066
rect 105986 19014 106038 19066
rect 106050 19014 106102 19066
rect 106114 19014 106166 19066
rect 106178 19014 106230 19066
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 106658 18470 106710 18522
rect 106722 18470 106774 18522
rect 106786 18470 106838 18522
rect 106850 18470 106902 18522
rect 106914 18470 106966 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 105922 17926 105974 17978
rect 105986 17926 106038 17978
rect 106050 17926 106102 17978
rect 106114 17926 106166 17978
rect 106178 17926 106230 17978
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 106658 17382 106710 17434
rect 106722 17382 106774 17434
rect 106786 17382 106838 17434
rect 106850 17382 106902 17434
rect 106914 17382 106966 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 105922 16838 105974 16890
rect 105986 16838 106038 16890
rect 106050 16838 106102 16890
rect 106114 16838 106166 16890
rect 106178 16838 106230 16890
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 106658 16294 106710 16346
rect 106722 16294 106774 16346
rect 106786 16294 106838 16346
rect 106850 16294 106902 16346
rect 106914 16294 106966 16346
rect 1308 16056 1360 16108
rect 9496 15920 9548 15972
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 105922 15750 105974 15802
rect 105986 15750 106038 15802
rect 106050 15750 106102 15802
rect 106114 15750 106166 15802
rect 106178 15750 106230 15802
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 106658 15206 106710 15258
rect 106722 15206 106774 15258
rect 106786 15206 106838 15258
rect 106850 15206 106902 15258
rect 106914 15206 106966 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 105922 14662 105974 14714
rect 105986 14662 106038 14714
rect 106050 14662 106102 14714
rect 106114 14662 106166 14714
rect 106178 14662 106230 14714
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 106658 14118 106710 14170
rect 106722 14118 106774 14170
rect 106786 14118 106838 14170
rect 106850 14118 106902 14170
rect 106914 14118 106966 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 105922 13574 105974 13626
rect 105986 13574 106038 13626
rect 106050 13574 106102 13626
rect 106114 13574 106166 13626
rect 106178 13574 106230 13626
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 106658 13030 106710 13082
rect 106722 13030 106774 13082
rect 106786 13030 106838 13082
rect 106850 13030 106902 13082
rect 106914 13030 106966 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 105922 12486 105974 12538
rect 105986 12486 106038 12538
rect 106050 12486 106102 12538
rect 106114 12486 106166 12538
rect 106178 12486 106230 12538
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 106658 11942 106710 11994
rect 106722 11942 106774 11994
rect 106786 11942 106838 11994
rect 106850 11942 106902 11994
rect 106914 11942 106966 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 105922 11398 105974 11450
rect 105986 11398 106038 11450
rect 106050 11398 106102 11450
rect 106114 11398 106166 11450
rect 106178 11398 106230 11450
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 106658 10854 106710 10906
rect 106722 10854 106774 10906
rect 106786 10854 106838 10906
rect 106850 10854 106902 10906
rect 106914 10854 106966 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 105922 10310 105974 10362
rect 105986 10310 106038 10362
rect 106050 10310 106102 10362
rect 106114 10310 106166 10362
rect 106178 10310 106230 10362
rect 90732 10004 90784 10056
rect 104716 10004 104768 10056
rect 90824 9936 90876 9988
rect 103796 9936 103848 9988
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 106658 9766 106710 9818
rect 106722 9766 106774 9818
rect 106786 9766 106838 9818
rect 106850 9766 106902 9818
rect 106914 9766 106966 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 105922 9222 105974 9274
rect 105986 9222 106038 9274
rect 106050 9222 106102 9274
rect 106114 9222 106166 9274
rect 106178 9222 106230 9274
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 106658 8678 106710 8730
rect 106722 8678 106774 8730
rect 106786 8678 106838 8730
rect 106850 8678 106902 8730
rect 106914 8678 106966 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 105922 8134 105974 8186
rect 105986 8134 106038 8186
rect 106050 8134 106102 8186
rect 106114 8134 106166 8186
rect 106178 8134 106230 8186
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 66314 7590 66366 7642
rect 66378 7590 66430 7642
rect 66442 7590 66494 7642
rect 66506 7590 66558 7642
rect 66570 7590 66622 7642
rect 97034 7590 97086 7642
rect 97098 7590 97150 7642
rect 97162 7590 97214 7642
rect 97226 7590 97278 7642
rect 97290 7590 97342 7642
rect 106658 7590 106710 7642
rect 106722 7590 106774 7642
rect 106786 7590 106838 7642
rect 106850 7590 106902 7642
rect 106914 7590 106966 7642
rect 16120 7531 16172 7540
rect 16120 7497 16129 7531
rect 16129 7497 16163 7531
rect 16163 7497 16172 7531
rect 16120 7488 16172 7497
rect 90640 7531 90692 7540
rect 90640 7497 90649 7531
rect 90649 7497 90683 7531
rect 90683 7497 90692 7531
rect 90640 7488 90692 7497
rect 90732 7531 90784 7540
rect 90732 7497 90741 7531
rect 90741 7497 90775 7531
rect 90775 7497 90784 7531
rect 90732 7488 90784 7497
rect 91008 7531 91060 7540
rect 91008 7497 91017 7531
rect 91017 7497 91051 7531
rect 91051 7497 91060 7531
rect 91008 7488 91060 7497
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 96374 7046 96426 7098
rect 96438 7046 96490 7098
rect 96502 7046 96554 7098
rect 96566 7046 96618 7098
rect 96630 7046 96682 7098
rect 105922 7046 105974 7098
rect 105986 7046 106038 7098
rect 106050 7046 106102 7098
rect 106114 7046 106166 7098
rect 106178 7046 106230 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 66314 6502 66366 6554
rect 66378 6502 66430 6554
rect 66442 6502 66494 6554
rect 66506 6502 66558 6554
rect 66570 6502 66622 6554
rect 97034 6502 97086 6554
rect 97098 6502 97150 6554
rect 97162 6502 97214 6554
rect 97226 6502 97278 6554
rect 97290 6502 97342 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 96374 5958 96426 6010
rect 96438 5958 96490 6010
rect 96502 5958 96554 6010
rect 96566 5958 96618 6010
rect 96630 5958 96682 6010
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 66314 5414 66366 5466
rect 66378 5414 66430 5466
rect 66442 5414 66494 5466
rect 66506 5414 66558 5466
rect 66570 5414 66622 5466
rect 97034 5414 97086 5466
rect 97098 5414 97150 5466
rect 97162 5414 97214 5466
rect 97226 5414 97278 5466
rect 97290 5414 97342 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 96374 4870 96426 4922
rect 96438 4870 96490 4922
rect 96502 4870 96554 4922
rect 96566 4870 96618 4922
rect 96630 4870 96682 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 66314 4326 66366 4378
rect 66378 4326 66430 4378
rect 66442 4326 66494 4378
rect 66506 4326 66558 4378
rect 66570 4326 66622 4378
rect 97034 4326 97086 4378
rect 97098 4326 97150 4378
rect 97162 4326 97214 4378
rect 97226 4326 97278 4378
rect 97290 4326 97342 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 96374 3782 96426 3834
rect 96438 3782 96490 3834
rect 96502 3782 96554 3834
rect 96566 3782 96618 3834
rect 96630 3782 96682 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 66314 3238 66366 3290
rect 66378 3238 66430 3290
rect 66442 3238 66494 3290
rect 66506 3238 66558 3290
rect 66570 3238 66622 3290
rect 97034 3238 97086 3290
rect 97098 3238 97150 3290
rect 97162 3238 97214 3290
rect 97226 3238 97278 3290
rect 97290 3238 97342 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 96374 2694 96426 2746
rect 96438 2694 96490 2746
rect 96502 2694 96554 2746
rect 96566 2694 96618 2746
rect 96630 2694 96682 2746
rect 23480 2635 23532 2644
rect 23480 2601 23489 2635
rect 23489 2601 23523 2635
rect 23523 2601 23532 2635
rect 23480 2592 23532 2601
rect 24768 2635 24820 2644
rect 24768 2601 24777 2635
rect 24777 2601 24811 2635
rect 24811 2601 24820 2635
rect 24768 2592 24820 2601
rect 25872 2635 25924 2644
rect 25872 2601 25881 2635
rect 25881 2601 25915 2635
rect 25915 2601 25924 2635
rect 25872 2592 25924 2601
rect 27160 2635 27212 2644
rect 27160 2601 27169 2635
rect 27169 2601 27203 2635
rect 27203 2601 27212 2635
rect 27160 2592 27212 2601
rect 28448 2635 28500 2644
rect 28448 2601 28457 2635
rect 28457 2601 28491 2635
rect 28491 2601 28500 2635
rect 28448 2592 28500 2601
rect 29276 2635 29328 2644
rect 29276 2601 29285 2635
rect 29285 2601 29319 2635
rect 29319 2601 29328 2635
rect 29276 2592 29328 2601
rect 30564 2635 30616 2644
rect 30564 2601 30573 2635
rect 30573 2601 30607 2635
rect 30607 2601 30616 2635
rect 30564 2592 30616 2601
rect 31668 2635 31720 2644
rect 31668 2601 31677 2635
rect 31677 2601 31711 2635
rect 31711 2601 31720 2635
rect 31668 2592 31720 2601
rect 32956 2635 33008 2644
rect 32956 2601 32965 2635
rect 32965 2601 32999 2635
rect 32999 2601 33008 2635
rect 32956 2592 33008 2601
rect 34244 2635 34296 2644
rect 34244 2601 34253 2635
rect 34253 2601 34287 2635
rect 34287 2601 34296 2635
rect 34244 2592 34296 2601
rect 35440 2592 35492 2644
rect 36360 2635 36412 2644
rect 36360 2601 36369 2635
rect 36369 2601 36403 2635
rect 36403 2601 36412 2635
rect 36360 2592 36412 2601
rect 37464 2635 37516 2644
rect 37464 2601 37473 2635
rect 37473 2601 37507 2635
rect 37507 2601 37516 2635
rect 37464 2592 37516 2601
rect 38752 2635 38804 2644
rect 38752 2601 38761 2635
rect 38761 2601 38795 2635
rect 38795 2601 38804 2635
rect 38752 2592 38804 2601
rect 39948 2592 40000 2644
rect 41328 2635 41380 2644
rect 41328 2601 41337 2635
rect 41337 2601 41371 2635
rect 41371 2601 41380 2635
rect 41328 2592 41380 2601
rect 42156 2635 42208 2644
rect 42156 2601 42165 2635
rect 42165 2601 42199 2635
rect 42199 2601 42208 2635
rect 42156 2592 42208 2601
rect 43444 2635 43496 2644
rect 43444 2601 43453 2635
rect 43453 2601 43487 2635
rect 43487 2601 43496 2635
rect 43444 2592 43496 2601
rect 23204 2295 23256 2304
rect 23204 2261 23213 2295
rect 23213 2261 23247 2295
rect 23247 2261 23256 2295
rect 23204 2252 23256 2261
rect 24492 2295 24544 2304
rect 24492 2261 24501 2295
rect 24501 2261 24535 2295
rect 24535 2261 24544 2295
rect 24492 2252 24544 2261
rect 25780 2295 25832 2304
rect 25780 2261 25789 2295
rect 25789 2261 25823 2295
rect 25823 2261 25832 2295
rect 25780 2252 25832 2261
rect 27068 2295 27120 2304
rect 27068 2261 27077 2295
rect 27077 2261 27111 2295
rect 27111 2261 27120 2295
rect 27068 2252 27120 2261
rect 28356 2295 28408 2304
rect 28356 2261 28365 2295
rect 28365 2261 28399 2295
rect 28399 2261 28408 2295
rect 28356 2252 28408 2261
rect 29000 2295 29052 2304
rect 29000 2261 29009 2295
rect 29009 2261 29043 2295
rect 29043 2261 29052 2295
rect 29000 2252 29052 2261
rect 30288 2295 30340 2304
rect 30288 2261 30297 2295
rect 30297 2261 30331 2295
rect 30331 2261 30340 2295
rect 30288 2252 30340 2261
rect 31576 2295 31628 2304
rect 31576 2261 31585 2295
rect 31585 2261 31619 2295
rect 31619 2261 31628 2295
rect 31576 2252 31628 2261
rect 32864 2295 32916 2304
rect 32864 2261 32873 2295
rect 32873 2261 32907 2295
rect 32907 2261 32916 2295
rect 32864 2252 32916 2261
rect 34152 2295 34204 2304
rect 34152 2261 34161 2295
rect 34161 2261 34195 2295
rect 34195 2261 34204 2295
rect 34152 2252 34204 2261
rect 35440 2295 35492 2304
rect 35440 2261 35449 2295
rect 35449 2261 35483 2295
rect 35483 2261 35492 2295
rect 35440 2252 35492 2261
rect 36084 2295 36136 2304
rect 36084 2261 36093 2295
rect 36093 2261 36127 2295
rect 36127 2261 36136 2295
rect 36084 2252 36136 2261
rect 37372 2295 37424 2304
rect 37372 2261 37381 2295
rect 37381 2261 37415 2295
rect 37415 2261 37424 2295
rect 37372 2252 37424 2261
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 39948 2295 40000 2304
rect 39948 2261 39957 2295
rect 39957 2261 39991 2295
rect 39991 2261 40000 2295
rect 39948 2252 40000 2261
rect 41236 2295 41288 2304
rect 41236 2261 41245 2295
rect 41245 2261 41279 2295
rect 41279 2261 41288 2295
rect 41236 2252 41288 2261
rect 41880 2295 41932 2304
rect 41880 2261 41889 2295
rect 41889 2261 41923 2295
rect 41923 2261 41932 2295
rect 41880 2252 41932 2261
rect 43168 2295 43220 2304
rect 43168 2261 43177 2295
rect 43177 2261 43211 2295
rect 43211 2261 43220 2295
rect 43168 2252 43220 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 66314 2150 66366 2202
rect 66378 2150 66430 2202
rect 66442 2150 66494 2202
rect 66506 2150 66558 2202
rect 66570 2150 66622 2202
rect 97034 2150 97086 2202
rect 97098 2150 97150 2202
rect 97162 2150 97214 2202
rect 97226 2150 97278 2202
rect 97290 2150 97342 2202
<< metal2 >>
rect 98550 129200 98606 130000
rect 98564 128382 98592 129200
rect 98552 128376 98604 128382
rect 98552 128318 98604 128324
rect 102140 128376 102192 128382
rect 102140 128318 102192 128324
rect 4874 127324 5182 127333
rect 4874 127322 4880 127324
rect 4936 127322 4960 127324
rect 5016 127322 5040 127324
rect 5096 127322 5120 127324
rect 5176 127322 5182 127324
rect 4936 127270 4938 127322
rect 5118 127270 5120 127322
rect 4874 127268 4880 127270
rect 4936 127268 4960 127270
rect 5016 127268 5040 127270
rect 5096 127268 5120 127270
rect 5176 127268 5182 127270
rect 4874 127259 5182 127268
rect 35594 127324 35902 127333
rect 35594 127322 35600 127324
rect 35656 127322 35680 127324
rect 35736 127322 35760 127324
rect 35816 127322 35840 127324
rect 35896 127322 35902 127324
rect 35656 127270 35658 127322
rect 35838 127270 35840 127322
rect 35594 127268 35600 127270
rect 35656 127268 35680 127270
rect 35736 127268 35760 127270
rect 35816 127268 35840 127270
rect 35896 127268 35902 127270
rect 35594 127259 35902 127268
rect 66314 127324 66622 127333
rect 66314 127322 66320 127324
rect 66376 127322 66400 127324
rect 66456 127322 66480 127324
rect 66536 127322 66560 127324
rect 66616 127322 66622 127324
rect 66376 127270 66378 127322
rect 66558 127270 66560 127322
rect 66314 127268 66320 127270
rect 66376 127268 66400 127270
rect 66456 127268 66480 127270
rect 66536 127268 66560 127270
rect 66616 127268 66622 127270
rect 66314 127259 66622 127268
rect 97034 127324 97342 127333
rect 97034 127322 97040 127324
rect 97096 127322 97120 127324
rect 97176 127322 97200 127324
rect 97256 127322 97280 127324
rect 97336 127322 97342 127324
rect 97096 127270 97098 127322
rect 97278 127270 97280 127322
rect 97034 127268 97040 127270
rect 97096 127268 97120 127270
rect 97176 127268 97200 127270
rect 97256 127268 97280 127270
rect 97336 127268 97342 127270
rect 97034 127259 97342 127268
rect 4214 126780 4522 126789
rect 4214 126778 4220 126780
rect 4276 126778 4300 126780
rect 4356 126778 4380 126780
rect 4436 126778 4460 126780
rect 4516 126778 4522 126780
rect 4276 126726 4278 126778
rect 4458 126726 4460 126778
rect 4214 126724 4220 126726
rect 4276 126724 4300 126726
rect 4356 126724 4380 126726
rect 4436 126724 4460 126726
rect 4516 126724 4522 126726
rect 4214 126715 4522 126724
rect 34934 126780 35242 126789
rect 34934 126778 34940 126780
rect 34996 126778 35020 126780
rect 35076 126778 35100 126780
rect 35156 126778 35180 126780
rect 35236 126778 35242 126780
rect 34996 126726 34998 126778
rect 35178 126726 35180 126778
rect 34934 126724 34940 126726
rect 34996 126724 35020 126726
rect 35076 126724 35100 126726
rect 35156 126724 35180 126726
rect 35236 126724 35242 126726
rect 34934 126715 35242 126724
rect 65654 126780 65962 126789
rect 65654 126778 65660 126780
rect 65716 126778 65740 126780
rect 65796 126778 65820 126780
rect 65876 126778 65900 126780
rect 65956 126778 65962 126780
rect 65716 126726 65718 126778
rect 65898 126726 65900 126778
rect 65654 126724 65660 126726
rect 65716 126724 65740 126726
rect 65796 126724 65820 126726
rect 65876 126724 65900 126726
rect 65956 126724 65962 126726
rect 65654 126715 65962 126724
rect 96374 126780 96682 126789
rect 96374 126778 96380 126780
rect 96436 126778 96460 126780
rect 96516 126778 96540 126780
rect 96596 126778 96620 126780
rect 96676 126778 96682 126780
rect 96436 126726 96438 126778
rect 96618 126726 96620 126778
rect 96374 126724 96380 126726
rect 96436 126724 96460 126726
rect 96516 126724 96540 126726
rect 96596 126724 96620 126726
rect 96676 126724 96682 126726
rect 96374 126715 96682 126724
rect 42340 126472 42392 126478
rect 42340 126414 42392 126420
rect 77298 126440 77354 126449
rect 36084 126404 36136 126410
rect 36084 126346 36136 126352
rect 36268 126404 36320 126410
rect 36268 126346 36320 126352
rect 37740 126404 37792 126410
rect 37740 126346 37792 126352
rect 41328 126404 41380 126410
rect 41328 126346 41380 126352
rect 4874 126236 5182 126245
rect 4874 126234 4880 126236
rect 4936 126234 4960 126236
rect 5016 126234 5040 126236
rect 5096 126234 5120 126236
rect 5176 126234 5182 126236
rect 4936 126182 4938 126234
rect 5118 126182 5120 126234
rect 4874 126180 4880 126182
rect 4936 126180 4960 126182
rect 5016 126180 5040 126182
rect 5096 126180 5120 126182
rect 5176 126180 5182 126182
rect 4874 126171 5182 126180
rect 35594 126236 35902 126245
rect 35594 126234 35600 126236
rect 35656 126234 35680 126236
rect 35736 126234 35760 126236
rect 35816 126234 35840 126236
rect 35896 126234 35902 126236
rect 35656 126182 35658 126234
rect 35838 126182 35840 126234
rect 35594 126180 35600 126182
rect 35656 126180 35680 126182
rect 35736 126180 35760 126182
rect 35816 126180 35840 126182
rect 35896 126180 35902 126182
rect 35594 126171 35902 126180
rect 9588 126132 9640 126138
rect 9588 126074 9640 126080
rect 8208 126064 8260 126070
rect 8208 126006 8260 126012
rect 8116 125996 8168 126002
rect 8116 125938 8168 125944
rect 7932 125928 7984 125934
rect 7932 125870 7984 125876
rect 7840 125860 7892 125866
rect 7840 125802 7892 125808
rect 4214 125692 4522 125701
rect 4214 125690 4220 125692
rect 4276 125690 4300 125692
rect 4356 125690 4380 125692
rect 4436 125690 4460 125692
rect 4516 125690 4522 125692
rect 4276 125638 4278 125690
rect 4458 125638 4460 125690
rect 4214 125636 4220 125638
rect 4276 125636 4300 125638
rect 4356 125636 4380 125638
rect 4436 125636 4460 125638
rect 4516 125636 4522 125638
rect 4214 125627 4522 125636
rect 4874 125148 5182 125157
rect 4874 125146 4880 125148
rect 4936 125146 4960 125148
rect 5016 125146 5040 125148
rect 5096 125146 5120 125148
rect 5176 125146 5182 125148
rect 4936 125094 4938 125146
rect 5118 125094 5120 125146
rect 4874 125092 4880 125094
rect 4936 125092 4960 125094
rect 5016 125092 5040 125094
rect 5096 125092 5120 125094
rect 5176 125092 5182 125094
rect 4874 125083 5182 125092
rect 4214 124604 4522 124613
rect 4214 124602 4220 124604
rect 4276 124602 4300 124604
rect 4356 124602 4380 124604
rect 4436 124602 4460 124604
rect 4516 124602 4522 124604
rect 4276 124550 4278 124602
rect 4458 124550 4460 124602
rect 4214 124548 4220 124550
rect 4276 124548 4300 124550
rect 4356 124548 4380 124550
rect 4436 124548 4460 124550
rect 4516 124548 4522 124550
rect 4214 124539 4522 124548
rect 4874 124060 5182 124069
rect 4874 124058 4880 124060
rect 4936 124058 4960 124060
rect 5016 124058 5040 124060
rect 5096 124058 5120 124060
rect 5176 124058 5182 124060
rect 4936 124006 4938 124058
rect 5118 124006 5120 124058
rect 4874 124004 4880 124006
rect 4936 124004 4960 124006
rect 5016 124004 5040 124006
rect 5096 124004 5120 124006
rect 5176 124004 5182 124006
rect 4874 123995 5182 124004
rect 4214 123516 4522 123525
rect 4214 123514 4220 123516
rect 4276 123514 4300 123516
rect 4356 123514 4380 123516
rect 4436 123514 4460 123516
rect 4516 123514 4522 123516
rect 4276 123462 4278 123514
rect 4458 123462 4460 123514
rect 4214 123460 4220 123462
rect 4276 123460 4300 123462
rect 4356 123460 4380 123462
rect 4436 123460 4460 123462
rect 4516 123460 4522 123462
rect 4214 123451 4522 123460
rect 4874 122972 5182 122981
rect 4874 122970 4880 122972
rect 4936 122970 4960 122972
rect 5016 122970 5040 122972
rect 5096 122970 5120 122972
rect 5176 122970 5182 122972
rect 4936 122918 4938 122970
rect 5118 122918 5120 122970
rect 4874 122916 4880 122918
rect 4936 122916 4960 122918
rect 5016 122916 5040 122918
rect 5096 122916 5120 122918
rect 5176 122916 5182 122918
rect 4874 122907 5182 122916
rect 4214 122428 4522 122437
rect 4214 122426 4220 122428
rect 4276 122426 4300 122428
rect 4356 122426 4380 122428
rect 4436 122426 4460 122428
rect 4516 122426 4522 122428
rect 4276 122374 4278 122426
rect 4458 122374 4460 122426
rect 4214 122372 4220 122374
rect 4276 122372 4300 122374
rect 4356 122372 4380 122374
rect 4436 122372 4460 122374
rect 4516 122372 4522 122374
rect 4214 122363 4522 122372
rect 4874 121884 5182 121893
rect 4874 121882 4880 121884
rect 4936 121882 4960 121884
rect 5016 121882 5040 121884
rect 5096 121882 5120 121884
rect 5176 121882 5182 121884
rect 4936 121830 4938 121882
rect 5118 121830 5120 121882
rect 4874 121828 4880 121830
rect 4936 121828 4960 121830
rect 5016 121828 5040 121830
rect 5096 121828 5120 121830
rect 5176 121828 5182 121830
rect 4874 121819 5182 121828
rect 4214 121340 4522 121349
rect 4214 121338 4220 121340
rect 4276 121338 4300 121340
rect 4356 121338 4380 121340
rect 4436 121338 4460 121340
rect 4516 121338 4522 121340
rect 4276 121286 4278 121338
rect 4458 121286 4460 121338
rect 4214 121284 4220 121286
rect 4276 121284 4300 121286
rect 4356 121284 4380 121286
rect 4436 121284 4460 121286
rect 4516 121284 4522 121286
rect 4214 121275 4522 121284
rect 4874 120796 5182 120805
rect 4874 120794 4880 120796
rect 4936 120794 4960 120796
rect 5016 120794 5040 120796
rect 5096 120794 5120 120796
rect 5176 120794 5182 120796
rect 4936 120742 4938 120794
rect 5118 120742 5120 120794
rect 4874 120740 4880 120742
rect 4936 120740 4960 120742
rect 5016 120740 5040 120742
rect 5096 120740 5120 120742
rect 5176 120740 5182 120742
rect 4874 120731 5182 120740
rect 4214 120252 4522 120261
rect 4214 120250 4220 120252
rect 4276 120250 4300 120252
rect 4356 120250 4380 120252
rect 4436 120250 4460 120252
rect 4516 120250 4522 120252
rect 4276 120198 4278 120250
rect 4458 120198 4460 120250
rect 4214 120196 4220 120198
rect 4276 120196 4300 120198
rect 4356 120196 4380 120198
rect 4436 120196 4460 120198
rect 4516 120196 4522 120198
rect 4214 120187 4522 120196
rect 4874 119708 5182 119717
rect 4874 119706 4880 119708
rect 4936 119706 4960 119708
rect 5016 119706 5040 119708
rect 5096 119706 5120 119708
rect 5176 119706 5182 119708
rect 4936 119654 4938 119706
rect 5118 119654 5120 119706
rect 4874 119652 4880 119654
rect 4936 119652 4960 119654
rect 5016 119652 5040 119654
rect 5096 119652 5120 119654
rect 5176 119652 5182 119654
rect 4874 119643 5182 119652
rect 4214 119164 4522 119173
rect 4214 119162 4220 119164
rect 4276 119162 4300 119164
rect 4356 119162 4380 119164
rect 4436 119162 4460 119164
rect 4516 119162 4522 119164
rect 4276 119110 4278 119162
rect 4458 119110 4460 119162
rect 4214 119108 4220 119110
rect 4276 119108 4300 119110
rect 4356 119108 4380 119110
rect 4436 119108 4460 119110
rect 4516 119108 4522 119110
rect 4214 119099 4522 119108
rect 4874 118620 5182 118629
rect 4874 118618 4880 118620
rect 4936 118618 4960 118620
rect 5016 118618 5040 118620
rect 5096 118618 5120 118620
rect 5176 118618 5182 118620
rect 4936 118566 4938 118618
rect 5118 118566 5120 118618
rect 4874 118564 4880 118566
rect 4936 118564 4960 118566
rect 5016 118564 5040 118566
rect 5096 118564 5120 118566
rect 5176 118564 5182 118566
rect 4874 118555 5182 118564
rect 4214 118076 4522 118085
rect 4214 118074 4220 118076
rect 4276 118074 4300 118076
rect 4356 118074 4380 118076
rect 4436 118074 4460 118076
rect 4516 118074 4522 118076
rect 4276 118022 4278 118074
rect 4458 118022 4460 118074
rect 4214 118020 4220 118022
rect 4276 118020 4300 118022
rect 4356 118020 4380 118022
rect 4436 118020 4460 118022
rect 4516 118020 4522 118022
rect 4214 118011 4522 118020
rect 4874 117532 5182 117541
rect 4874 117530 4880 117532
rect 4936 117530 4960 117532
rect 5016 117530 5040 117532
rect 5096 117530 5120 117532
rect 5176 117530 5182 117532
rect 4936 117478 4938 117530
rect 5118 117478 5120 117530
rect 4874 117476 4880 117478
rect 4936 117476 4960 117478
rect 5016 117476 5040 117478
rect 5096 117476 5120 117478
rect 5176 117476 5182 117478
rect 4874 117467 5182 117476
rect 4214 116988 4522 116997
rect 4214 116986 4220 116988
rect 4276 116986 4300 116988
rect 4356 116986 4380 116988
rect 4436 116986 4460 116988
rect 4516 116986 4522 116988
rect 4276 116934 4278 116986
rect 4458 116934 4460 116986
rect 4214 116932 4220 116934
rect 4276 116932 4300 116934
rect 4356 116932 4380 116934
rect 4436 116932 4460 116934
rect 4516 116932 4522 116934
rect 4214 116923 4522 116932
rect 4874 116444 5182 116453
rect 4874 116442 4880 116444
rect 4936 116442 4960 116444
rect 5016 116442 5040 116444
rect 5096 116442 5120 116444
rect 5176 116442 5182 116444
rect 4936 116390 4938 116442
rect 5118 116390 5120 116442
rect 4874 116388 4880 116390
rect 4936 116388 4960 116390
rect 5016 116388 5040 116390
rect 5096 116388 5120 116390
rect 5176 116388 5182 116390
rect 4874 116379 5182 116388
rect 4214 115900 4522 115909
rect 4214 115898 4220 115900
rect 4276 115898 4300 115900
rect 4356 115898 4380 115900
rect 4436 115898 4460 115900
rect 4516 115898 4522 115900
rect 4276 115846 4278 115898
rect 4458 115846 4460 115898
rect 4214 115844 4220 115846
rect 4276 115844 4300 115846
rect 4356 115844 4380 115846
rect 4436 115844 4460 115846
rect 4516 115844 4522 115846
rect 4214 115835 4522 115844
rect 4874 115356 5182 115365
rect 4874 115354 4880 115356
rect 4936 115354 4960 115356
rect 5016 115354 5040 115356
rect 5096 115354 5120 115356
rect 5176 115354 5182 115356
rect 4936 115302 4938 115354
rect 5118 115302 5120 115354
rect 4874 115300 4880 115302
rect 4936 115300 4960 115302
rect 5016 115300 5040 115302
rect 5096 115300 5120 115302
rect 5176 115300 5182 115302
rect 4874 115291 5182 115300
rect 4214 114812 4522 114821
rect 4214 114810 4220 114812
rect 4276 114810 4300 114812
rect 4356 114810 4380 114812
rect 4436 114810 4460 114812
rect 4516 114810 4522 114812
rect 4276 114758 4278 114810
rect 4458 114758 4460 114810
rect 4214 114756 4220 114758
rect 4276 114756 4300 114758
rect 4356 114756 4380 114758
rect 4436 114756 4460 114758
rect 4516 114756 4522 114758
rect 4214 114747 4522 114756
rect 4874 114268 5182 114277
rect 4874 114266 4880 114268
rect 4936 114266 4960 114268
rect 5016 114266 5040 114268
rect 5096 114266 5120 114268
rect 5176 114266 5182 114268
rect 4936 114214 4938 114266
rect 5118 114214 5120 114266
rect 4874 114212 4880 114214
rect 4936 114212 4960 114214
rect 5016 114212 5040 114214
rect 5096 114212 5120 114214
rect 5176 114212 5182 114214
rect 4874 114203 5182 114212
rect 4214 113724 4522 113733
rect 4214 113722 4220 113724
rect 4276 113722 4300 113724
rect 4356 113722 4380 113724
rect 4436 113722 4460 113724
rect 4516 113722 4522 113724
rect 4276 113670 4278 113722
rect 4458 113670 4460 113722
rect 4214 113668 4220 113670
rect 4276 113668 4300 113670
rect 4356 113668 4380 113670
rect 4436 113668 4460 113670
rect 4516 113668 4522 113670
rect 4214 113659 4522 113668
rect 4874 113180 5182 113189
rect 4874 113178 4880 113180
rect 4936 113178 4960 113180
rect 5016 113178 5040 113180
rect 5096 113178 5120 113180
rect 5176 113178 5182 113180
rect 4936 113126 4938 113178
rect 5118 113126 5120 113178
rect 4874 113124 4880 113126
rect 4936 113124 4960 113126
rect 5016 113124 5040 113126
rect 5096 113124 5120 113126
rect 5176 113124 5182 113126
rect 4874 113115 5182 113124
rect 4214 112636 4522 112645
rect 4214 112634 4220 112636
rect 4276 112634 4300 112636
rect 4356 112634 4380 112636
rect 4436 112634 4460 112636
rect 4516 112634 4522 112636
rect 4276 112582 4278 112634
rect 4458 112582 4460 112634
rect 4214 112580 4220 112582
rect 4276 112580 4300 112582
rect 4356 112580 4380 112582
rect 4436 112580 4460 112582
rect 4516 112580 4522 112582
rect 4214 112571 4522 112580
rect 4874 112092 5182 112101
rect 4874 112090 4880 112092
rect 4936 112090 4960 112092
rect 5016 112090 5040 112092
rect 5096 112090 5120 112092
rect 5176 112090 5182 112092
rect 4936 112038 4938 112090
rect 5118 112038 5120 112090
rect 4874 112036 4880 112038
rect 4936 112036 4960 112038
rect 5016 112036 5040 112038
rect 5096 112036 5120 112038
rect 5176 112036 5182 112038
rect 4874 112027 5182 112036
rect 4214 111548 4522 111557
rect 4214 111546 4220 111548
rect 4276 111546 4300 111548
rect 4356 111546 4380 111548
rect 4436 111546 4460 111548
rect 4516 111546 4522 111548
rect 4276 111494 4278 111546
rect 4458 111494 4460 111546
rect 4214 111492 4220 111494
rect 4276 111492 4300 111494
rect 4356 111492 4380 111494
rect 4436 111492 4460 111494
rect 4516 111492 4522 111494
rect 4214 111483 4522 111492
rect 4874 111004 5182 111013
rect 4874 111002 4880 111004
rect 4936 111002 4960 111004
rect 5016 111002 5040 111004
rect 5096 111002 5120 111004
rect 5176 111002 5182 111004
rect 4936 110950 4938 111002
rect 5118 110950 5120 111002
rect 4874 110948 4880 110950
rect 4936 110948 4960 110950
rect 5016 110948 5040 110950
rect 5096 110948 5120 110950
rect 5176 110948 5182 110950
rect 4874 110939 5182 110948
rect 4214 110460 4522 110469
rect 4214 110458 4220 110460
rect 4276 110458 4300 110460
rect 4356 110458 4380 110460
rect 4436 110458 4460 110460
rect 4516 110458 4522 110460
rect 4276 110406 4278 110458
rect 4458 110406 4460 110458
rect 4214 110404 4220 110406
rect 4276 110404 4300 110406
rect 4356 110404 4380 110406
rect 4436 110404 4460 110406
rect 4516 110404 4522 110406
rect 4214 110395 4522 110404
rect 4874 109916 5182 109925
rect 4874 109914 4880 109916
rect 4936 109914 4960 109916
rect 5016 109914 5040 109916
rect 5096 109914 5120 109916
rect 5176 109914 5182 109916
rect 4936 109862 4938 109914
rect 5118 109862 5120 109914
rect 4874 109860 4880 109862
rect 4936 109860 4960 109862
rect 5016 109860 5040 109862
rect 5096 109860 5120 109862
rect 5176 109860 5182 109862
rect 4874 109851 5182 109860
rect 4214 109372 4522 109381
rect 4214 109370 4220 109372
rect 4276 109370 4300 109372
rect 4356 109370 4380 109372
rect 4436 109370 4460 109372
rect 4516 109370 4522 109372
rect 4276 109318 4278 109370
rect 4458 109318 4460 109370
rect 4214 109316 4220 109318
rect 4276 109316 4300 109318
rect 4356 109316 4380 109318
rect 4436 109316 4460 109318
rect 4516 109316 4522 109318
rect 4214 109307 4522 109316
rect 4874 108828 5182 108837
rect 4874 108826 4880 108828
rect 4936 108826 4960 108828
rect 5016 108826 5040 108828
rect 5096 108826 5120 108828
rect 5176 108826 5182 108828
rect 4936 108774 4938 108826
rect 5118 108774 5120 108826
rect 4874 108772 4880 108774
rect 4936 108772 4960 108774
rect 5016 108772 5040 108774
rect 5096 108772 5120 108774
rect 5176 108772 5182 108774
rect 4874 108763 5182 108772
rect 4214 108284 4522 108293
rect 4214 108282 4220 108284
rect 4276 108282 4300 108284
rect 4356 108282 4380 108284
rect 4436 108282 4460 108284
rect 4516 108282 4522 108284
rect 4276 108230 4278 108282
rect 4458 108230 4460 108282
rect 4214 108228 4220 108230
rect 4276 108228 4300 108230
rect 4356 108228 4380 108230
rect 4436 108228 4460 108230
rect 4516 108228 4522 108230
rect 4214 108219 4522 108228
rect 4874 107740 5182 107749
rect 4874 107738 4880 107740
rect 4936 107738 4960 107740
rect 5016 107738 5040 107740
rect 5096 107738 5120 107740
rect 5176 107738 5182 107740
rect 4936 107686 4938 107738
rect 5118 107686 5120 107738
rect 4874 107684 4880 107686
rect 4936 107684 4960 107686
rect 5016 107684 5040 107686
rect 5096 107684 5120 107686
rect 5176 107684 5182 107686
rect 4874 107675 5182 107684
rect 4214 107196 4522 107205
rect 4214 107194 4220 107196
rect 4276 107194 4300 107196
rect 4356 107194 4380 107196
rect 4436 107194 4460 107196
rect 4516 107194 4522 107196
rect 4276 107142 4278 107194
rect 4458 107142 4460 107194
rect 4214 107140 4220 107142
rect 4276 107140 4300 107142
rect 4356 107140 4380 107142
rect 4436 107140 4460 107142
rect 4516 107140 4522 107142
rect 4214 107131 4522 107140
rect 4874 106652 5182 106661
rect 4874 106650 4880 106652
rect 4936 106650 4960 106652
rect 5016 106650 5040 106652
rect 5096 106650 5120 106652
rect 5176 106650 5182 106652
rect 4936 106598 4938 106650
rect 5118 106598 5120 106650
rect 4874 106596 4880 106598
rect 4936 106596 4960 106598
rect 5016 106596 5040 106598
rect 5096 106596 5120 106598
rect 5176 106596 5182 106598
rect 4874 106587 5182 106596
rect 4214 106108 4522 106117
rect 4214 106106 4220 106108
rect 4276 106106 4300 106108
rect 4356 106106 4380 106108
rect 4436 106106 4460 106108
rect 4516 106106 4522 106108
rect 4276 106054 4278 106106
rect 4458 106054 4460 106106
rect 4214 106052 4220 106054
rect 4276 106052 4300 106054
rect 4356 106052 4380 106054
rect 4436 106052 4460 106054
rect 4516 106052 4522 106054
rect 4214 106043 4522 106052
rect 4874 105564 5182 105573
rect 4874 105562 4880 105564
rect 4936 105562 4960 105564
rect 5016 105562 5040 105564
rect 5096 105562 5120 105564
rect 5176 105562 5182 105564
rect 4936 105510 4938 105562
rect 5118 105510 5120 105562
rect 4874 105508 4880 105510
rect 4936 105508 4960 105510
rect 5016 105508 5040 105510
rect 5096 105508 5120 105510
rect 5176 105508 5182 105510
rect 4874 105499 5182 105508
rect 4214 105020 4522 105029
rect 4214 105018 4220 105020
rect 4276 105018 4300 105020
rect 4356 105018 4380 105020
rect 4436 105018 4460 105020
rect 4516 105018 4522 105020
rect 4276 104966 4278 105018
rect 4458 104966 4460 105018
rect 4214 104964 4220 104966
rect 4276 104964 4300 104966
rect 4356 104964 4380 104966
rect 4436 104964 4460 104966
rect 4516 104964 4522 104966
rect 4214 104955 4522 104964
rect 4874 104476 5182 104485
rect 4874 104474 4880 104476
rect 4936 104474 4960 104476
rect 5016 104474 5040 104476
rect 5096 104474 5120 104476
rect 5176 104474 5182 104476
rect 4936 104422 4938 104474
rect 5118 104422 5120 104474
rect 4874 104420 4880 104422
rect 4936 104420 4960 104422
rect 5016 104420 5040 104422
rect 5096 104420 5120 104422
rect 5176 104420 5182 104422
rect 4874 104411 5182 104420
rect 4214 103932 4522 103941
rect 4214 103930 4220 103932
rect 4276 103930 4300 103932
rect 4356 103930 4380 103932
rect 4436 103930 4460 103932
rect 4516 103930 4522 103932
rect 4276 103878 4278 103930
rect 4458 103878 4460 103930
rect 4214 103876 4220 103878
rect 4276 103876 4300 103878
rect 4356 103876 4380 103878
rect 4436 103876 4460 103878
rect 4516 103876 4522 103878
rect 4214 103867 4522 103876
rect 4874 103388 5182 103397
rect 4874 103386 4880 103388
rect 4936 103386 4960 103388
rect 5016 103386 5040 103388
rect 5096 103386 5120 103388
rect 5176 103386 5182 103388
rect 4936 103334 4938 103386
rect 5118 103334 5120 103386
rect 4874 103332 4880 103334
rect 4936 103332 4960 103334
rect 5016 103332 5040 103334
rect 5096 103332 5120 103334
rect 5176 103332 5182 103334
rect 4874 103323 5182 103332
rect 4214 102844 4522 102853
rect 4214 102842 4220 102844
rect 4276 102842 4300 102844
rect 4356 102842 4380 102844
rect 4436 102842 4460 102844
rect 4516 102842 4522 102844
rect 4276 102790 4278 102842
rect 4458 102790 4460 102842
rect 4214 102788 4220 102790
rect 4276 102788 4300 102790
rect 4356 102788 4380 102790
rect 4436 102788 4460 102790
rect 4516 102788 4522 102790
rect 4214 102779 4522 102788
rect 4874 102300 5182 102309
rect 4874 102298 4880 102300
rect 4936 102298 4960 102300
rect 5016 102298 5040 102300
rect 5096 102298 5120 102300
rect 5176 102298 5182 102300
rect 4936 102246 4938 102298
rect 5118 102246 5120 102298
rect 4874 102244 4880 102246
rect 4936 102244 4960 102246
rect 5016 102244 5040 102246
rect 5096 102244 5120 102246
rect 5176 102244 5182 102246
rect 4874 102235 5182 102244
rect 4214 101756 4522 101765
rect 4214 101754 4220 101756
rect 4276 101754 4300 101756
rect 4356 101754 4380 101756
rect 4436 101754 4460 101756
rect 4516 101754 4522 101756
rect 4276 101702 4278 101754
rect 4458 101702 4460 101754
rect 4214 101700 4220 101702
rect 4276 101700 4300 101702
rect 4356 101700 4380 101702
rect 4436 101700 4460 101702
rect 4516 101700 4522 101702
rect 4214 101691 4522 101700
rect 1216 101448 1268 101454
rect 1214 101416 1216 101425
rect 1268 101416 1270 101425
rect 1214 101351 1270 101360
rect 4874 101212 5182 101221
rect 4874 101210 4880 101212
rect 4936 101210 4960 101212
rect 5016 101210 5040 101212
rect 5096 101210 5120 101212
rect 5176 101210 5182 101212
rect 4936 101158 4938 101210
rect 5118 101158 5120 101210
rect 4874 101156 4880 101158
rect 4936 101156 4960 101158
rect 5016 101156 5040 101158
rect 5096 101156 5120 101158
rect 5176 101156 5182 101158
rect 4874 101147 5182 101156
rect 4214 100668 4522 100677
rect 4214 100666 4220 100668
rect 4276 100666 4300 100668
rect 4356 100666 4380 100668
rect 4436 100666 4460 100668
rect 4516 100666 4522 100668
rect 4276 100614 4278 100666
rect 4458 100614 4460 100666
rect 4214 100612 4220 100614
rect 4276 100612 4300 100614
rect 4356 100612 4380 100614
rect 4436 100612 4460 100614
rect 4516 100612 4522 100614
rect 4214 100603 4522 100612
rect 4874 100124 5182 100133
rect 4874 100122 4880 100124
rect 4936 100122 4960 100124
rect 5016 100122 5040 100124
rect 5096 100122 5120 100124
rect 5176 100122 5182 100124
rect 4936 100070 4938 100122
rect 5118 100070 5120 100122
rect 4874 100068 4880 100070
rect 4936 100068 4960 100070
rect 5016 100068 5040 100070
rect 5096 100068 5120 100070
rect 5176 100068 5182 100070
rect 4874 100059 5182 100068
rect 1400 99884 1452 99890
rect 1400 99826 1452 99832
rect 1412 99385 1440 99826
rect 4214 99580 4522 99589
rect 4214 99578 4220 99580
rect 4276 99578 4300 99580
rect 4356 99578 4380 99580
rect 4436 99578 4460 99580
rect 4516 99578 4522 99580
rect 4276 99526 4278 99578
rect 4458 99526 4460 99578
rect 4214 99524 4220 99526
rect 4276 99524 4300 99526
rect 4356 99524 4380 99526
rect 4436 99524 4460 99526
rect 4516 99524 4522 99526
rect 4214 99515 4522 99524
rect 1398 99376 1454 99385
rect 1398 99311 1454 99320
rect 4874 99036 5182 99045
rect 4874 99034 4880 99036
rect 4936 99034 4960 99036
rect 5016 99034 5040 99036
rect 5096 99034 5120 99036
rect 5176 99034 5182 99036
rect 4936 98982 4938 99034
rect 5118 98982 5120 99034
rect 4874 98980 4880 98982
rect 4936 98980 4960 98982
rect 5016 98980 5040 98982
rect 5096 98980 5120 98982
rect 5176 98980 5182 98982
rect 4874 98971 5182 98980
rect 1308 98796 1360 98802
rect 1308 98738 1360 98744
rect 1320 98705 1348 98738
rect 1306 98696 1362 98705
rect 1306 98631 1362 98640
rect 4214 98492 4522 98501
rect 4214 98490 4220 98492
rect 4276 98490 4300 98492
rect 4356 98490 4380 98492
rect 4436 98490 4460 98492
rect 4516 98490 4522 98492
rect 4276 98438 4278 98490
rect 4458 98438 4460 98490
rect 4214 98436 4220 98438
rect 4276 98436 4300 98438
rect 4356 98436 4380 98438
rect 4436 98436 4460 98438
rect 4516 98436 4522 98438
rect 4214 98427 4522 98436
rect 4874 97948 5182 97957
rect 4874 97946 4880 97948
rect 4936 97946 4960 97948
rect 5016 97946 5040 97948
rect 5096 97946 5120 97948
rect 5176 97946 5182 97948
rect 4936 97894 4938 97946
rect 5118 97894 5120 97946
rect 4874 97892 4880 97894
rect 4936 97892 4960 97894
rect 5016 97892 5040 97894
rect 5096 97892 5120 97894
rect 5176 97892 5182 97894
rect 4874 97883 5182 97892
rect 4214 97404 4522 97413
rect 4214 97402 4220 97404
rect 4276 97402 4300 97404
rect 4356 97402 4380 97404
rect 4436 97402 4460 97404
rect 4516 97402 4522 97404
rect 4276 97350 4278 97402
rect 4458 97350 4460 97402
rect 4214 97348 4220 97350
rect 4276 97348 4300 97350
rect 4356 97348 4380 97350
rect 4436 97348 4460 97350
rect 4516 97348 4522 97350
rect 4214 97339 4522 97348
rect 1308 97096 1360 97102
rect 1308 97038 1360 97044
rect 1320 96665 1348 97038
rect 4874 96860 5182 96869
rect 4874 96858 4880 96860
rect 4936 96858 4960 96860
rect 5016 96858 5040 96860
rect 5096 96858 5120 96860
rect 5176 96858 5182 96860
rect 4936 96806 4938 96858
rect 5118 96806 5120 96858
rect 4874 96804 4880 96806
rect 4936 96804 4960 96806
rect 5016 96804 5040 96806
rect 5096 96804 5120 96806
rect 5176 96804 5182 96806
rect 4874 96795 5182 96804
rect 1306 96656 1362 96665
rect 1306 96591 1362 96600
rect 4214 96316 4522 96325
rect 4214 96314 4220 96316
rect 4276 96314 4300 96316
rect 4356 96314 4380 96316
rect 4436 96314 4460 96316
rect 4516 96314 4522 96316
rect 4276 96262 4278 96314
rect 4458 96262 4460 96314
rect 4214 96260 4220 96262
rect 4276 96260 4300 96262
rect 4356 96260 4380 96262
rect 4436 96260 4460 96262
rect 4516 96260 4522 96262
rect 4214 96251 4522 96260
rect 1216 96008 1268 96014
rect 1214 95976 1216 95985
rect 1268 95976 1270 95985
rect 1214 95911 1270 95920
rect 4874 95772 5182 95781
rect 4874 95770 4880 95772
rect 4936 95770 4960 95772
rect 5016 95770 5040 95772
rect 5096 95770 5120 95772
rect 5176 95770 5182 95772
rect 4936 95718 4938 95770
rect 5118 95718 5120 95770
rect 4874 95716 4880 95718
rect 4936 95716 4960 95718
rect 5016 95716 5040 95718
rect 5096 95716 5120 95718
rect 5176 95716 5182 95718
rect 4874 95707 5182 95716
rect 4214 95228 4522 95237
rect 4214 95226 4220 95228
rect 4276 95226 4300 95228
rect 4356 95226 4380 95228
rect 4436 95226 4460 95228
rect 4516 95226 4522 95228
rect 4276 95174 4278 95226
rect 4458 95174 4460 95226
rect 4214 95172 4220 95174
rect 4276 95172 4300 95174
rect 4356 95172 4380 95174
rect 4436 95172 4460 95174
rect 4516 95172 4522 95174
rect 4214 95163 4522 95172
rect 4874 94684 5182 94693
rect 4874 94682 4880 94684
rect 4936 94682 4960 94684
rect 5016 94682 5040 94684
rect 5096 94682 5120 94684
rect 5176 94682 5182 94684
rect 4936 94630 4938 94682
rect 5118 94630 5120 94682
rect 4874 94628 4880 94630
rect 4936 94628 4960 94630
rect 5016 94628 5040 94630
rect 5096 94628 5120 94630
rect 5176 94628 5182 94630
rect 4874 94619 5182 94628
rect 1308 94444 1360 94450
rect 1308 94386 1360 94392
rect 1320 93945 1348 94386
rect 4214 94140 4522 94149
rect 4214 94138 4220 94140
rect 4276 94138 4300 94140
rect 4356 94138 4380 94140
rect 4436 94138 4460 94140
rect 4516 94138 4522 94140
rect 4276 94086 4278 94138
rect 4458 94086 4460 94138
rect 4214 94084 4220 94086
rect 4276 94084 4300 94086
rect 4356 94084 4380 94086
rect 4436 94084 4460 94086
rect 4516 94084 4522 94086
rect 4214 94075 4522 94084
rect 1306 93936 1362 93945
rect 1306 93871 1362 93880
rect 4874 93596 5182 93605
rect 4874 93594 4880 93596
rect 4936 93594 4960 93596
rect 5016 93594 5040 93596
rect 5096 93594 5120 93596
rect 5176 93594 5182 93596
rect 4936 93542 4938 93594
rect 5118 93542 5120 93594
rect 4874 93540 4880 93542
rect 4936 93540 4960 93542
rect 5016 93540 5040 93542
rect 5096 93540 5120 93542
rect 5176 93540 5182 93542
rect 4874 93531 5182 93540
rect 4214 93052 4522 93061
rect 4214 93050 4220 93052
rect 4276 93050 4300 93052
rect 4356 93050 4380 93052
rect 4436 93050 4460 93052
rect 4516 93050 4522 93052
rect 4276 92998 4278 93050
rect 4458 92998 4460 93050
rect 4214 92996 4220 92998
rect 4276 92996 4300 92998
rect 4356 92996 4380 92998
rect 4436 92996 4460 92998
rect 4516 92996 4522 92998
rect 4214 92987 4522 92996
rect 4874 92508 5182 92517
rect 4874 92506 4880 92508
rect 4936 92506 4960 92508
rect 5016 92506 5040 92508
rect 5096 92506 5120 92508
rect 5176 92506 5182 92508
rect 4936 92454 4938 92506
rect 5118 92454 5120 92506
rect 4874 92452 4880 92454
rect 4936 92452 4960 92454
rect 5016 92452 5040 92454
rect 5096 92452 5120 92454
rect 5176 92452 5182 92454
rect 4874 92443 5182 92452
rect 4214 91964 4522 91973
rect 4214 91962 4220 91964
rect 4276 91962 4300 91964
rect 4356 91962 4380 91964
rect 4436 91962 4460 91964
rect 4516 91962 4522 91964
rect 4276 91910 4278 91962
rect 4458 91910 4460 91962
rect 4214 91908 4220 91910
rect 4276 91908 4300 91910
rect 4356 91908 4380 91910
rect 4436 91908 4460 91910
rect 4516 91908 4522 91910
rect 4214 91899 4522 91908
rect 4874 91420 5182 91429
rect 4874 91418 4880 91420
rect 4936 91418 4960 91420
rect 5016 91418 5040 91420
rect 5096 91418 5120 91420
rect 5176 91418 5182 91420
rect 4936 91366 4938 91418
rect 5118 91366 5120 91418
rect 4874 91364 4880 91366
rect 4936 91364 4960 91366
rect 5016 91364 5040 91366
rect 5096 91364 5120 91366
rect 5176 91364 5182 91366
rect 4874 91355 5182 91364
rect 4214 90876 4522 90885
rect 4214 90874 4220 90876
rect 4276 90874 4300 90876
rect 4356 90874 4380 90876
rect 4436 90874 4460 90876
rect 4516 90874 4522 90876
rect 4276 90822 4278 90874
rect 4458 90822 4460 90874
rect 4214 90820 4220 90822
rect 4276 90820 4300 90822
rect 4356 90820 4380 90822
rect 4436 90820 4460 90822
rect 4516 90820 4522 90822
rect 4214 90811 4522 90820
rect 4874 90332 5182 90341
rect 4874 90330 4880 90332
rect 4936 90330 4960 90332
rect 5016 90330 5040 90332
rect 5096 90330 5120 90332
rect 5176 90330 5182 90332
rect 4936 90278 4938 90330
rect 5118 90278 5120 90330
rect 4874 90276 4880 90278
rect 4936 90276 4960 90278
rect 5016 90276 5040 90278
rect 5096 90276 5120 90278
rect 5176 90276 5182 90278
rect 4874 90267 5182 90276
rect 4214 89788 4522 89797
rect 4214 89786 4220 89788
rect 4276 89786 4300 89788
rect 4356 89786 4380 89788
rect 4436 89786 4460 89788
rect 4516 89786 4522 89788
rect 4276 89734 4278 89786
rect 4458 89734 4460 89786
rect 4214 89732 4220 89734
rect 4276 89732 4300 89734
rect 4356 89732 4380 89734
rect 4436 89732 4460 89734
rect 4516 89732 4522 89734
rect 4214 89723 4522 89732
rect 4874 89244 5182 89253
rect 4874 89242 4880 89244
rect 4936 89242 4960 89244
rect 5016 89242 5040 89244
rect 5096 89242 5120 89244
rect 5176 89242 5182 89244
rect 4936 89190 4938 89242
rect 5118 89190 5120 89242
rect 4874 89188 4880 89190
rect 4936 89188 4960 89190
rect 5016 89188 5040 89190
rect 5096 89188 5120 89190
rect 5176 89188 5182 89190
rect 4874 89179 5182 89188
rect 4214 88700 4522 88709
rect 4214 88698 4220 88700
rect 4276 88698 4300 88700
rect 4356 88698 4380 88700
rect 4436 88698 4460 88700
rect 4516 88698 4522 88700
rect 4276 88646 4278 88698
rect 4458 88646 4460 88698
rect 4214 88644 4220 88646
rect 4276 88644 4300 88646
rect 4356 88644 4380 88646
rect 4436 88644 4460 88646
rect 4516 88644 4522 88646
rect 4214 88635 4522 88644
rect 4874 88156 5182 88165
rect 4874 88154 4880 88156
rect 4936 88154 4960 88156
rect 5016 88154 5040 88156
rect 5096 88154 5120 88156
rect 5176 88154 5182 88156
rect 4936 88102 4938 88154
rect 5118 88102 5120 88154
rect 4874 88100 4880 88102
rect 4936 88100 4960 88102
rect 5016 88100 5040 88102
rect 5096 88100 5120 88102
rect 5176 88100 5182 88102
rect 4874 88091 5182 88100
rect 4214 87612 4522 87621
rect 4214 87610 4220 87612
rect 4276 87610 4300 87612
rect 4356 87610 4380 87612
rect 4436 87610 4460 87612
rect 4516 87610 4522 87612
rect 4276 87558 4278 87610
rect 4458 87558 4460 87610
rect 4214 87556 4220 87558
rect 4276 87556 4300 87558
rect 4356 87556 4380 87558
rect 4436 87556 4460 87558
rect 4516 87556 4522 87558
rect 4214 87547 4522 87556
rect 4874 87068 5182 87077
rect 4874 87066 4880 87068
rect 4936 87066 4960 87068
rect 5016 87066 5040 87068
rect 5096 87066 5120 87068
rect 5176 87066 5182 87068
rect 4936 87014 4938 87066
rect 5118 87014 5120 87066
rect 4874 87012 4880 87014
rect 4936 87012 4960 87014
rect 5016 87012 5040 87014
rect 5096 87012 5120 87014
rect 5176 87012 5182 87014
rect 4874 87003 5182 87012
rect 4214 86524 4522 86533
rect 4214 86522 4220 86524
rect 4276 86522 4300 86524
rect 4356 86522 4380 86524
rect 4436 86522 4460 86524
rect 4516 86522 4522 86524
rect 4276 86470 4278 86522
rect 4458 86470 4460 86522
rect 4214 86468 4220 86470
rect 4276 86468 4300 86470
rect 4356 86468 4380 86470
rect 4436 86468 4460 86470
rect 4516 86468 4522 86470
rect 4214 86459 4522 86468
rect 4874 85980 5182 85989
rect 4874 85978 4880 85980
rect 4936 85978 4960 85980
rect 5016 85978 5040 85980
rect 5096 85978 5120 85980
rect 5176 85978 5182 85980
rect 4936 85926 4938 85978
rect 5118 85926 5120 85978
rect 4874 85924 4880 85926
rect 4936 85924 4960 85926
rect 5016 85924 5040 85926
rect 5096 85924 5120 85926
rect 5176 85924 5182 85926
rect 4874 85915 5182 85924
rect 4214 85436 4522 85445
rect 4214 85434 4220 85436
rect 4276 85434 4300 85436
rect 4356 85434 4380 85436
rect 4436 85434 4460 85436
rect 4516 85434 4522 85436
rect 4276 85382 4278 85434
rect 4458 85382 4460 85434
rect 4214 85380 4220 85382
rect 4276 85380 4300 85382
rect 4356 85380 4380 85382
rect 4436 85380 4460 85382
rect 4516 85380 4522 85382
rect 4214 85371 4522 85380
rect 4874 84892 5182 84901
rect 4874 84890 4880 84892
rect 4936 84890 4960 84892
rect 5016 84890 5040 84892
rect 5096 84890 5120 84892
rect 5176 84890 5182 84892
rect 4936 84838 4938 84890
rect 5118 84838 5120 84890
rect 4874 84836 4880 84838
rect 4936 84836 4960 84838
rect 5016 84836 5040 84838
rect 5096 84836 5120 84838
rect 5176 84836 5182 84838
rect 4874 84827 5182 84836
rect 4214 84348 4522 84357
rect 4214 84346 4220 84348
rect 4276 84346 4300 84348
rect 4356 84346 4380 84348
rect 4436 84346 4460 84348
rect 4516 84346 4522 84348
rect 4276 84294 4278 84346
rect 4458 84294 4460 84346
rect 4214 84292 4220 84294
rect 4276 84292 4300 84294
rect 4356 84292 4380 84294
rect 4436 84292 4460 84294
rect 4516 84292 4522 84294
rect 4214 84283 4522 84292
rect 4874 83804 5182 83813
rect 4874 83802 4880 83804
rect 4936 83802 4960 83804
rect 5016 83802 5040 83804
rect 5096 83802 5120 83804
rect 5176 83802 5182 83804
rect 4936 83750 4938 83802
rect 5118 83750 5120 83802
rect 4874 83748 4880 83750
rect 4936 83748 4960 83750
rect 5016 83748 5040 83750
rect 5096 83748 5120 83750
rect 5176 83748 5182 83750
rect 4874 83739 5182 83748
rect 4214 83260 4522 83269
rect 4214 83258 4220 83260
rect 4276 83258 4300 83260
rect 4356 83258 4380 83260
rect 4436 83258 4460 83260
rect 4516 83258 4522 83260
rect 4276 83206 4278 83258
rect 4458 83206 4460 83258
rect 4214 83204 4220 83206
rect 4276 83204 4300 83206
rect 4356 83204 4380 83206
rect 4436 83204 4460 83206
rect 4516 83204 4522 83206
rect 4214 83195 4522 83204
rect 4874 82716 5182 82725
rect 4874 82714 4880 82716
rect 4936 82714 4960 82716
rect 5016 82714 5040 82716
rect 5096 82714 5120 82716
rect 5176 82714 5182 82716
rect 4936 82662 4938 82714
rect 5118 82662 5120 82714
rect 4874 82660 4880 82662
rect 4936 82660 4960 82662
rect 5016 82660 5040 82662
rect 5096 82660 5120 82662
rect 5176 82660 5182 82662
rect 4874 82651 5182 82660
rect 4214 82172 4522 82181
rect 4214 82170 4220 82172
rect 4276 82170 4300 82172
rect 4356 82170 4380 82172
rect 4436 82170 4460 82172
rect 4516 82170 4522 82172
rect 4276 82118 4278 82170
rect 4458 82118 4460 82170
rect 4214 82116 4220 82118
rect 4276 82116 4300 82118
rect 4356 82116 4380 82118
rect 4436 82116 4460 82118
rect 4516 82116 4522 82118
rect 4214 82107 4522 82116
rect 4874 81628 5182 81637
rect 4874 81626 4880 81628
rect 4936 81626 4960 81628
rect 5016 81626 5040 81628
rect 5096 81626 5120 81628
rect 5176 81626 5182 81628
rect 4936 81574 4938 81626
rect 5118 81574 5120 81626
rect 4874 81572 4880 81574
rect 4936 81572 4960 81574
rect 5016 81572 5040 81574
rect 5096 81572 5120 81574
rect 5176 81572 5182 81574
rect 4874 81563 5182 81572
rect 4214 81084 4522 81093
rect 4214 81082 4220 81084
rect 4276 81082 4300 81084
rect 4356 81082 4380 81084
rect 4436 81082 4460 81084
rect 4516 81082 4522 81084
rect 4276 81030 4278 81082
rect 4458 81030 4460 81082
rect 4214 81028 4220 81030
rect 4276 81028 4300 81030
rect 4356 81028 4380 81030
rect 4436 81028 4460 81030
rect 4516 81028 4522 81030
rect 4214 81019 4522 81028
rect 4874 80540 5182 80549
rect 4874 80538 4880 80540
rect 4936 80538 4960 80540
rect 5016 80538 5040 80540
rect 5096 80538 5120 80540
rect 5176 80538 5182 80540
rect 4936 80486 4938 80538
rect 5118 80486 5120 80538
rect 4874 80484 4880 80486
rect 4936 80484 4960 80486
rect 5016 80484 5040 80486
rect 5096 80484 5120 80486
rect 5176 80484 5182 80486
rect 4874 80475 5182 80484
rect 4214 79996 4522 80005
rect 4214 79994 4220 79996
rect 4276 79994 4300 79996
rect 4356 79994 4380 79996
rect 4436 79994 4460 79996
rect 4516 79994 4522 79996
rect 4276 79942 4278 79994
rect 4458 79942 4460 79994
rect 4214 79940 4220 79942
rect 4276 79940 4300 79942
rect 4356 79940 4380 79942
rect 4436 79940 4460 79942
rect 4516 79940 4522 79942
rect 4214 79931 4522 79940
rect 4874 79452 5182 79461
rect 4874 79450 4880 79452
rect 4936 79450 4960 79452
rect 5016 79450 5040 79452
rect 5096 79450 5120 79452
rect 5176 79450 5182 79452
rect 4936 79398 4938 79450
rect 5118 79398 5120 79450
rect 4874 79396 4880 79398
rect 4936 79396 4960 79398
rect 5016 79396 5040 79398
rect 5096 79396 5120 79398
rect 5176 79396 5182 79398
rect 4874 79387 5182 79396
rect 4214 78908 4522 78917
rect 4214 78906 4220 78908
rect 4276 78906 4300 78908
rect 4356 78906 4380 78908
rect 4436 78906 4460 78908
rect 4516 78906 4522 78908
rect 4276 78854 4278 78906
rect 4458 78854 4460 78906
rect 4214 78852 4220 78854
rect 4276 78852 4300 78854
rect 4356 78852 4380 78854
rect 4436 78852 4460 78854
rect 4516 78852 4522 78854
rect 4214 78843 4522 78852
rect 1308 78532 1360 78538
rect 1308 78474 1360 78480
rect 7564 78532 7616 78538
rect 7564 78474 7616 78480
rect 1320 78305 1348 78474
rect 4874 78364 5182 78373
rect 4874 78362 4880 78364
rect 4936 78362 4960 78364
rect 5016 78362 5040 78364
rect 5096 78362 5120 78364
rect 5176 78362 5182 78364
rect 4936 78310 4938 78362
rect 5118 78310 5120 78362
rect 4874 78308 4880 78310
rect 4936 78308 4960 78310
rect 5016 78308 5040 78310
rect 5096 78308 5120 78310
rect 5176 78308 5182 78310
rect 1306 78296 1362 78305
rect 4874 78299 5182 78308
rect 1306 78231 1362 78240
rect 1308 78124 1360 78130
rect 1308 78066 1360 78072
rect 1320 77625 1348 78066
rect 4214 77820 4522 77829
rect 4214 77818 4220 77820
rect 4276 77818 4300 77820
rect 4356 77818 4380 77820
rect 4436 77818 4460 77820
rect 4516 77818 4522 77820
rect 4276 77766 4278 77818
rect 4458 77766 4460 77818
rect 4214 77764 4220 77766
rect 4276 77764 4300 77766
rect 4356 77764 4380 77766
rect 4436 77764 4460 77766
rect 4516 77764 4522 77766
rect 4214 77755 4522 77764
rect 1306 77616 1362 77625
rect 1306 77551 1362 77560
rect 4874 77276 5182 77285
rect 4874 77274 4880 77276
rect 4936 77274 4960 77276
rect 5016 77274 5040 77276
rect 5096 77274 5120 77276
rect 5176 77274 5182 77276
rect 4936 77222 4938 77274
rect 5118 77222 5120 77274
rect 4874 77220 4880 77222
rect 4936 77220 4960 77222
rect 5016 77220 5040 77222
rect 5096 77220 5120 77222
rect 5176 77220 5182 77222
rect 4874 77211 5182 77220
rect 1216 77036 1268 77042
rect 1216 76978 1268 76984
rect 1228 76945 1256 76978
rect 1214 76936 1270 76945
rect 1214 76871 1270 76880
rect 4214 76732 4522 76741
rect 4214 76730 4220 76732
rect 4276 76730 4300 76732
rect 4356 76730 4380 76732
rect 4436 76730 4460 76732
rect 4516 76730 4522 76732
rect 4276 76678 4278 76730
rect 4458 76678 4460 76730
rect 4214 76676 4220 76678
rect 4276 76676 4300 76678
rect 4356 76676 4380 76678
rect 4436 76676 4460 76678
rect 4516 76676 4522 76678
rect 4214 76667 4522 76676
rect 1216 76356 1268 76362
rect 1216 76298 1268 76304
rect 1228 76265 1256 76298
rect 1214 76256 1270 76265
rect 1214 76191 1270 76200
rect 4874 76188 5182 76197
rect 4874 76186 4880 76188
rect 4936 76186 4960 76188
rect 5016 76186 5040 76188
rect 5096 76186 5120 76188
rect 5176 76186 5182 76188
rect 4936 76134 4938 76186
rect 5118 76134 5120 76186
rect 4874 76132 4880 76134
rect 4936 76132 4960 76134
rect 5016 76132 5040 76134
rect 5096 76132 5120 76134
rect 5176 76132 5182 76134
rect 4874 76123 5182 76132
rect 5540 76084 5592 76090
rect 5540 76026 5592 76032
rect 1400 75948 1452 75954
rect 1400 75890 1452 75896
rect 1412 75585 1440 75890
rect 4214 75644 4522 75653
rect 4214 75642 4220 75644
rect 4276 75642 4300 75644
rect 4356 75642 4380 75644
rect 4436 75642 4460 75644
rect 4516 75642 4522 75644
rect 4276 75590 4278 75642
rect 4458 75590 4460 75642
rect 4214 75588 4220 75590
rect 4276 75588 4300 75590
rect 4356 75588 4380 75590
rect 4436 75588 4460 75590
rect 4516 75588 4522 75590
rect 1398 75576 1454 75585
rect 4214 75579 4522 75588
rect 5552 75585 5580 76026
rect 1398 75511 1454 75520
rect 5538 75576 5594 75585
rect 5538 75511 5594 75520
rect 1308 75268 1360 75274
rect 1308 75210 1360 75216
rect 6920 75268 6972 75274
rect 6920 75210 6972 75216
rect 1320 74905 1348 75210
rect 4874 75100 5182 75109
rect 4874 75098 4880 75100
rect 4936 75098 4960 75100
rect 5016 75098 5040 75100
rect 5096 75098 5120 75100
rect 5176 75098 5182 75100
rect 4936 75046 4938 75098
rect 5118 75046 5120 75098
rect 4874 75044 4880 75046
rect 4936 75044 4960 75046
rect 5016 75044 5040 75046
rect 5096 75044 5120 75046
rect 5176 75044 5182 75046
rect 4874 75035 5182 75044
rect 1306 74896 1362 74905
rect 1306 74831 1362 74840
rect 4214 74556 4522 74565
rect 4214 74554 4220 74556
rect 4276 74554 4300 74556
rect 4356 74554 4380 74556
rect 4436 74554 4460 74556
rect 4516 74554 4522 74556
rect 4276 74502 4278 74554
rect 4458 74502 4460 74554
rect 4214 74500 4220 74502
rect 4276 74500 4300 74502
rect 4356 74500 4380 74502
rect 4436 74500 4460 74502
rect 4516 74500 4522 74502
rect 4214 74491 4522 74500
rect 1214 74216 1270 74225
rect 1214 74151 1216 74160
rect 1268 74151 1270 74160
rect 1216 74122 1268 74128
rect 1860 74112 1912 74118
rect 1860 74054 1912 74060
rect 1308 73772 1360 73778
rect 1308 73714 1360 73720
rect 1320 73545 1348 73714
rect 1306 73536 1362 73545
rect 1306 73471 1362 73480
rect 1492 73092 1544 73098
rect 1492 73034 1544 73040
rect 1504 72865 1532 73034
rect 1490 72856 1546 72865
rect 1490 72791 1546 72800
rect 1308 72684 1360 72690
rect 1308 72626 1360 72632
rect 1320 72185 1348 72626
rect 1306 72176 1362 72185
rect 1306 72111 1362 72120
rect 1872 71738 1900 74054
rect 4874 74012 5182 74021
rect 4874 74010 4880 74012
rect 4936 74010 4960 74012
rect 5016 74010 5040 74012
rect 5096 74010 5120 74012
rect 5176 74010 5182 74012
rect 4936 73958 4938 74010
rect 5118 73958 5120 74010
rect 4874 73956 4880 73958
rect 4936 73956 4960 73958
rect 5016 73956 5040 73958
rect 5096 73956 5120 73958
rect 5176 73956 5182 73958
rect 4874 73947 5182 73956
rect 4214 73468 4522 73477
rect 4214 73466 4220 73468
rect 4276 73466 4300 73468
rect 4356 73466 4380 73468
rect 4436 73466 4460 73468
rect 4516 73466 4522 73468
rect 4276 73414 4278 73466
rect 4458 73414 4460 73466
rect 4214 73412 4220 73414
rect 4276 73412 4300 73414
rect 4356 73412 4380 73414
rect 4436 73412 4460 73414
rect 4516 73412 4522 73414
rect 4214 73403 4522 73412
rect 4874 72924 5182 72933
rect 4874 72922 4880 72924
rect 4936 72922 4960 72924
rect 5016 72922 5040 72924
rect 5096 72922 5120 72924
rect 5176 72922 5182 72924
rect 4936 72870 4938 72922
rect 5118 72870 5120 72922
rect 4874 72868 4880 72870
rect 4936 72868 4960 72870
rect 5016 72868 5040 72870
rect 5096 72868 5120 72870
rect 5176 72868 5182 72870
rect 4874 72859 5182 72868
rect 4214 72380 4522 72389
rect 4214 72378 4220 72380
rect 4276 72378 4300 72380
rect 4356 72378 4380 72380
rect 4436 72378 4460 72380
rect 4516 72378 4522 72380
rect 4276 72326 4278 72378
rect 4458 72326 4460 72378
rect 4214 72324 4220 72326
rect 4276 72324 4300 72326
rect 4356 72324 4380 72326
rect 4436 72324 4460 72326
rect 4516 72324 4522 72326
rect 4214 72315 4522 72324
rect 4874 71836 5182 71845
rect 4874 71834 4880 71836
rect 4936 71834 4960 71836
rect 5016 71834 5040 71836
rect 5096 71834 5120 71836
rect 5176 71834 5182 71836
rect 4936 71782 4938 71834
rect 5118 71782 5120 71834
rect 4874 71780 4880 71782
rect 4936 71780 4960 71782
rect 5016 71780 5040 71782
rect 5096 71780 5120 71782
rect 5176 71780 5182 71782
rect 4874 71771 5182 71780
rect 1860 71732 1912 71738
rect 1860 71674 1912 71680
rect 1216 71596 1268 71602
rect 1216 71538 1268 71544
rect 1228 71505 1256 71538
rect 1214 71496 1270 71505
rect 1214 71431 1270 71440
rect 1860 71392 1912 71398
rect 1860 71334 1912 71340
rect 1308 70916 1360 70922
rect 1308 70858 1360 70864
rect 1320 70825 1348 70858
rect 1306 70816 1362 70825
rect 1306 70751 1362 70760
rect 1872 70038 1900 71334
rect 4214 71292 4522 71301
rect 4214 71290 4220 71292
rect 4276 71290 4300 71292
rect 4356 71290 4380 71292
rect 4436 71290 4460 71292
rect 4516 71290 4522 71292
rect 4276 71238 4278 71290
rect 4458 71238 4460 71290
rect 4214 71236 4220 71238
rect 4276 71236 4300 71238
rect 4356 71236 4380 71238
rect 4436 71236 4460 71238
rect 4516 71236 4522 71238
rect 4214 71227 4522 71236
rect 2228 70848 2280 70854
rect 2228 70790 2280 70796
rect 2240 70446 2268 70790
rect 4874 70748 5182 70757
rect 4874 70746 4880 70748
rect 4936 70746 4960 70748
rect 5016 70746 5040 70748
rect 5096 70746 5120 70748
rect 5176 70746 5182 70748
rect 4936 70694 4938 70746
rect 5118 70694 5120 70746
rect 4874 70692 4880 70694
rect 4936 70692 4960 70694
rect 5016 70692 5040 70694
rect 5096 70692 5120 70694
rect 5176 70692 5182 70694
rect 4874 70683 5182 70692
rect 2228 70440 2280 70446
rect 2228 70382 2280 70388
rect 2240 70145 2268 70382
rect 4214 70204 4522 70213
rect 4214 70202 4220 70204
rect 4276 70202 4300 70204
rect 4356 70202 4380 70204
rect 4436 70202 4460 70204
rect 4516 70202 4522 70204
rect 4276 70150 4278 70202
rect 4458 70150 4460 70202
rect 4214 70148 4220 70150
rect 4276 70148 4300 70150
rect 4356 70148 4380 70150
rect 4436 70148 4460 70150
rect 4516 70148 4522 70150
rect 2226 70136 2282 70145
rect 4214 70139 4522 70148
rect 2226 70071 2282 70080
rect 1860 70032 1912 70038
rect 1860 69974 1912 69980
rect 1308 69828 1360 69834
rect 1308 69770 1360 69776
rect 1320 69465 1348 69770
rect 4874 69660 5182 69669
rect 4874 69658 4880 69660
rect 4936 69658 4960 69660
rect 5016 69658 5040 69660
rect 5096 69658 5120 69660
rect 5176 69658 5182 69660
rect 4936 69606 4938 69658
rect 5118 69606 5120 69658
rect 4874 69604 4880 69606
rect 4936 69604 4960 69606
rect 5016 69604 5040 69606
rect 5096 69604 5120 69606
rect 5176 69604 5182 69606
rect 4874 69595 5182 69604
rect 1306 69456 1362 69465
rect 6932 69426 6960 75210
rect 7576 69494 7604 78474
rect 7656 77988 7708 77994
rect 7656 77930 7708 77936
rect 7668 69562 7696 77930
rect 7656 69556 7708 69562
rect 7656 69498 7708 69504
rect 7564 69488 7616 69494
rect 7564 69430 7616 69436
rect 1306 69391 1362 69400
rect 6920 69420 6972 69426
rect 6920 69362 6972 69368
rect 4214 69116 4522 69125
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69051 4522 69060
rect 1214 68776 1270 68785
rect 1214 68711 1216 68720
rect 1268 68711 1270 68720
rect 1216 68682 1268 68688
rect 4874 68572 5182 68581
rect 4874 68570 4880 68572
rect 4936 68570 4960 68572
rect 5016 68570 5040 68572
rect 5096 68570 5120 68572
rect 5176 68570 5182 68572
rect 4936 68518 4938 68570
rect 5118 68518 5120 68570
rect 4874 68516 4880 68518
rect 4936 68516 4960 68518
rect 5016 68516 5040 68518
rect 5096 68516 5120 68518
rect 5176 68516 5182 68518
rect 4874 68507 5182 68516
rect 7852 68474 7880 125802
rect 7840 68468 7892 68474
rect 7840 68410 7892 68416
rect 7944 68406 7972 125870
rect 8024 125724 8076 125730
rect 8024 125666 8076 125672
rect 7932 68400 7984 68406
rect 7932 68342 7984 68348
rect 1308 68332 1360 68338
rect 1308 68274 1360 68280
rect 1320 68105 1348 68274
rect 2044 68264 2096 68270
rect 2044 68206 2096 68212
rect 1306 68096 1362 68105
rect 1306 68031 1362 68040
rect 2056 67930 2084 68206
rect 4214 68028 4522 68037
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67963 4522 67972
rect 2044 67924 2096 67930
rect 2044 67866 2096 67872
rect 1676 67856 1728 67862
rect 1676 67798 1728 67804
rect 1124 67652 1176 67658
rect 1124 67594 1176 67600
rect 1136 67425 1164 67594
rect 1122 67416 1178 67425
rect 1122 67351 1178 67360
rect 848 67040 900 67046
rect 848 66982 900 66988
rect 860 66881 888 66982
rect 846 66872 902 66881
rect 846 66807 902 66816
rect 848 65952 900 65958
rect 846 65920 848 65929
rect 900 65920 902 65929
rect 846 65855 902 65864
rect 846 65512 902 65521
rect 846 65447 902 65456
rect 860 65414 888 65447
rect 848 65408 900 65414
rect 848 65350 900 65356
rect 1400 64932 1452 64938
rect 1400 64874 1452 64880
rect 1412 64705 1440 64874
rect 1398 64696 1454 64705
rect 1398 64631 1454 64640
rect 848 64320 900 64326
rect 848 64262 900 64268
rect 860 64161 888 64262
rect 846 64152 902 64161
rect 846 64087 902 64096
rect 848 63504 900 63510
rect 846 63472 848 63481
rect 900 63472 902 63481
rect 846 63407 902 63416
rect 846 62792 902 62801
rect 846 62727 848 62736
rect 900 62727 902 62736
rect 848 62698 900 62704
rect 1492 62212 1544 62218
rect 1492 62154 1544 62160
rect 1504 61985 1532 62154
rect 1490 61976 1546 61985
rect 1490 61911 1546 61920
rect 1688 61878 1716 67798
rect 4874 67484 5182 67493
rect 4874 67482 4880 67484
rect 4936 67482 4960 67484
rect 5016 67482 5040 67484
rect 5096 67482 5120 67484
rect 5176 67482 5182 67484
rect 4936 67430 4938 67482
rect 5118 67430 5120 67482
rect 4874 67428 4880 67430
rect 4936 67428 4960 67430
rect 5016 67428 5040 67430
rect 5096 67428 5120 67430
rect 5176 67428 5182 67430
rect 4874 67419 5182 67428
rect 8036 67289 8064 125666
rect 8022 67280 8078 67289
rect 8022 67215 8078 67224
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 2780 66836 2832 66842
rect 2780 66778 2832 66784
rect 1860 64320 1912 64326
rect 1860 64262 1912 64268
rect 1872 62490 1900 64262
rect 2792 63510 2820 66778
rect 3424 66768 3476 66774
rect 8128 66745 8156 125938
rect 8220 67425 8248 126006
rect 9496 125792 9548 125798
rect 9496 125734 9548 125740
rect 8392 101584 8444 101590
rect 8392 101526 8444 101532
rect 8404 101289 8432 101526
rect 8390 101280 8446 101289
rect 8390 101215 8446 101224
rect 8392 99748 8444 99754
rect 8392 99690 8444 99696
rect 8404 99521 8432 99690
rect 8390 99512 8446 99521
rect 8390 99447 8446 99456
rect 8392 98660 8444 98666
rect 8392 98602 8444 98608
rect 8404 98433 8432 98602
rect 8390 98424 8446 98433
rect 8390 98359 8446 98368
rect 8392 97232 8444 97238
rect 8392 97174 8444 97180
rect 8404 96801 8432 97174
rect 8390 96792 8446 96801
rect 8390 96727 8446 96736
rect 8392 96144 8444 96150
rect 8392 96086 8444 96092
rect 8404 95713 8432 96086
rect 8390 95704 8446 95713
rect 8390 95639 8446 95648
rect 8392 94308 8444 94314
rect 8392 94250 8444 94256
rect 8404 93945 8432 94250
rect 8390 93936 8446 93945
rect 8390 93871 8446 93880
rect 8944 76900 8996 76906
rect 8944 76842 8996 76848
rect 8852 76356 8904 76362
rect 8852 76298 8904 76304
rect 8392 70440 8444 70446
rect 8392 70382 8444 70388
rect 8404 67862 8432 70382
rect 8864 69601 8892 76298
rect 8956 69737 8984 76842
rect 9508 74534 9536 125734
rect 9324 74506 9536 74534
rect 9128 73772 9180 73778
rect 9128 73714 9180 73720
rect 9036 73228 9088 73234
rect 9036 73170 9088 73176
rect 9048 69902 9076 73170
rect 9036 69896 9088 69902
rect 9036 69838 9088 69844
rect 8942 69728 8998 69737
rect 8942 69663 8998 69672
rect 8850 69592 8906 69601
rect 8850 69527 8906 69536
rect 8392 67856 8444 67862
rect 8392 67798 8444 67804
rect 8206 67416 8262 67425
rect 8206 67351 8262 67360
rect 9140 67153 9168 73714
rect 9220 70984 9272 70990
rect 9220 70926 9272 70932
rect 9232 69873 9260 70926
rect 9218 69864 9274 69873
rect 9218 69799 9274 69808
rect 9324 68338 9352 74506
rect 9600 73778 9628 126074
rect 36096 124273 36124 126346
rect 36280 125798 36308 126346
rect 37648 126336 37700 126342
rect 37648 126278 37700 126284
rect 37660 125866 37688 126278
rect 37648 125860 37700 125866
rect 37648 125802 37700 125808
rect 36268 125792 36320 125798
rect 36268 125734 36320 125740
rect 37752 124273 37780 126346
rect 40960 126336 41012 126342
rect 40960 126278 41012 126284
rect 40972 125934 41000 126278
rect 40960 125928 41012 125934
rect 40960 125870 41012 125876
rect 41340 124273 41368 126346
rect 41420 126336 41472 126342
rect 41420 126278 41472 126284
rect 41432 126002 41460 126278
rect 41420 125996 41472 126002
rect 41420 125938 41472 125944
rect 36082 124264 36138 124273
rect 36082 124199 36138 124208
rect 37738 124264 37794 124273
rect 37738 124199 37794 124208
rect 41326 124264 41382 124273
rect 41326 124199 41382 124208
rect 42352 124137 42380 126414
rect 45192 126404 45244 126410
rect 45192 126346 45244 126352
rect 48504 126404 48556 126410
rect 48504 126346 48556 126352
rect 49700 126404 49752 126410
rect 49700 126346 49752 126352
rect 56784 126404 56836 126410
rect 56784 126346 56836 126352
rect 59360 126404 59412 126410
rect 59360 126346 59412 126352
rect 61844 126404 61896 126410
rect 61844 126346 61896 126352
rect 63960 126404 64012 126410
rect 63960 126346 64012 126352
rect 64420 126404 64472 126410
rect 64420 126346 64472 126352
rect 66076 126404 66128 126410
rect 66076 126346 66128 126352
rect 68560 126404 68612 126410
rect 68560 126346 68612 126352
rect 71412 126404 71464 126410
rect 77298 126375 77300 126384
rect 71412 126346 71464 126352
rect 77352 126375 77354 126384
rect 77300 126346 77352 126352
rect 45100 126336 45152 126342
rect 45100 126278 45152 126284
rect 45112 126070 45140 126278
rect 45100 126064 45152 126070
rect 45204 126041 45232 126346
rect 48412 126336 48464 126342
rect 48412 126278 48464 126284
rect 45100 126006 45152 126012
rect 45190 126032 45246 126041
rect 45190 125967 45246 125976
rect 48424 125730 48452 126278
rect 48412 125724 48464 125730
rect 48412 125666 48464 125672
rect 48516 124273 48544 126346
rect 49608 126336 49660 126342
rect 49608 126278 49660 126284
rect 49620 126138 49648 126278
rect 49608 126132 49660 126138
rect 49608 126074 49660 126080
rect 49712 125633 49740 126346
rect 56796 126041 56824 126346
rect 56782 126032 56838 126041
rect 56782 125967 56838 125976
rect 59372 125633 59400 126346
rect 59728 126336 59780 126342
rect 59728 126278 59780 126284
rect 59740 126138 59768 126278
rect 59728 126132 59780 126138
rect 59728 126074 59780 126080
rect 61856 125769 61884 126346
rect 62212 126336 62264 126342
rect 62212 126278 62264 126284
rect 62224 126070 62252 126278
rect 62212 126064 62264 126070
rect 62212 126006 62264 126012
rect 61842 125760 61898 125769
rect 61842 125695 61898 125704
rect 63972 125633 64000 126346
rect 64328 126336 64380 126342
rect 64328 126278 64380 126284
rect 64340 126002 64368 126278
rect 64328 125996 64380 126002
rect 64328 125938 64380 125944
rect 49698 125624 49754 125633
rect 49698 125559 49754 125568
rect 59358 125624 59414 125633
rect 59358 125559 59414 125568
rect 63958 125624 64014 125633
rect 63958 125559 64014 125568
rect 64432 125225 64460 126346
rect 65984 126336 66036 126342
rect 65984 126278 66036 126284
rect 65996 125934 66024 126278
rect 65984 125928 66036 125934
rect 65984 125870 66036 125876
rect 64418 125216 64474 125225
rect 64418 125151 64474 125160
rect 66088 124273 66116 126346
rect 67088 126336 67140 126342
rect 67088 126278 67140 126284
rect 66314 126236 66622 126245
rect 66314 126234 66320 126236
rect 66376 126234 66400 126236
rect 66456 126234 66480 126236
rect 66536 126234 66560 126236
rect 66616 126234 66622 126236
rect 66376 126182 66378 126234
rect 66558 126182 66560 126234
rect 66314 126180 66320 126182
rect 66376 126180 66400 126182
rect 66456 126180 66480 126182
rect 66536 126180 66560 126182
rect 66616 126180 66622 126182
rect 66314 126171 66622 126180
rect 67100 125866 67128 126278
rect 67088 125860 67140 125866
rect 67088 125802 67140 125808
rect 68572 124273 68600 126346
rect 70860 126336 70912 126342
rect 70860 126278 70912 126284
rect 70872 125730 70900 126278
rect 70860 125724 70912 125730
rect 70860 125666 70912 125672
rect 71424 124273 71452 126346
rect 71780 126336 71832 126342
rect 71780 126278 71832 126284
rect 86316 126336 86368 126342
rect 86316 126278 86368 126284
rect 87328 126336 87380 126342
rect 87328 126278 87380 126284
rect 96068 126336 96120 126342
rect 96068 126278 96120 126284
rect 71792 125798 71820 126278
rect 71780 125792 71832 125798
rect 71780 125734 71832 125740
rect 48502 124264 48558 124273
rect 48502 124199 48558 124208
rect 66074 124264 66130 124273
rect 66074 124199 66130 124208
rect 68558 124264 68614 124273
rect 68558 124199 68614 124208
rect 71410 124264 71466 124273
rect 71410 124199 71466 124208
rect 42338 124128 42394 124137
rect 42338 124063 42394 124072
rect 86328 124001 86356 126278
rect 86314 123992 86370 124001
rect 86314 123927 86370 123936
rect 87340 123865 87368 126278
rect 96080 123865 96108 126278
rect 97034 126236 97342 126245
rect 97034 126234 97040 126236
rect 97096 126234 97120 126236
rect 97176 126234 97200 126236
rect 97256 126234 97280 126236
rect 97336 126234 97342 126236
rect 97096 126182 97098 126234
rect 97278 126182 97280 126234
rect 97034 126180 97040 126182
rect 97096 126180 97120 126182
rect 97176 126180 97200 126182
rect 97256 126180 97280 126182
rect 97336 126180 97342 126182
rect 97034 126171 97342 126180
rect 87326 123856 87382 123865
rect 87326 123791 87382 123800
rect 96066 123856 96122 123865
rect 96066 123791 96122 123800
rect 87340 123758 87368 123791
rect 87328 123752 87380 123758
rect 87328 123694 87380 123700
rect 102046 83388 102102 83397
rect 101968 83346 102046 83374
rect 9588 73772 9640 73778
rect 9588 73714 9640 73720
rect 9588 73636 9640 73642
rect 9588 73578 9640 73584
rect 9496 72548 9548 72554
rect 9496 72490 9548 72496
rect 9404 71732 9456 71738
rect 9404 71674 9456 71680
rect 9416 69465 9444 71674
rect 9508 69834 9536 72490
rect 9600 69970 9628 73578
rect 38660 70032 38712 70038
rect 38660 69974 38712 69980
rect 73620 70032 73672 70038
rect 73620 69974 73672 69980
rect 9588 69964 9640 69970
rect 9588 69906 9640 69912
rect 38672 69873 38700 69974
rect 43260 69964 43312 69970
rect 43260 69906 43312 69912
rect 71780 69964 71832 69970
rect 71780 69906 71832 69912
rect 40960 69896 41012 69902
rect 37462 69864 37518 69873
rect 9496 69828 9548 69834
rect 37462 69799 37518 69808
rect 38658 69864 38714 69873
rect 38658 69799 38714 69808
rect 39762 69864 39818 69873
rect 39762 69799 39764 69808
rect 9496 69770 9548 69776
rect 37476 69766 37504 69799
rect 37464 69760 37516 69766
rect 37464 69702 37516 69708
rect 23294 69592 23350 69601
rect 23294 69527 23350 69536
rect 23478 69592 23534 69601
rect 23478 69527 23534 69536
rect 24674 69592 24730 69601
rect 24674 69527 24730 69536
rect 25778 69592 25834 69601
rect 25778 69527 25834 69536
rect 26974 69592 27030 69601
rect 26974 69527 27030 69536
rect 28078 69592 28134 69601
rect 28078 69527 28134 69536
rect 30470 69592 30526 69601
rect 30470 69527 30526 69536
rect 31758 69592 31814 69601
rect 31758 69527 31814 69536
rect 32862 69592 32918 69601
rect 32862 69527 32864 69536
rect 9402 69456 9458 69465
rect 9402 69391 9458 69400
rect 23308 69329 23336 69527
rect 23294 69320 23350 69329
rect 23294 69255 23350 69264
rect 9312 68332 9364 68338
rect 9312 68274 9364 68280
rect 23492 67930 23520 69527
rect 24688 67930 24716 69527
rect 25792 68134 25820 69527
rect 25780 68128 25832 68134
rect 25780 68070 25832 68076
rect 25792 67930 25820 68070
rect 26988 67930 27016 69527
rect 23480 67924 23532 67930
rect 23480 67866 23532 67872
rect 24676 67924 24728 67930
rect 24676 67866 24728 67872
rect 25780 67924 25832 67930
rect 25780 67866 25832 67872
rect 26976 67924 27028 67930
rect 26976 67866 27028 67872
rect 28092 67794 28120 69527
rect 29550 69320 29606 69329
rect 29550 69255 29606 69264
rect 29564 67930 29592 69255
rect 30484 68202 30512 69527
rect 30472 68196 30524 68202
rect 30472 68138 30524 68144
rect 30484 67930 30512 68138
rect 31772 67930 31800 69527
rect 32916 69527 32918 69536
rect 33966 69592 34022 69601
rect 33966 69527 34022 69536
rect 35162 69592 35218 69601
rect 35162 69527 35218 69536
rect 36358 69592 36414 69601
rect 36358 69527 36414 69536
rect 32864 69498 32916 69504
rect 32876 67930 32904 69498
rect 33600 68468 33652 68474
rect 33600 68410 33652 68416
rect 29552 67924 29604 67930
rect 29552 67866 29604 67872
rect 30472 67924 30524 67930
rect 30472 67866 30524 67872
rect 31760 67924 31812 67930
rect 31760 67866 31812 67872
rect 32864 67924 32916 67930
rect 32864 67866 32916 67872
rect 10324 67788 10376 67794
rect 10324 67730 10376 67736
rect 28080 67788 28132 67794
rect 28080 67730 28132 67736
rect 9126 67144 9182 67153
rect 9126 67079 9182 67088
rect 3424 66710 3476 66716
rect 8114 66736 8170 66745
rect 2780 63504 2832 63510
rect 2780 63446 2832 63452
rect 3436 63034 3464 66710
rect 8114 66671 8170 66680
rect 4874 66396 5182 66405
rect 4874 66394 4880 66396
rect 4936 66394 4960 66396
rect 5016 66394 5040 66396
rect 5096 66394 5120 66396
rect 5176 66394 5182 66396
rect 4936 66342 4938 66394
rect 5118 66342 5120 66394
rect 4874 66340 4880 66342
rect 4936 66340 4960 66342
rect 5016 66340 5040 66342
rect 5096 66340 5120 66342
rect 5176 66340 5182 66342
rect 4874 66331 5182 66340
rect 9588 66292 9640 66298
rect 9588 66234 9640 66240
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 4874 65308 5182 65317
rect 4874 65306 4880 65308
rect 4936 65306 4960 65308
rect 5016 65306 5040 65308
rect 5096 65306 5120 65308
rect 5176 65306 5182 65308
rect 4936 65254 4938 65306
rect 5118 65254 5120 65306
rect 4874 65252 4880 65254
rect 4936 65252 4960 65254
rect 5016 65252 5040 65254
rect 5096 65252 5120 65254
rect 5176 65252 5182 65254
rect 4874 65243 5182 65252
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 4874 64220 5182 64229
rect 4874 64218 4880 64220
rect 4936 64218 4960 64220
rect 5016 64218 5040 64220
rect 5096 64218 5120 64220
rect 5176 64218 5182 64220
rect 4936 64166 4938 64218
rect 5118 64166 5120 64218
rect 4874 64164 4880 64166
rect 4936 64164 4960 64166
rect 5016 64164 5040 64166
rect 5096 64164 5120 64166
rect 5176 64164 5182 64166
rect 4874 64155 5182 64164
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 4874 63132 5182 63141
rect 4874 63130 4880 63132
rect 4936 63130 4960 63132
rect 5016 63130 5040 63132
rect 5096 63130 5120 63132
rect 5176 63130 5182 63132
rect 4936 63078 4938 63130
rect 5118 63078 5120 63130
rect 4874 63076 4880 63078
rect 4936 63076 4960 63078
rect 5016 63076 5040 63078
rect 5096 63076 5120 63078
rect 5176 63076 5182 63078
rect 4874 63067 5182 63076
rect 3424 63028 3476 63034
rect 3424 62970 3476 62976
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 1860 62484 1912 62490
rect 1860 62426 1912 62432
rect 4874 62044 5182 62053
rect 4874 62042 4880 62044
rect 4936 62042 4960 62044
rect 5016 62042 5040 62044
rect 5096 62042 5120 62044
rect 5176 62042 5182 62044
rect 4936 61990 4938 62042
rect 5118 61990 5120 62042
rect 4874 61988 4880 61990
rect 4936 61988 4960 61990
rect 5016 61988 5040 61990
rect 5096 61988 5120 61990
rect 5176 61988 5182 61990
rect 4874 61979 5182 61988
rect 1676 61872 1728 61878
rect 1676 61814 1728 61820
rect 1308 61804 1360 61810
rect 1308 61746 1360 61752
rect 1320 61305 1348 61746
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 1306 61296 1362 61305
rect 1306 61231 1362 61240
rect 4874 60956 5182 60965
rect 4874 60954 4880 60956
rect 4936 60954 4960 60956
rect 5016 60954 5040 60956
rect 5096 60954 5120 60956
rect 5176 60954 5182 60956
rect 4936 60902 4938 60954
rect 5118 60902 5120 60954
rect 4874 60900 4880 60902
rect 4936 60900 4960 60902
rect 5016 60900 5040 60902
rect 5096 60900 5120 60902
rect 5176 60900 5182 60902
rect 4874 60891 5182 60900
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 4874 59868 5182 59877
rect 4874 59866 4880 59868
rect 4936 59866 4960 59868
rect 5016 59866 5040 59868
rect 5096 59866 5120 59868
rect 5176 59866 5182 59868
rect 4936 59814 4938 59866
rect 5118 59814 5120 59866
rect 4874 59812 4880 59814
rect 4936 59812 4960 59814
rect 5016 59812 5040 59814
rect 5096 59812 5120 59814
rect 5176 59812 5182 59814
rect 4874 59803 5182 59812
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 4874 58780 5182 58789
rect 4874 58778 4880 58780
rect 4936 58778 4960 58780
rect 5016 58778 5040 58780
rect 5096 58778 5120 58780
rect 5176 58778 5182 58780
rect 4936 58726 4938 58778
rect 5118 58726 5120 58778
rect 4874 58724 4880 58726
rect 4936 58724 4960 58726
rect 5016 58724 5040 58726
rect 5096 58724 5120 58726
rect 5176 58724 5182 58726
rect 4874 58715 5182 58724
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 4874 57692 5182 57701
rect 4874 57690 4880 57692
rect 4936 57690 4960 57692
rect 5016 57690 5040 57692
rect 5096 57690 5120 57692
rect 5176 57690 5182 57692
rect 4936 57638 4938 57690
rect 5118 57638 5120 57690
rect 4874 57636 4880 57638
rect 4936 57636 4960 57638
rect 5016 57636 5040 57638
rect 5096 57636 5120 57638
rect 5176 57636 5182 57638
rect 4874 57627 5182 57636
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4874 56604 5182 56613
rect 4874 56602 4880 56604
rect 4936 56602 4960 56604
rect 5016 56602 5040 56604
rect 5096 56602 5120 56604
rect 5176 56602 5182 56604
rect 4936 56550 4938 56602
rect 5118 56550 5120 56602
rect 4874 56548 4880 56550
rect 4936 56548 4960 56550
rect 5016 56548 5040 56550
rect 5096 56548 5120 56550
rect 5176 56548 5182 56550
rect 4874 56539 5182 56548
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4874 55516 5182 55525
rect 4874 55514 4880 55516
rect 4936 55514 4960 55516
rect 5016 55514 5040 55516
rect 5096 55514 5120 55516
rect 5176 55514 5182 55516
rect 4936 55462 4938 55514
rect 5118 55462 5120 55514
rect 4874 55460 4880 55462
rect 4936 55460 4960 55462
rect 5016 55460 5040 55462
rect 5096 55460 5120 55462
rect 5176 55460 5182 55462
rect 4874 55451 5182 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4874 54428 5182 54437
rect 4874 54426 4880 54428
rect 4936 54426 4960 54428
rect 5016 54426 5040 54428
rect 5096 54426 5120 54428
rect 5176 54426 5182 54428
rect 4936 54374 4938 54426
rect 5118 54374 5120 54426
rect 4874 54372 4880 54374
rect 4936 54372 4960 54374
rect 5016 54372 5040 54374
rect 5096 54372 5120 54374
rect 5176 54372 5182 54374
rect 4874 54363 5182 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4874 53340 5182 53349
rect 4874 53338 4880 53340
rect 4936 53338 4960 53340
rect 5016 53338 5040 53340
rect 5096 53338 5120 53340
rect 5176 53338 5182 53340
rect 4936 53286 4938 53338
rect 5118 53286 5120 53338
rect 4874 53284 4880 53286
rect 4936 53284 4960 53286
rect 5016 53284 5040 53286
rect 5096 53284 5120 53286
rect 5176 53284 5182 53286
rect 4874 53275 5182 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4874 52252 5182 52261
rect 4874 52250 4880 52252
rect 4936 52250 4960 52252
rect 5016 52250 5040 52252
rect 5096 52250 5120 52252
rect 5176 52250 5182 52252
rect 4936 52198 4938 52250
rect 5118 52198 5120 52250
rect 4874 52196 4880 52198
rect 4936 52196 4960 52198
rect 5016 52196 5040 52198
rect 5096 52196 5120 52198
rect 5176 52196 5182 52198
rect 4874 52187 5182 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4874 51164 5182 51173
rect 4874 51162 4880 51164
rect 4936 51162 4960 51164
rect 5016 51162 5040 51164
rect 5096 51162 5120 51164
rect 5176 51162 5182 51164
rect 4936 51110 4938 51162
rect 5118 51110 5120 51162
rect 4874 51108 4880 51110
rect 4936 51108 4960 51110
rect 5016 51108 5040 51110
rect 5096 51108 5120 51110
rect 5176 51108 5182 51110
rect 4874 51099 5182 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4874 50076 5182 50085
rect 4874 50074 4880 50076
rect 4936 50074 4960 50076
rect 5016 50074 5040 50076
rect 5096 50074 5120 50076
rect 5176 50074 5182 50076
rect 4936 50022 4938 50074
rect 5118 50022 5120 50074
rect 4874 50020 4880 50022
rect 4936 50020 4960 50022
rect 5016 50020 5040 50022
rect 5096 50020 5120 50022
rect 5176 50020 5182 50022
rect 4874 50011 5182 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4874 48988 5182 48997
rect 4874 48986 4880 48988
rect 4936 48986 4960 48988
rect 5016 48986 5040 48988
rect 5096 48986 5120 48988
rect 5176 48986 5182 48988
rect 4936 48934 4938 48986
rect 5118 48934 5120 48986
rect 4874 48932 4880 48934
rect 4936 48932 4960 48934
rect 5016 48932 5040 48934
rect 5096 48932 5120 48934
rect 5176 48932 5182 48934
rect 4874 48923 5182 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4874 47900 5182 47909
rect 4874 47898 4880 47900
rect 4936 47898 4960 47900
rect 5016 47898 5040 47900
rect 5096 47898 5120 47900
rect 5176 47898 5182 47900
rect 4936 47846 4938 47898
rect 5118 47846 5120 47898
rect 4874 47844 4880 47846
rect 4936 47844 4960 47846
rect 5016 47844 5040 47846
rect 5096 47844 5120 47846
rect 5176 47844 5182 47846
rect 4874 47835 5182 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 5540 41744 5592 41750
rect 5540 41686 5592 41692
rect 1216 41608 1268 41614
rect 1214 41576 1216 41585
rect 1268 41576 1270 41585
rect 1214 41511 1270 41520
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 5552 41313 5580 41686
rect 5538 41304 5594 41313
rect 5538 41239 5594 41248
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 5540 40180 5592 40186
rect 5540 40122 5592 40128
rect 1400 40044 1452 40050
rect 1400 39986 1452 39992
rect 1412 39545 1440 39986
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 5552 39681 5580 40122
rect 5538 39672 5594 39681
rect 5538 39607 5594 39616
rect 1398 39536 1454 39545
rect 1398 39471 1454 39480
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 8392 38480 8444 38486
rect 8390 38448 8392 38457
rect 8444 38448 8446 38457
rect 8390 38383 8446 38392
rect 1216 38344 1268 38350
rect 1216 38286 1268 38292
rect 1228 38185 1256 38286
rect 1214 38176 1270 38185
rect 1214 38111 1270 38120
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 1400 37256 1452 37262
rect 1400 37198 1452 37204
rect 1412 36825 1440 37198
rect 9496 37188 9548 37194
rect 9496 37130 9548 37136
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 1398 36816 1454 36825
rect 1398 36751 1454 36760
rect 9508 36733 9536 37130
rect 9494 36724 9550 36733
rect 9494 36659 9550 36668
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 9496 35828 9548 35834
rect 9496 35770 9548 35776
rect 1308 35692 1360 35698
rect 9508 35650 9536 35770
rect 1308 35634 1360 35640
rect 9494 35641 9550 35650
rect 1320 35465 1348 35634
rect 9494 35576 9550 35585
rect 1306 35456 1362 35465
rect 1306 35391 1362 35400
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 5540 34740 5592 34746
rect 5540 34682 5592 34688
rect 1400 34604 1452 34610
rect 1400 34546 1452 34552
rect 1412 34105 1440 34546
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 1398 34096 1454 34105
rect 1398 34031 1454 34040
rect 5552 33969 5580 34682
rect 5538 33960 5594 33969
rect 5538 33895 5594 33904
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 1308 16108 1360 16114
rect 1308 16050 1360 16056
rect 1320 15745 1348 16050
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 1306 15736 1362 15745
rect 4214 15739 4522 15748
rect 1306 15671 1362 15680
rect 9508 15490 9536 15914
rect 9494 15481 9550 15490
rect 9494 15416 9550 15425
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 9600 9897 9628 66234
rect 10336 64326 10364 67730
rect 29000 67720 29052 67726
rect 16394 67688 16450 67697
rect 29000 67662 29052 67668
rect 16394 67623 16396 67632
rect 16448 67623 16450 67632
rect 22100 67652 22152 67658
rect 16396 67594 16448 67600
rect 22100 67594 22152 67600
rect 16408 66314 16436 67594
rect 18880 67380 18932 67386
rect 18880 67322 18932 67328
rect 17316 67244 17368 67250
rect 17316 67186 17368 67192
rect 17328 66706 17356 67186
rect 18892 66774 18920 67322
rect 20352 67176 20404 67182
rect 22112 67130 22140 67594
rect 22376 67584 22428 67590
rect 22376 67526 22428 67532
rect 20352 67118 20404 67124
rect 20260 67040 20312 67046
rect 19338 67008 19394 67017
rect 20260 66982 20312 66988
rect 19338 66943 19394 66952
rect 18880 66768 18932 66774
rect 18880 66710 18932 66716
rect 19352 66706 19380 66943
rect 17316 66700 17368 66706
rect 17316 66642 17368 66648
rect 19340 66700 19392 66706
rect 19340 66642 19392 66648
rect 20272 66502 20300 66982
rect 20364 66881 20392 67118
rect 21836 67102 22140 67130
rect 21272 67040 21324 67046
rect 21272 66982 21324 66988
rect 20350 66872 20406 66881
rect 20350 66807 20406 66816
rect 20260 66496 20312 66502
rect 20260 66438 20312 66444
rect 20444 66496 20496 66502
rect 20444 66438 20496 66444
rect 16408 66298 16528 66314
rect 16396 66292 16528 66298
rect 16448 66286 16528 66292
rect 16396 66234 16448 66240
rect 16500 66144 16528 66286
rect 20272 66162 20300 66438
rect 20456 66298 20484 66438
rect 20444 66292 20496 66298
rect 20444 66234 20496 66240
rect 21284 66162 21312 66982
rect 21836 66570 21864 67102
rect 22008 67040 22060 67046
rect 22008 66982 22060 66988
rect 22020 66570 22048 66982
rect 22388 66638 22416 67526
rect 24676 67380 24728 67386
rect 24676 67322 24728 67328
rect 24308 67312 24360 67318
rect 24308 67254 24360 67260
rect 23296 67040 23348 67046
rect 23296 66982 23348 66988
rect 23308 66842 23336 66982
rect 24320 66842 24348 67254
rect 23296 66836 23348 66842
rect 23296 66778 23348 66784
rect 24308 66836 24360 66842
rect 24308 66778 24360 66784
rect 22376 66632 22428 66638
rect 22376 66574 22428 66580
rect 24688 66570 24716 67322
rect 29012 67250 29040 67662
rect 31024 67584 31076 67590
rect 31024 67526 31076 67532
rect 32864 67584 32916 67590
rect 32864 67526 32916 67532
rect 29000 67244 29052 67250
rect 29000 67186 29052 67192
rect 25044 67176 25096 67182
rect 25044 67118 25096 67124
rect 25056 66706 25084 67118
rect 25780 67040 25832 67046
rect 29012 67017 29040 67186
rect 29092 67176 29144 67182
rect 29092 67118 29144 67124
rect 25780 66982 25832 66988
rect 28998 67008 29054 67017
rect 25044 66700 25096 66706
rect 25044 66642 25096 66648
rect 25792 66638 25820 66982
rect 28998 66943 29054 66952
rect 27066 66872 27122 66881
rect 27066 66807 27122 66816
rect 27080 66774 27108 66807
rect 27068 66768 27120 66774
rect 27068 66710 27120 66716
rect 29012 66638 29040 66943
rect 29104 66774 29132 67118
rect 31036 67046 31064 67526
rect 31208 67244 31260 67250
rect 31208 67186 31260 67192
rect 32772 67244 32824 67250
rect 32772 67186 32824 67192
rect 30564 67040 30616 67046
rect 30564 66982 30616 66988
rect 31024 67040 31076 67046
rect 31024 66982 31076 66988
rect 29734 66872 29790 66881
rect 29734 66807 29736 66816
rect 29788 66807 29790 66816
rect 29736 66778 29788 66784
rect 29092 66768 29144 66774
rect 29092 66710 29144 66716
rect 25780 66632 25832 66638
rect 25780 66574 25832 66580
rect 29000 66632 29052 66638
rect 29000 66574 29052 66580
rect 21824 66564 21876 66570
rect 21824 66506 21876 66512
rect 22008 66564 22060 66570
rect 22008 66506 22060 66512
rect 24676 66564 24728 66570
rect 24676 66506 24728 66512
rect 22020 66230 22048 66506
rect 26148 66496 26200 66502
rect 26148 66438 26200 66444
rect 22008 66224 22060 66230
rect 23756 66224 23808 66230
rect 22008 66166 22060 66172
rect 23584 66172 23756 66178
rect 23584 66166 23808 66172
rect 23584 66162 23796 66166
rect 16580 66156 16632 66162
rect 16500 66116 16580 66144
rect 16580 66098 16632 66104
rect 20260 66156 20312 66162
rect 20260 66098 20312 66104
rect 21272 66156 21324 66162
rect 21272 66098 21324 66104
rect 23572 66156 23796 66162
rect 23624 66150 23796 66156
rect 23572 66098 23624 66104
rect 22376 66088 22428 66094
rect 22020 66036 22376 66042
rect 22020 66030 22428 66036
rect 22020 66014 22416 66030
rect 22020 64462 22048 66014
rect 26160 64938 26188 66438
rect 29104 66298 29132 66710
rect 30104 66496 30156 66502
rect 30104 66438 30156 66444
rect 30116 66298 30144 66438
rect 29092 66292 29144 66298
rect 29092 66234 29144 66240
rect 30104 66292 30156 66298
rect 30104 66234 30156 66240
rect 30116 65550 30144 66234
rect 30576 66230 30604 66982
rect 31024 66564 31076 66570
rect 31024 66506 31076 66512
rect 31036 66230 31064 66506
rect 31220 66230 31248 67186
rect 32784 66774 32812 67186
rect 32876 67114 32904 67526
rect 33508 67244 33560 67250
rect 33508 67186 33560 67192
rect 32956 67176 33008 67182
rect 32956 67118 33008 67124
rect 32864 67108 32916 67114
rect 32864 67050 32916 67056
rect 32772 66768 32824 66774
rect 32772 66710 32824 66716
rect 31944 66496 31996 66502
rect 31944 66438 31996 66444
rect 32772 66496 32824 66502
rect 32772 66438 32824 66444
rect 31956 66298 31984 66438
rect 31944 66292 31996 66298
rect 31944 66234 31996 66240
rect 30564 66224 30616 66230
rect 30564 66166 30616 66172
rect 31024 66224 31076 66230
rect 31024 66166 31076 66172
rect 31208 66224 31260 66230
rect 31208 66166 31260 66172
rect 32784 66094 32812 66438
rect 32968 66298 32996 67118
rect 33520 67046 33548 67186
rect 33508 67040 33560 67046
rect 33508 66982 33560 66988
rect 33048 66768 33100 66774
rect 33048 66710 33100 66716
rect 33060 66638 33088 66710
rect 33048 66632 33100 66638
rect 33046 66600 33048 66609
rect 33100 66600 33102 66609
rect 33046 66535 33102 66544
rect 32956 66292 33008 66298
rect 32956 66234 33008 66240
rect 32772 66088 32824 66094
rect 32772 66030 32824 66036
rect 30104 65544 30156 65550
rect 33520 65521 33548 66982
rect 33612 66706 33640 68410
rect 33692 68400 33744 68406
rect 33692 68342 33744 68348
rect 33704 67250 33732 68342
rect 33980 67930 34008 69527
rect 35176 69426 35204 69527
rect 36372 69494 36400 69527
rect 36360 69488 36412 69494
rect 36360 69430 36412 69436
rect 35164 69420 35216 69426
rect 35164 69362 35216 69368
rect 35176 67930 35204 69362
rect 35992 68332 36044 68338
rect 35992 68274 36044 68280
rect 33968 67924 34020 67930
rect 33968 67866 34020 67872
rect 35164 67924 35216 67930
rect 35164 67866 35216 67872
rect 35594 67484 35902 67493
rect 35594 67482 35600 67484
rect 35656 67482 35680 67484
rect 35736 67482 35760 67484
rect 35816 67482 35840 67484
rect 35896 67482 35902 67484
rect 35656 67430 35658 67482
rect 35838 67430 35840 67482
rect 35594 67428 35600 67430
rect 35656 67428 35680 67430
rect 35736 67428 35760 67430
rect 35816 67428 35840 67430
rect 35896 67428 35902 67430
rect 35594 67419 35902 67428
rect 36004 67386 36032 68274
rect 36372 67930 36400 69430
rect 37476 67930 37504 69702
rect 38672 67930 38700 69799
rect 39816 69799 39818 69808
rect 40958 69864 40960 69873
rect 43272 69873 43300 69906
rect 70952 69896 71004 69902
rect 41012 69864 41014 69873
rect 40958 69799 41014 69808
rect 43258 69864 43314 69873
rect 70952 69838 71004 69844
rect 43258 69799 43314 69808
rect 69296 69828 69348 69834
rect 39764 69770 39816 69776
rect 39776 67930 39804 69770
rect 40972 67930 41000 69799
rect 42154 69592 42210 69601
rect 42154 69527 42210 69536
rect 42168 68678 42196 69527
rect 42156 68672 42208 68678
rect 42156 68614 42208 68620
rect 42168 67930 42196 68614
rect 43272 67930 43300 69799
rect 69296 69770 69348 69776
rect 68468 69760 68520 69766
rect 68468 69702 68520 69708
rect 66996 69692 67048 69698
rect 66996 69634 67048 69640
rect 65654 68028 65962 68037
rect 65654 68026 65660 68028
rect 65716 68026 65740 68028
rect 65796 68026 65820 68028
rect 65876 68026 65900 68028
rect 65956 68026 65962 68028
rect 65716 67974 65718 68026
rect 65898 67974 65900 68026
rect 65654 67972 65660 67974
rect 65716 67972 65740 67974
rect 65796 67972 65820 67974
rect 65876 67972 65900 67974
rect 65956 67972 65962 67974
rect 65654 67963 65962 67972
rect 36360 67924 36412 67930
rect 36360 67866 36412 67872
rect 37464 67924 37516 67930
rect 37464 67866 37516 67872
rect 38660 67924 38712 67930
rect 38660 67866 38712 67872
rect 39764 67924 39816 67930
rect 39764 67866 39816 67872
rect 40960 67924 41012 67930
rect 40960 67866 41012 67872
rect 42156 67924 42208 67930
rect 42156 67866 42208 67872
rect 43260 67924 43312 67930
rect 43260 67866 43312 67872
rect 38660 67584 38712 67590
rect 38660 67526 38712 67532
rect 40406 67552 40462 67561
rect 38672 67386 38700 67526
rect 40406 67487 40462 67496
rect 35348 67380 35400 67386
rect 35348 67322 35400 67328
rect 35992 67380 36044 67386
rect 35992 67322 36044 67328
rect 38660 67380 38712 67386
rect 38660 67322 38712 67328
rect 39948 67380 40000 67386
rect 39948 67322 40000 67328
rect 33692 67244 33744 67250
rect 33692 67186 33744 67192
rect 34244 67176 34296 67182
rect 34244 67118 34296 67124
rect 34256 66774 34284 67118
rect 34934 66940 35242 66949
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66875 35242 66884
rect 34244 66768 34296 66774
rect 34244 66710 34296 66716
rect 33600 66700 33652 66706
rect 33600 66642 33652 66648
rect 33876 66700 33928 66706
rect 33876 66642 33928 66648
rect 33612 66502 33640 66642
rect 33888 66609 33916 66642
rect 35360 66609 35388 67322
rect 39028 67244 39080 67250
rect 39028 67186 39080 67192
rect 35992 66632 36044 66638
rect 33874 66600 33930 66609
rect 33874 66535 33930 66544
rect 35346 66600 35402 66609
rect 35992 66574 36044 66580
rect 35346 66535 35402 66544
rect 33600 66496 33652 66502
rect 33600 66438 33652 66444
rect 35594 66396 35902 66405
rect 35594 66394 35600 66396
rect 35656 66394 35680 66396
rect 35736 66394 35760 66396
rect 35816 66394 35840 66396
rect 35896 66394 35902 66396
rect 35656 66342 35658 66394
rect 35838 66342 35840 66394
rect 35594 66340 35600 66342
rect 35656 66340 35680 66342
rect 35736 66340 35760 66342
rect 35816 66340 35840 66342
rect 35896 66340 35902 66342
rect 35594 66331 35902 66340
rect 34934 65852 35242 65861
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65787 35242 65796
rect 30104 65486 30156 65492
rect 33506 65512 33562 65521
rect 33506 65447 33562 65456
rect 26148 64932 26200 64938
rect 26148 64874 26200 64880
rect 22008 64456 22060 64462
rect 22008 64398 22060 64404
rect 10324 64320 10376 64326
rect 10324 64262 10376 64268
rect 36004 64161 36032 66574
rect 39040 66337 39068 67186
rect 39120 67176 39172 67182
rect 39120 67118 39172 67124
rect 39132 66745 39160 67118
rect 39396 67108 39448 67114
rect 39396 67050 39448 67056
rect 39118 66736 39174 66745
rect 39118 66671 39174 66680
rect 39026 66328 39082 66337
rect 39408 66298 39436 67050
rect 39960 67046 39988 67322
rect 40420 67182 40448 67487
rect 66314 67484 66622 67493
rect 66314 67482 66320 67484
rect 66376 67482 66400 67484
rect 66456 67482 66480 67484
rect 66536 67482 66560 67484
rect 66616 67482 66622 67484
rect 66376 67430 66378 67482
rect 66558 67430 66560 67482
rect 66314 67428 66320 67430
rect 66376 67428 66400 67430
rect 66456 67428 66480 67430
rect 66536 67428 66560 67430
rect 66616 67428 66622 67430
rect 66314 67419 66622 67428
rect 67008 67386 67036 69634
rect 68284 67584 68336 67590
rect 68284 67526 68336 67532
rect 47860 67380 47912 67386
rect 47860 67322 47912 67328
rect 66996 67380 67048 67386
rect 66996 67322 67048 67328
rect 45744 67312 45796 67318
rect 46664 67312 46716 67318
rect 45744 67254 45796 67260
rect 46662 67280 46664 67289
rect 46716 67280 46718 67289
rect 40408 67176 40460 67182
rect 44456 67176 44508 67182
rect 40408 67118 40460 67124
rect 44454 67144 44456 67153
rect 44508 67144 44510 67153
rect 40420 67046 40448 67118
rect 44454 67079 44510 67088
rect 39948 67040 40000 67046
rect 39948 66982 40000 66988
rect 40408 67040 40460 67046
rect 40408 66982 40460 66988
rect 43996 67040 44048 67046
rect 43996 66982 44048 66988
rect 44008 66842 44036 66982
rect 43996 66836 44048 66842
rect 43996 66778 44048 66784
rect 39026 66263 39082 66272
rect 39396 66292 39448 66298
rect 39396 66234 39448 66240
rect 45756 66201 45784 67254
rect 46662 67215 46718 67224
rect 47492 67244 47544 67250
rect 47492 67186 47544 67192
rect 45742 66192 45798 66201
rect 45742 66127 45798 66136
rect 47504 64161 47532 67186
rect 47872 66609 47900 67322
rect 62394 67280 62450 67289
rect 62394 67215 62396 67224
rect 62448 67215 62450 67224
rect 62396 67186 62448 67192
rect 68296 67182 68324 67526
rect 68480 67318 68508 69702
rect 69018 67552 69074 67561
rect 69018 67487 69074 67496
rect 69032 67386 69060 67487
rect 69020 67380 69072 67386
rect 69020 67322 69072 67328
rect 68468 67312 68520 67318
rect 68468 67254 68520 67260
rect 68560 67244 68612 67250
rect 68560 67186 68612 67192
rect 68284 67176 68336 67182
rect 62210 67144 62266 67153
rect 60740 67108 60792 67114
rect 68284 67118 68336 67124
rect 62210 67079 62212 67088
rect 60740 67050 60792 67056
rect 62264 67079 62266 67088
rect 63408 67108 63460 67114
rect 62212 67050 62264 67056
rect 63408 67050 63460 67056
rect 67548 67108 67600 67114
rect 67548 67050 67600 67056
rect 53656 66768 53708 66774
rect 53656 66710 53708 66716
rect 47858 66600 47914 66609
rect 47858 66535 47914 66544
rect 53668 65958 53696 66710
rect 57888 66496 57940 66502
rect 57888 66438 57940 66444
rect 57900 66230 57928 66438
rect 57888 66224 57940 66230
rect 57888 66166 57940 66172
rect 60752 66162 60780 67050
rect 60740 66156 60792 66162
rect 60740 66098 60792 66104
rect 53656 65952 53708 65958
rect 53654 65920 53656 65929
rect 53708 65920 53710 65929
rect 53654 65855 53710 65864
rect 63420 64161 63448 67050
rect 66168 67040 66220 67046
rect 66168 66982 66220 66988
rect 65654 66940 65962 66949
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66875 65962 66884
rect 65654 65852 65962 65861
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65787 65962 65796
rect 35990 64152 36046 64161
rect 35990 64087 36046 64096
rect 47490 64152 47546 64161
rect 47490 64087 47546 64096
rect 63406 64152 63462 64161
rect 63406 64087 63462 64096
rect 66180 64025 66208 66982
rect 67560 66745 67588 67050
rect 67546 66736 67602 66745
rect 68296 66706 68324 67118
rect 68572 66842 68600 67186
rect 68560 66836 68612 66842
rect 68560 66778 68612 66784
rect 67546 66671 67602 66680
rect 68284 66700 68336 66706
rect 68284 66642 68336 66648
rect 67638 66600 67694 66609
rect 67638 66535 67640 66544
rect 67692 66535 67694 66544
rect 67640 66506 67692 66512
rect 69308 66502 69336 69770
rect 69754 68232 69810 68241
rect 69754 68167 69810 68176
rect 69768 67930 69796 68167
rect 69756 67924 69808 67930
rect 69756 67866 69808 67872
rect 69664 67584 69716 67590
rect 69664 67526 69716 67532
rect 69676 67266 69704 67526
rect 69768 67386 69796 67866
rect 69848 67584 69900 67590
rect 69848 67526 69900 67532
rect 69756 67380 69808 67386
rect 69756 67322 69808 67328
rect 69480 67244 69532 67250
rect 69676 67238 69796 67266
rect 69480 67186 69532 67192
rect 69492 67046 69520 67186
rect 69768 67182 69796 67238
rect 69756 67176 69808 67182
rect 69756 67118 69808 67124
rect 69480 67040 69532 67046
rect 69480 66982 69532 66988
rect 69860 66502 69888 67526
rect 70964 67386 70992 69838
rect 70952 67380 71004 67386
rect 70952 67322 71004 67328
rect 69940 67176 69992 67182
rect 69940 67118 69992 67124
rect 70032 67176 70084 67182
rect 70032 67118 70084 67124
rect 69952 66570 69980 67118
rect 70044 66706 70072 67118
rect 70400 67108 70452 67114
rect 70400 67050 70452 67056
rect 70584 67108 70636 67114
rect 70584 67050 70636 67056
rect 70412 67017 70440 67050
rect 70398 67008 70454 67017
rect 70398 66943 70454 66952
rect 70032 66700 70084 66706
rect 70032 66642 70084 66648
rect 70596 66638 70624 67050
rect 70964 66774 70992 67322
rect 71792 67250 71820 69906
rect 73632 67250 73660 69974
rect 90362 69864 90418 69873
rect 90362 69799 90418 69808
rect 88616 68808 88668 68814
rect 88616 68750 88668 68756
rect 88340 68400 88392 68406
rect 88340 68342 88392 68348
rect 88352 67930 88380 68342
rect 88340 67924 88392 67930
rect 88340 67866 88392 67872
rect 85672 67720 85724 67726
rect 85672 67662 85724 67668
rect 87512 67720 87564 67726
rect 87512 67662 87564 67668
rect 79966 67552 80022 67561
rect 79966 67487 80022 67496
rect 75366 67416 75422 67425
rect 73988 67380 74040 67386
rect 75366 67351 75368 67360
rect 73988 67322 74040 67328
rect 75420 67351 75422 67360
rect 75460 67380 75512 67386
rect 75368 67322 75420 67328
rect 75460 67322 75512 67328
rect 75828 67380 75880 67386
rect 75828 67322 75880 67328
rect 71780 67244 71832 67250
rect 71780 67186 71832 67192
rect 71872 67244 71924 67250
rect 71872 67186 71924 67192
rect 73620 67244 73672 67250
rect 73620 67186 73672 67192
rect 73712 67244 73764 67250
rect 73712 67186 73764 67192
rect 71792 66774 71820 67186
rect 70952 66768 71004 66774
rect 70952 66710 71004 66716
rect 71780 66768 71832 66774
rect 71780 66710 71832 66716
rect 70308 66632 70360 66638
rect 70308 66574 70360 66580
rect 70584 66632 70636 66638
rect 70584 66574 70636 66580
rect 69940 66564 69992 66570
rect 69940 66506 69992 66512
rect 69296 66496 69348 66502
rect 69296 66438 69348 66444
rect 69848 66496 69900 66502
rect 69848 66438 69900 66444
rect 66314 66396 66622 66405
rect 66314 66394 66320 66396
rect 66376 66394 66400 66396
rect 66456 66394 66480 66396
rect 66536 66394 66560 66396
rect 66616 66394 66622 66396
rect 66376 66342 66378 66394
rect 66558 66342 66560 66394
rect 66314 66340 66320 66342
rect 66376 66340 66400 66342
rect 66456 66340 66480 66342
rect 66536 66340 66560 66342
rect 66616 66340 66622 66342
rect 66314 66331 66622 66340
rect 70320 66298 70348 66574
rect 70308 66292 70360 66298
rect 70308 66234 70360 66240
rect 66166 64016 66222 64025
rect 66166 63951 66222 63960
rect 71884 63889 71912 67186
rect 73724 66337 73752 67186
rect 73710 66328 73766 66337
rect 73710 66263 73766 66272
rect 74000 66094 74028 67322
rect 73988 66088 74040 66094
rect 73988 66030 74040 66036
rect 75472 64161 75500 67322
rect 75644 67244 75696 67250
rect 75644 67186 75696 67192
rect 75656 67046 75684 67186
rect 75644 67040 75696 67046
rect 75644 66982 75696 66988
rect 75840 66842 75868 67322
rect 76196 67244 76248 67250
rect 76196 67186 76248 67192
rect 77392 67244 77444 67250
rect 77392 67186 77444 67192
rect 77576 67244 77628 67250
rect 77576 67186 77628 67192
rect 75828 66836 75880 66842
rect 75828 66778 75880 66784
rect 76208 66706 76236 67186
rect 76196 66700 76248 66706
rect 76196 66642 76248 66648
rect 75920 66632 75972 66638
rect 75920 66574 75972 66580
rect 75932 65618 75960 66574
rect 75920 65612 75972 65618
rect 75920 65554 75972 65560
rect 77404 64190 77432 67186
rect 77588 66502 77616 67186
rect 77944 67108 77996 67114
rect 77944 67050 77996 67056
rect 77956 66638 77984 67050
rect 79784 67040 79836 67046
rect 79784 66982 79836 66988
rect 79876 67040 79928 67046
rect 79876 66982 79928 66988
rect 79796 66638 79824 66982
rect 79888 66842 79916 66982
rect 79980 66858 80008 67487
rect 85212 67176 85264 67182
rect 85212 67118 85264 67124
rect 85580 67176 85632 67182
rect 85580 67118 85632 67124
rect 83096 67040 83148 67046
rect 85224 67028 85252 67118
rect 85224 67000 85344 67028
rect 85592 67017 85620 67118
rect 83096 66982 83148 66988
rect 79980 66842 80192 66858
rect 83108 66842 83136 66982
rect 79876 66836 79928 66842
rect 79980 66836 80204 66842
rect 79980 66830 80152 66836
rect 79876 66778 79928 66784
rect 80152 66778 80204 66784
rect 83096 66836 83148 66842
rect 83096 66778 83148 66784
rect 84842 66736 84898 66745
rect 79968 66700 80020 66706
rect 79968 66642 80020 66648
rect 83372 66700 83424 66706
rect 84842 66671 84844 66680
rect 83372 66642 83424 66648
rect 84896 66671 84898 66680
rect 84844 66642 84896 66648
rect 77944 66632 77996 66638
rect 77944 66574 77996 66580
rect 79784 66632 79836 66638
rect 79784 66574 79836 66580
rect 77576 66496 77628 66502
rect 77576 66438 77628 66444
rect 79980 66450 80008 66642
rect 80152 66496 80204 66502
rect 79980 66444 80152 66450
rect 79980 66438 80204 66444
rect 77588 66298 77616 66438
rect 79980 66422 80192 66438
rect 80164 66298 80192 66422
rect 77576 66292 77628 66298
rect 77576 66234 77628 66240
rect 80152 66292 80204 66298
rect 80152 66234 80204 66240
rect 83384 66230 83412 66642
rect 84660 66632 84712 66638
rect 84658 66600 84660 66609
rect 84712 66600 84714 66609
rect 85316 66570 85344 67000
rect 85578 67008 85634 67017
rect 85578 66943 85634 66952
rect 85684 66774 85712 67662
rect 86224 67652 86276 67658
rect 86224 67594 86276 67600
rect 86236 67046 86264 67594
rect 87524 67250 87552 67662
rect 88628 67250 88656 68750
rect 89168 68264 89220 68270
rect 89168 68206 89220 68212
rect 88892 68128 88944 68134
rect 88892 68070 88944 68076
rect 88904 67930 88932 68070
rect 89180 67930 89208 68206
rect 88892 67924 88944 67930
rect 88892 67866 88944 67872
rect 89168 67924 89220 67930
rect 89168 67866 89220 67872
rect 90376 67794 90404 69799
rect 96894 69592 96950 69601
rect 96894 69527 96950 69536
rect 90822 68776 90878 68785
rect 90822 68711 90878 68720
rect 95884 68740 95936 68746
rect 90640 68332 90692 68338
rect 90640 68274 90692 68280
rect 90364 67788 90416 67794
rect 90364 67730 90416 67736
rect 89076 67720 89128 67726
rect 89076 67662 89128 67668
rect 86960 67244 87012 67250
rect 86960 67186 87012 67192
rect 87512 67244 87564 67250
rect 87512 67186 87564 67192
rect 88524 67244 88576 67250
rect 88524 67186 88576 67192
rect 88616 67244 88668 67250
rect 88616 67186 88668 67192
rect 86224 67040 86276 67046
rect 86224 66982 86276 66988
rect 85672 66768 85724 66774
rect 85394 66736 85450 66745
rect 85672 66710 85724 66716
rect 86236 66706 86264 66982
rect 85394 66671 85396 66680
rect 85448 66671 85450 66680
rect 86224 66700 86276 66706
rect 85396 66642 85448 66648
rect 86224 66642 86276 66648
rect 84658 66535 84714 66544
rect 85304 66564 85356 66570
rect 85304 66506 85356 66512
rect 84936 66496 84988 66502
rect 84936 66438 84988 66444
rect 83372 66224 83424 66230
rect 83372 66166 83424 66172
rect 84948 65521 84976 66438
rect 86236 66094 86264 66642
rect 86972 66450 87000 67186
rect 88432 67108 88484 67114
rect 88432 67050 88484 67056
rect 87604 67040 87656 67046
rect 87604 66982 87656 66988
rect 87788 67040 87840 67046
rect 87788 66982 87840 66988
rect 86512 66422 87000 66450
rect 86512 66162 86540 66422
rect 86960 66292 87012 66298
rect 86960 66234 87012 66240
rect 86500 66156 86552 66162
rect 86500 66098 86552 66104
rect 86224 66088 86276 66094
rect 86224 66030 86276 66036
rect 86592 66020 86644 66026
rect 86592 65962 86644 65968
rect 85580 65952 85632 65958
rect 85580 65894 85632 65900
rect 86500 65952 86552 65958
rect 86500 65894 86552 65900
rect 86604 65906 86632 65962
rect 86776 65952 86828 65958
rect 86604 65900 86776 65906
rect 86604 65894 86828 65900
rect 84934 65512 84990 65521
rect 85592 65482 85620 65894
rect 86512 65618 86540 65894
rect 86604 65878 86816 65894
rect 86972 65754 87000 66234
rect 86960 65748 87012 65754
rect 86960 65690 87012 65696
rect 86500 65612 86552 65618
rect 86500 65554 86552 65560
rect 84934 65447 84990 65456
rect 85580 65476 85632 65482
rect 85580 65418 85632 65424
rect 87616 65074 87644 66982
rect 87800 65686 87828 66982
rect 88340 66836 88392 66842
rect 88340 66778 88392 66784
rect 88352 66722 88380 66778
rect 87892 66694 88380 66722
rect 88444 66706 88472 67050
rect 88432 66700 88484 66706
rect 87892 66502 87920 66694
rect 88432 66642 88484 66648
rect 88340 66564 88392 66570
rect 88340 66506 88392 66512
rect 87880 66496 87932 66502
rect 87972 66496 88024 66502
rect 87880 66438 87932 66444
rect 87970 66464 87972 66473
rect 88024 66464 88026 66473
rect 87970 66399 88026 66408
rect 88352 66298 88380 66506
rect 88444 66298 88472 66642
rect 88536 66473 88564 67186
rect 88522 66464 88578 66473
rect 88522 66399 88578 66408
rect 88340 66292 88392 66298
rect 88340 66234 88392 66240
rect 88432 66292 88484 66298
rect 88432 66234 88484 66240
rect 88064 66156 88116 66162
rect 88064 66098 88116 66104
rect 88432 66156 88484 66162
rect 88432 66098 88484 66104
rect 87788 65680 87840 65686
rect 87788 65622 87840 65628
rect 88076 65618 88104 66098
rect 88444 65958 88472 66098
rect 88432 65952 88484 65958
rect 88432 65894 88484 65900
rect 88064 65612 88116 65618
rect 88064 65554 88116 65560
rect 87604 65068 87656 65074
rect 87604 65010 87656 65016
rect 88536 64462 88564 66399
rect 88628 66162 88656 67186
rect 89088 66620 89116 67662
rect 89812 67652 89864 67658
rect 89812 67594 89864 67600
rect 89260 67584 89312 67590
rect 89260 67526 89312 67532
rect 89272 67250 89300 67526
rect 89352 67380 89404 67386
rect 89352 67322 89404 67328
rect 89260 67244 89312 67250
rect 89260 67186 89312 67192
rect 89364 67046 89392 67322
rect 89536 67244 89588 67250
rect 89536 67186 89588 67192
rect 89352 67040 89404 67046
rect 89352 66982 89404 66988
rect 89548 66722 89576 67186
rect 89824 67114 89852 67594
rect 90652 67590 90680 68274
rect 90732 68196 90784 68202
rect 90732 68138 90784 68144
rect 90744 67930 90772 68138
rect 90836 67930 90864 68711
rect 95884 68682 95936 68688
rect 93584 68400 93636 68406
rect 93584 68342 93636 68348
rect 91560 68196 91612 68202
rect 91560 68138 91612 68144
rect 90732 67924 90784 67930
rect 90732 67866 90784 67872
rect 90824 67924 90876 67930
rect 90824 67866 90876 67872
rect 90916 67856 90968 67862
rect 90916 67798 90968 67804
rect 91008 67856 91060 67862
rect 91008 67798 91060 67804
rect 90928 67697 90956 67798
rect 90914 67688 90970 67697
rect 90914 67623 90970 67632
rect 90640 67584 90692 67590
rect 90824 67584 90876 67590
rect 90640 67526 90692 67532
rect 90822 67552 90824 67561
rect 90916 67584 90968 67590
rect 90876 67552 90878 67561
rect 90916 67526 90968 67532
rect 90822 67487 90878 67496
rect 89812 67108 89864 67114
rect 89812 67050 89864 67056
rect 89548 66694 89760 66722
rect 89628 66632 89680 66638
rect 89088 66592 89628 66620
rect 89088 66162 89116 66592
rect 89628 66574 89680 66580
rect 89732 66450 89760 66694
rect 90928 66502 90956 67526
rect 89640 66422 89760 66450
rect 90272 66496 90324 66502
rect 90272 66438 90324 66444
rect 90916 66496 90968 66502
rect 90916 66438 90968 66444
rect 89640 66298 89668 66422
rect 89628 66292 89680 66298
rect 89628 66234 89680 66240
rect 89812 66224 89864 66230
rect 89732 66184 89812 66212
rect 89732 66178 89760 66184
rect 88616 66156 88668 66162
rect 88616 66098 88668 66104
rect 89076 66156 89128 66162
rect 89076 66098 89128 66104
rect 89640 66150 89760 66178
rect 89812 66166 89864 66172
rect 89640 65686 89668 66150
rect 90284 65958 90312 66438
rect 90928 66094 90956 66438
rect 91020 66337 91048 67798
rect 91468 67720 91520 67726
rect 91572 67674 91600 68138
rect 93492 68128 93544 68134
rect 93492 68070 93544 68076
rect 91520 67668 91600 67674
rect 91468 67662 91600 67668
rect 93400 67720 93452 67726
rect 93400 67662 93452 67668
rect 91480 67646 91600 67662
rect 91572 67318 91600 67646
rect 91744 67652 91796 67658
rect 91744 67594 91796 67600
rect 92664 67652 92716 67658
rect 92664 67594 92716 67600
rect 91560 67312 91612 67318
rect 91560 67254 91612 67260
rect 91006 66328 91062 66337
rect 91006 66263 91062 66272
rect 90916 66088 90968 66094
rect 90916 66030 90968 66036
rect 90272 65952 90324 65958
rect 90272 65894 90324 65900
rect 91192 65952 91244 65958
rect 91192 65894 91244 65900
rect 91204 65686 91232 65894
rect 89628 65680 89680 65686
rect 89628 65622 89680 65628
rect 91192 65680 91244 65686
rect 91192 65622 91244 65628
rect 91756 65618 91784 67594
rect 92112 67380 92164 67386
rect 92112 67322 92164 67328
rect 92020 67244 92072 67250
rect 92124 67232 92152 67322
rect 92072 67204 92152 67232
rect 92020 67186 92072 67192
rect 92296 67176 92348 67182
rect 92296 67118 92348 67124
rect 92020 67040 92072 67046
rect 92020 66982 92072 66988
rect 92032 66842 92060 66982
rect 92020 66836 92072 66842
rect 92020 66778 92072 66784
rect 92308 66094 92336 67118
rect 92676 66162 92704 67594
rect 93308 67380 93360 67386
rect 93308 67322 93360 67328
rect 93216 66632 93268 66638
rect 93320 66620 93348 67322
rect 93412 67114 93440 67662
rect 93504 67164 93532 68070
rect 93596 67318 93624 68342
rect 95700 68332 95752 68338
rect 95700 68274 95752 68280
rect 94044 68264 94096 68270
rect 94044 68206 94096 68212
rect 93952 67652 94004 67658
rect 93952 67594 94004 67600
rect 93676 67584 93728 67590
rect 93676 67526 93728 67532
rect 93768 67584 93820 67590
rect 93768 67526 93820 67532
rect 93584 67312 93636 67318
rect 93584 67254 93636 67260
rect 93504 67136 93624 67164
rect 93400 67108 93452 67114
rect 93400 67050 93452 67056
rect 93268 66592 93348 66620
rect 93216 66574 93268 66580
rect 93032 66496 93084 66502
rect 93032 66438 93084 66444
rect 93044 66230 93072 66438
rect 93320 66298 93348 66592
rect 93596 66570 93624 67136
rect 93688 67046 93716 67526
rect 93780 67182 93808 67526
rect 93768 67176 93820 67182
rect 93768 67118 93820 67124
rect 93676 67040 93728 67046
rect 93676 66982 93728 66988
rect 93492 66564 93544 66570
rect 93492 66506 93544 66512
rect 93584 66564 93636 66570
rect 93584 66506 93636 66512
rect 93308 66292 93360 66298
rect 93308 66234 93360 66240
rect 92940 66224 92992 66230
rect 92940 66166 92992 66172
rect 93032 66224 93084 66230
rect 93032 66166 93084 66172
rect 92664 66156 92716 66162
rect 92664 66098 92716 66104
rect 92296 66088 92348 66094
rect 92296 66030 92348 66036
rect 92952 66042 92980 66166
rect 93504 66094 93532 66506
rect 93964 66162 93992 67594
rect 94056 66706 94084 68206
rect 95608 68128 95660 68134
rect 95608 68070 95660 68076
rect 94136 67924 94188 67930
rect 94136 67866 94188 67872
rect 95056 67924 95108 67930
rect 95056 67866 95108 67872
rect 94148 67726 94176 67866
rect 94964 67856 95016 67862
rect 94964 67798 95016 67804
rect 94136 67720 94188 67726
rect 94136 67662 94188 67668
rect 94778 67552 94834 67561
rect 94778 67487 94834 67496
rect 94792 67182 94820 67487
rect 94504 67176 94556 67182
rect 94504 67118 94556 67124
rect 94780 67176 94832 67182
rect 94780 67118 94832 67124
rect 94516 66842 94544 67118
rect 94976 66842 95004 67798
rect 95068 67726 95096 67866
rect 95620 67833 95648 68070
rect 95606 67824 95662 67833
rect 95606 67759 95662 67768
rect 95620 67726 95648 67759
rect 95056 67720 95108 67726
rect 95332 67720 95384 67726
rect 95056 67662 95108 67668
rect 95330 67688 95332 67697
rect 95608 67720 95660 67726
rect 95384 67688 95386 67697
rect 95608 67662 95660 67668
rect 95330 67623 95386 67632
rect 95712 67590 95740 68274
rect 95700 67584 95752 67590
rect 95792 67584 95844 67590
rect 95700 67526 95752 67532
rect 95790 67552 95792 67561
rect 95844 67552 95846 67561
rect 94504 66836 94556 66842
rect 94504 66778 94556 66784
rect 94964 66836 95016 66842
rect 94964 66778 95016 66784
rect 94044 66700 94096 66706
rect 94044 66642 94096 66648
rect 94516 66162 94544 66778
rect 94976 66570 95004 66778
rect 95712 66570 95740 67526
rect 95790 67487 95846 67496
rect 95896 67386 95924 68682
rect 96068 68196 96120 68202
rect 96068 68138 96120 68144
rect 95976 67584 96028 67590
rect 95976 67526 96028 67532
rect 95792 67380 95844 67386
rect 95792 67322 95844 67328
rect 95884 67380 95936 67386
rect 95884 67322 95936 67328
rect 94964 66564 95016 66570
rect 94964 66506 95016 66512
rect 95700 66564 95752 66570
rect 95700 66506 95752 66512
rect 95804 66502 95832 67322
rect 94872 66496 94924 66502
rect 94872 66438 94924 66444
rect 95792 66496 95844 66502
rect 95792 66438 95844 66444
rect 93952 66156 94004 66162
rect 93952 66098 94004 66104
rect 94504 66156 94556 66162
rect 94504 66098 94556 66104
rect 93492 66088 93544 66094
rect 92952 66014 93072 66042
rect 93492 66030 93544 66036
rect 93964 66026 93992 66098
rect 94884 66026 94912 66438
rect 95988 66094 96016 67526
rect 96080 66774 96108 68138
rect 96160 68128 96212 68134
rect 96160 68070 96212 68076
rect 96172 66842 96200 68070
rect 96374 68028 96682 68037
rect 96374 68026 96380 68028
rect 96436 68026 96460 68028
rect 96516 68026 96540 68028
rect 96596 68026 96620 68028
rect 96676 68026 96682 68028
rect 96436 67974 96438 68026
rect 96618 67974 96620 68026
rect 96374 67972 96380 67974
rect 96436 67972 96460 67974
rect 96516 67972 96540 67974
rect 96596 67972 96620 67974
rect 96676 67972 96682 67974
rect 96374 67963 96682 67972
rect 96620 67720 96672 67726
rect 96618 67688 96620 67697
rect 96672 67688 96674 67697
rect 96618 67623 96674 67632
rect 96710 67552 96766 67561
rect 96710 67487 96766 67496
rect 96724 67386 96752 67487
rect 96712 67380 96764 67386
rect 96712 67322 96764 67328
rect 96712 67244 96764 67250
rect 96712 67186 96764 67192
rect 96724 67046 96752 67186
rect 96804 67176 96856 67182
rect 96804 67118 96856 67124
rect 96252 67040 96304 67046
rect 96252 66982 96304 66988
rect 96712 67040 96764 67046
rect 96712 66982 96764 66988
rect 96264 66842 96292 66982
rect 96374 66940 96682 66949
rect 96374 66938 96380 66940
rect 96436 66938 96460 66940
rect 96516 66938 96540 66940
rect 96596 66938 96620 66940
rect 96676 66938 96682 66940
rect 96436 66886 96438 66938
rect 96618 66886 96620 66938
rect 96374 66884 96380 66886
rect 96436 66884 96460 66886
rect 96516 66884 96540 66886
rect 96596 66884 96620 66886
rect 96676 66884 96682 66886
rect 96374 66875 96682 66884
rect 96160 66836 96212 66842
rect 96160 66778 96212 66784
rect 96252 66836 96304 66842
rect 96252 66778 96304 66784
rect 96068 66768 96120 66774
rect 96068 66710 96120 66716
rect 96172 66638 96200 66778
rect 96160 66632 96212 66638
rect 96160 66574 96212 66580
rect 96160 66496 96212 66502
rect 96160 66438 96212 66444
rect 96068 66224 96120 66230
rect 96068 66166 96120 66172
rect 95976 66088 96028 66094
rect 95976 66030 96028 66036
rect 93044 65958 93072 66014
rect 93952 66020 94004 66026
rect 93952 65962 94004 65968
rect 94872 66020 94924 66026
rect 94872 65962 94924 65968
rect 93032 65952 93084 65958
rect 93032 65894 93084 65900
rect 93492 65952 93544 65958
rect 93492 65894 93544 65900
rect 93044 65754 93072 65894
rect 93032 65748 93084 65754
rect 93032 65690 93084 65696
rect 91744 65612 91796 65618
rect 91744 65554 91796 65560
rect 93504 65414 93532 65894
rect 93492 65408 93544 65414
rect 93492 65350 93544 65356
rect 96080 65210 96108 66166
rect 96068 65204 96120 65210
rect 96068 65146 96120 65152
rect 88524 64456 88576 64462
rect 88524 64398 88576 64404
rect 77392 64184 77444 64190
rect 75458 64152 75514 64161
rect 77392 64126 77444 64132
rect 75458 64087 75514 64096
rect 96172 63889 96200 66438
rect 96264 66144 96292 66778
rect 96724 66774 96752 66982
rect 96436 66768 96488 66774
rect 96436 66710 96488 66716
rect 96712 66768 96764 66774
rect 96712 66710 96764 66716
rect 96448 66230 96476 66710
rect 96620 66632 96672 66638
rect 96620 66574 96672 66580
rect 96436 66224 96488 66230
rect 96436 66166 96488 66172
rect 96344 66156 96396 66162
rect 96264 66116 96344 66144
rect 96344 66098 96396 66104
rect 96632 65958 96660 66574
rect 96712 66292 96764 66298
rect 96712 66234 96764 66240
rect 96620 65952 96672 65958
rect 96620 65894 96672 65900
rect 96374 65852 96682 65861
rect 96374 65850 96380 65852
rect 96436 65850 96460 65852
rect 96516 65850 96540 65852
rect 96596 65850 96620 65852
rect 96676 65850 96682 65852
rect 96436 65798 96438 65850
rect 96618 65798 96620 65850
rect 96374 65796 96380 65798
rect 96436 65796 96460 65798
rect 96516 65796 96540 65798
rect 96596 65796 96620 65798
rect 96676 65796 96682 65798
rect 96374 65787 96682 65796
rect 96724 65550 96752 66234
rect 96816 65958 96844 67118
rect 96908 66502 96936 69527
rect 97172 68672 97224 68678
rect 97172 68614 97224 68620
rect 97184 67930 97212 68614
rect 97172 67924 97224 67930
rect 97172 67866 97224 67872
rect 99196 67856 99248 67862
rect 96986 67824 97042 67833
rect 99196 67798 99248 67804
rect 96986 67759 96988 67768
rect 97040 67759 97042 67768
rect 96988 67730 97040 67736
rect 98184 67584 98236 67590
rect 98184 67526 98236 67532
rect 97034 67484 97342 67493
rect 97034 67482 97040 67484
rect 97096 67482 97120 67484
rect 97176 67482 97200 67484
rect 97256 67482 97280 67484
rect 97336 67482 97342 67484
rect 97096 67430 97098 67482
rect 97278 67430 97280 67482
rect 97034 67428 97040 67430
rect 97096 67428 97120 67430
rect 97176 67428 97200 67430
rect 97256 67428 97280 67430
rect 97336 67428 97342 67430
rect 97034 67419 97342 67428
rect 98196 67318 98224 67526
rect 98184 67312 98236 67318
rect 98184 67254 98236 67260
rect 99208 67250 99236 67798
rect 99748 67380 99800 67386
rect 99748 67322 99800 67328
rect 99380 67312 99432 67318
rect 99760 67266 99788 67322
rect 101968 67318 101996 83346
rect 102046 83323 102102 83332
rect 102048 75200 102100 75206
rect 102048 75142 102100 75148
rect 102060 67794 102088 75142
rect 102048 67788 102100 67794
rect 102048 67730 102100 67736
rect 99432 67260 99788 67266
rect 99380 67254 99788 67260
rect 101772 67312 101824 67318
rect 101772 67254 101824 67260
rect 101956 67312 102008 67318
rect 102152 67289 102180 128318
rect 105922 126780 106230 126789
rect 105922 126778 105928 126780
rect 105984 126778 106008 126780
rect 106064 126778 106088 126780
rect 106144 126778 106168 126780
rect 106224 126778 106230 126780
rect 105984 126726 105986 126778
rect 106166 126726 106168 126778
rect 105922 126724 105928 126726
rect 105984 126724 106008 126726
rect 106064 126724 106088 126726
rect 106144 126724 106168 126726
rect 106224 126724 106230 126726
rect 105922 126715 106230 126724
rect 102600 126472 102652 126478
rect 102600 126414 102652 126420
rect 102324 126404 102376 126410
rect 102324 126346 102376 126352
rect 102232 125724 102284 125730
rect 102232 125666 102284 125672
rect 102244 67561 102272 125666
rect 102230 67552 102286 67561
rect 102230 67487 102286 67496
rect 101956 67254 102008 67260
rect 102138 67280 102194 67289
rect 99196 67244 99248 67250
rect 99196 67186 99248 67192
rect 99392 67238 99788 67254
rect 98368 66632 98420 66638
rect 98368 66574 98420 66580
rect 98276 66564 98328 66570
rect 98276 66506 98328 66512
rect 96896 66496 96948 66502
rect 96896 66438 96948 66444
rect 97034 66396 97342 66405
rect 97034 66394 97040 66396
rect 97096 66394 97120 66396
rect 97176 66394 97200 66396
rect 97256 66394 97280 66396
rect 97336 66394 97342 66396
rect 97096 66342 97098 66394
rect 97278 66342 97280 66394
rect 97034 66340 97040 66342
rect 97096 66340 97120 66342
rect 97176 66340 97200 66342
rect 97256 66340 97280 66342
rect 97336 66340 97342 66342
rect 97034 66331 97342 66340
rect 98288 66298 98316 66506
rect 98276 66292 98328 66298
rect 98276 66234 98328 66240
rect 98380 66230 98408 66574
rect 99208 66298 99236 67186
rect 99392 66842 99420 67238
rect 99564 67176 99616 67182
rect 99564 67118 99616 67124
rect 99380 66836 99432 66842
rect 99380 66778 99432 66784
rect 99472 66836 99524 66842
rect 99472 66778 99524 66784
rect 99392 66298 99420 66778
rect 99484 66638 99512 66778
rect 99472 66632 99524 66638
rect 99472 66574 99524 66580
rect 99196 66292 99248 66298
rect 99196 66234 99248 66240
rect 99380 66292 99432 66298
rect 99380 66234 99432 66240
rect 98368 66224 98420 66230
rect 98368 66166 98420 66172
rect 99576 66026 99604 67118
rect 101784 66638 101812 67254
rect 102138 67215 102194 67224
rect 101864 67040 101916 67046
rect 101864 66982 101916 66988
rect 101876 66638 101904 66982
rect 102336 66745 102364 126346
rect 102416 126064 102468 126070
rect 102416 126006 102468 126012
rect 102428 68241 102456 126006
rect 102508 125860 102560 125866
rect 102508 125802 102560 125808
rect 102520 69834 102548 125802
rect 102508 69828 102560 69834
rect 102508 69770 102560 69776
rect 102612 69766 102640 126414
rect 106658 126236 106966 126245
rect 106658 126234 106664 126236
rect 106720 126234 106744 126236
rect 106800 126234 106824 126236
rect 106880 126234 106904 126236
rect 106960 126234 106966 126236
rect 106720 126182 106722 126234
rect 106902 126182 106904 126234
rect 106658 126180 106664 126182
rect 106720 126180 106744 126182
rect 106800 126180 106824 126182
rect 106880 126180 106904 126182
rect 106960 126180 106966 126182
rect 106658 126171 106966 126180
rect 103520 126132 103572 126138
rect 103520 126074 103572 126080
rect 102692 125996 102744 126002
rect 102692 125938 102744 125944
rect 102704 69970 102732 125938
rect 102782 123856 102838 123865
rect 102782 123791 102838 123800
rect 102796 77518 102824 123791
rect 103058 82240 103114 82249
rect 103058 82175 103114 82184
rect 102784 77512 102836 77518
rect 102784 77454 102836 77460
rect 102692 69964 102744 69970
rect 102692 69906 102744 69912
rect 102600 69760 102652 69766
rect 102600 69702 102652 69708
rect 102414 68232 102470 68241
rect 102414 68167 102470 68176
rect 102600 68196 102652 68202
rect 102600 68138 102652 68144
rect 102612 67590 102640 68138
rect 102600 67584 102652 67590
rect 102600 67526 102652 67532
rect 102796 67386 102824 77454
rect 102784 67380 102836 67386
rect 102784 67322 102836 67328
rect 103072 67114 103100 82175
rect 103532 69698 103560 126074
rect 103612 125928 103664 125934
rect 103612 125870 103664 125876
rect 103624 69902 103652 125870
rect 103704 125792 103756 125798
rect 103704 125734 103756 125740
rect 103716 70038 103744 125734
rect 105922 125692 106230 125701
rect 105922 125690 105928 125692
rect 105984 125690 106008 125692
rect 106064 125690 106088 125692
rect 106144 125690 106168 125692
rect 106224 125690 106230 125692
rect 105984 125638 105986 125690
rect 106166 125638 106168 125690
rect 105922 125636 105928 125638
rect 105984 125636 106008 125638
rect 106064 125636 106088 125638
rect 106144 125636 106168 125638
rect 106224 125636 106230 125638
rect 105922 125627 106230 125636
rect 106658 125148 106966 125157
rect 106658 125146 106664 125148
rect 106720 125146 106744 125148
rect 106800 125146 106824 125148
rect 106880 125146 106904 125148
rect 106960 125146 106966 125148
rect 106720 125094 106722 125146
rect 106902 125094 106904 125146
rect 106658 125092 106664 125094
rect 106720 125092 106744 125094
rect 106800 125092 106824 125094
rect 106880 125092 106904 125094
rect 106960 125092 106966 125094
rect 106658 125083 106966 125092
rect 105922 124604 106230 124613
rect 105922 124602 105928 124604
rect 105984 124602 106008 124604
rect 106064 124602 106088 124604
rect 106144 124602 106168 124604
rect 106224 124602 106230 124604
rect 105984 124550 105986 124602
rect 106166 124550 106168 124602
rect 105922 124548 105928 124550
rect 105984 124548 106008 124550
rect 106064 124548 106088 124550
rect 106144 124548 106168 124550
rect 106224 124548 106230 124550
rect 105922 124539 106230 124548
rect 106658 124060 106966 124069
rect 106658 124058 106664 124060
rect 106720 124058 106744 124060
rect 106800 124058 106824 124060
rect 106880 124058 106904 124060
rect 106960 124058 106966 124060
rect 106720 124006 106722 124058
rect 106902 124006 106904 124058
rect 106658 124004 106664 124006
rect 106720 124004 106744 124006
rect 106800 124004 106824 124006
rect 106880 124004 106904 124006
rect 106960 124004 106966 124006
rect 104714 123992 104770 124001
rect 106658 123995 106966 124004
rect 104714 123927 104770 123936
rect 104440 123752 104492 123758
rect 104440 123694 104492 123700
rect 104348 119944 104400 119950
rect 104348 119886 104400 119892
rect 104360 119785 104388 119886
rect 104346 119776 104402 119785
rect 104346 119711 104402 119720
rect 104452 85338 104480 123694
rect 104728 86426 104756 123927
rect 105922 123516 106230 123525
rect 105922 123514 105928 123516
rect 105984 123514 106008 123516
rect 106064 123514 106088 123516
rect 106144 123514 106168 123516
rect 106224 123514 106230 123516
rect 105984 123462 105986 123514
rect 106166 123462 106168 123514
rect 105922 123460 105928 123462
rect 105984 123460 106008 123462
rect 106064 123460 106088 123462
rect 106144 123460 106168 123462
rect 106224 123460 106230 123462
rect 105922 123451 106230 123460
rect 106658 122972 106966 122981
rect 106658 122970 106664 122972
rect 106720 122970 106744 122972
rect 106800 122970 106824 122972
rect 106880 122970 106904 122972
rect 106960 122970 106966 122972
rect 106720 122918 106722 122970
rect 106902 122918 106904 122970
rect 106658 122916 106664 122918
rect 106720 122916 106744 122918
rect 106800 122916 106824 122918
rect 106880 122916 106904 122918
rect 106960 122916 106966 122918
rect 106658 122907 106966 122916
rect 105922 122428 106230 122437
rect 105922 122426 105928 122428
rect 105984 122426 106008 122428
rect 106064 122426 106088 122428
rect 106144 122426 106168 122428
rect 106224 122426 106230 122428
rect 105984 122374 105986 122426
rect 106166 122374 106168 122426
rect 105922 122372 105928 122374
rect 105984 122372 106008 122374
rect 106064 122372 106088 122374
rect 106144 122372 106168 122374
rect 106224 122372 106230 122374
rect 105922 122363 106230 122372
rect 106658 121884 106966 121893
rect 106658 121882 106664 121884
rect 106720 121882 106744 121884
rect 106800 121882 106824 121884
rect 106880 121882 106904 121884
rect 106960 121882 106966 121884
rect 106720 121830 106722 121882
rect 106902 121830 106904 121882
rect 106658 121828 106664 121830
rect 106720 121828 106744 121830
rect 106800 121828 106824 121830
rect 106880 121828 106904 121830
rect 106960 121828 106966 121830
rect 106658 121819 106966 121828
rect 105922 121340 106230 121349
rect 105922 121338 105928 121340
rect 105984 121338 106008 121340
rect 106064 121338 106088 121340
rect 106144 121338 106168 121340
rect 106224 121338 106230 121340
rect 105984 121286 105986 121338
rect 106166 121286 106168 121338
rect 105922 121284 105928 121286
rect 105984 121284 106008 121286
rect 106064 121284 106088 121286
rect 106144 121284 106168 121286
rect 106224 121284 106230 121286
rect 105922 121275 106230 121284
rect 106658 120796 106966 120805
rect 106658 120794 106664 120796
rect 106720 120794 106744 120796
rect 106800 120794 106824 120796
rect 106880 120794 106904 120796
rect 106960 120794 106966 120796
rect 106720 120742 106722 120794
rect 106902 120742 106904 120794
rect 106658 120740 106664 120742
rect 106720 120740 106744 120742
rect 106800 120740 106824 120742
rect 106880 120740 106904 120742
rect 106960 120740 106966 120742
rect 106658 120731 106966 120740
rect 105922 120252 106230 120261
rect 105922 120250 105928 120252
rect 105984 120250 106008 120252
rect 106064 120250 106088 120252
rect 106144 120250 106168 120252
rect 106224 120250 106230 120252
rect 105984 120198 105986 120250
rect 106166 120198 106168 120250
rect 105922 120196 105928 120198
rect 105984 120196 106008 120198
rect 106064 120196 106088 120198
rect 106144 120196 106168 120198
rect 106224 120196 106230 120198
rect 105922 120187 106230 120196
rect 106658 119708 106966 119717
rect 106658 119706 106664 119708
rect 106720 119706 106744 119708
rect 106800 119706 106824 119708
rect 106880 119706 106904 119708
rect 106960 119706 106966 119708
rect 106720 119654 106722 119706
rect 106902 119654 106904 119706
rect 106658 119652 106664 119654
rect 106720 119652 106744 119654
rect 106800 119652 106824 119654
rect 106880 119652 106904 119654
rect 106960 119652 106966 119654
rect 106658 119643 106966 119652
rect 105922 119164 106230 119173
rect 105922 119162 105928 119164
rect 105984 119162 106008 119164
rect 106064 119162 106088 119164
rect 106144 119162 106168 119164
rect 106224 119162 106230 119164
rect 105984 119110 105986 119162
rect 106166 119110 106168 119162
rect 105922 119108 105928 119110
rect 105984 119108 106008 119110
rect 106064 119108 106088 119110
rect 106144 119108 106168 119110
rect 106224 119108 106230 119110
rect 105922 119099 106230 119108
rect 106658 118620 106966 118629
rect 106658 118618 106664 118620
rect 106720 118618 106744 118620
rect 106800 118618 106824 118620
rect 106880 118618 106904 118620
rect 106960 118618 106966 118620
rect 106720 118566 106722 118618
rect 106902 118566 106904 118618
rect 106658 118564 106664 118566
rect 106720 118564 106744 118566
rect 106800 118564 106824 118566
rect 106880 118564 106904 118566
rect 106960 118564 106966 118566
rect 106658 118555 106966 118564
rect 105922 118076 106230 118085
rect 105922 118074 105928 118076
rect 105984 118074 106008 118076
rect 106064 118074 106088 118076
rect 106144 118074 106168 118076
rect 106224 118074 106230 118076
rect 105984 118022 105986 118074
rect 106166 118022 106168 118074
rect 105922 118020 105928 118022
rect 105984 118020 106008 118022
rect 106064 118020 106088 118022
rect 106144 118020 106168 118022
rect 106224 118020 106230 118022
rect 105922 118011 106230 118020
rect 106658 117532 106966 117541
rect 106658 117530 106664 117532
rect 106720 117530 106744 117532
rect 106800 117530 106824 117532
rect 106880 117530 106904 117532
rect 106960 117530 106966 117532
rect 106720 117478 106722 117530
rect 106902 117478 106904 117530
rect 106658 117476 106664 117478
rect 106720 117476 106744 117478
rect 106800 117476 106824 117478
rect 106880 117476 106904 117478
rect 106960 117476 106966 117478
rect 106658 117467 106966 117476
rect 105922 116988 106230 116997
rect 105922 116986 105928 116988
rect 105984 116986 106008 116988
rect 106064 116986 106088 116988
rect 106144 116986 106168 116988
rect 106224 116986 106230 116988
rect 105984 116934 105986 116986
rect 106166 116934 106168 116986
rect 105922 116932 105928 116934
rect 105984 116932 106008 116934
rect 106064 116932 106088 116934
rect 106144 116932 106168 116934
rect 106224 116932 106230 116934
rect 105922 116923 106230 116932
rect 106658 116444 106966 116453
rect 106658 116442 106664 116444
rect 106720 116442 106744 116444
rect 106800 116442 106824 116444
rect 106880 116442 106904 116444
rect 106960 116442 106966 116444
rect 106720 116390 106722 116442
rect 106902 116390 106904 116442
rect 106658 116388 106664 116390
rect 106720 116388 106744 116390
rect 106800 116388 106824 116390
rect 106880 116388 106904 116390
rect 106960 116388 106966 116390
rect 106658 116379 106966 116388
rect 105922 115900 106230 115909
rect 105922 115898 105928 115900
rect 105984 115898 106008 115900
rect 106064 115898 106088 115900
rect 106144 115898 106168 115900
rect 106224 115898 106230 115900
rect 105984 115846 105986 115898
rect 106166 115846 106168 115898
rect 105922 115844 105928 115846
rect 105984 115844 106008 115846
rect 106064 115844 106088 115846
rect 106144 115844 106168 115846
rect 106224 115844 106230 115846
rect 105922 115835 106230 115844
rect 106658 115356 106966 115365
rect 106658 115354 106664 115356
rect 106720 115354 106744 115356
rect 106800 115354 106824 115356
rect 106880 115354 106904 115356
rect 106960 115354 106966 115356
rect 106720 115302 106722 115354
rect 106902 115302 106904 115354
rect 106658 115300 106664 115302
rect 106720 115300 106744 115302
rect 106800 115300 106824 115302
rect 106880 115300 106904 115302
rect 106960 115300 106966 115302
rect 106658 115291 106966 115300
rect 105922 114812 106230 114821
rect 105922 114810 105928 114812
rect 105984 114810 106008 114812
rect 106064 114810 106088 114812
rect 106144 114810 106168 114812
rect 106224 114810 106230 114812
rect 105984 114758 105986 114810
rect 106166 114758 106168 114810
rect 105922 114756 105928 114758
rect 105984 114756 106008 114758
rect 106064 114756 106088 114758
rect 106144 114756 106168 114758
rect 106224 114756 106230 114758
rect 105922 114747 106230 114756
rect 106658 114268 106966 114277
rect 106658 114266 106664 114268
rect 106720 114266 106744 114268
rect 106800 114266 106824 114268
rect 106880 114266 106904 114268
rect 106960 114266 106966 114268
rect 106720 114214 106722 114266
rect 106902 114214 106904 114266
rect 106658 114212 106664 114214
rect 106720 114212 106744 114214
rect 106800 114212 106824 114214
rect 106880 114212 106904 114214
rect 106960 114212 106966 114214
rect 106658 114203 106966 114212
rect 105922 113724 106230 113733
rect 105922 113722 105928 113724
rect 105984 113722 106008 113724
rect 106064 113722 106088 113724
rect 106144 113722 106168 113724
rect 106224 113722 106230 113724
rect 105984 113670 105986 113722
rect 106166 113670 106168 113722
rect 105922 113668 105928 113670
rect 105984 113668 106008 113670
rect 106064 113668 106088 113670
rect 106144 113668 106168 113670
rect 106224 113668 106230 113670
rect 105922 113659 106230 113668
rect 106658 113180 106966 113189
rect 106658 113178 106664 113180
rect 106720 113178 106744 113180
rect 106800 113178 106824 113180
rect 106880 113178 106904 113180
rect 106960 113178 106966 113180
rect 106720 113126 106722 113178
rect 106902 113126 106904 113178
rect 106658 113124 106664 113126
rect 106720 113124 106744 113126
rect 106800 113124 106824 113126
rect 106880 113124 106904 113126
rect 106960 113124 106966 113126
rect 106658 113115 106966 113124
rect 105922 112636 106230 112645
rect 105922 112634 105928 112636
rect 105984 112634 106008 112636
rect 106064 112634 106088 112636
rect 106144 112634 106168 112636
rect 106224 112634 106230 112636
rect 105984 112582 105986 112634
rect 106166 112582 106168 112634
rect 105922 112580 105928 112582
rect 105984 112580 106008 112582
rect 106064 112580 106088 112582
rect 106144 112580 106168 112582
rect 106224 112580 106230 112582
rect 105922 112571 106230 112580
rect 106658 112092 106966 112101
rect 106658 112090 106664 112092
rect 106720 112090 106744 112092
rect 106800 112090 106824 112092
rect 106880 112090 106904 112092
rect 106960 112090 106966 112092
rect 106720 112038 106722 112090
rect 106902 112038 106904 112090
rect 106658 112036 106664 112038
rect 106720 112036 106744 112038
rect 106800 112036 106824 112038
rect 106880 112036 106904 112038
rect 106960 112036 106966 112038
rect 106658 112027 106966 112036
rect 105922 111548 106230 111557
rect 105922 111546 105928 111548
rect 105984 111546 106008 111548
rect 106064 111546 106088 111548
rect 106144 111546 106168 111548
rect 106224 111546 106230 111548
rect 105984 111494 105986 111546
rect 106166 111494 106168 111546
rect 105922 111492 105928 111494
rect 105984 111492 106008 111494
rect 106064 111492 106088 111494
rect 106144 111492 106168 111494
rect 106224 111492 106230 111494
rect 105922 111483 106230 111492
rect 106658 111004 106966 111013
rect 106658 111002 106664 111004
rect 106720 111002 106744 111004
rect 106800 111002 106824 111004
rect 106880 111002 106904 111004
rect 106960 111002 106966 111004
rect 106720 110950 106722 111002
rect 106902 110950 106904 111002
rect 106658 110948 106664 110950
rect 106720 110948 106744 110950
rect 106800 110948 106824 110950
rect 106880 110948 106904 110950
rect 106960 110948 106966 110950
rect 106658 110939 106966 110948
rect 105922 110460 106230 110469
rect 105922 110458 105928 110460
rect 105984 110458 106008 110460
rect 106064 110458 106088 110460
rect 106144 110458 106168 110460
rect 106224 110458 106230 110460
rect 105984 110406 105986 110458
rect 106166 110406 106168 110458
rect 105922 110404 105928 110406
rect 105984 110404 106008 110406
rect 106064 110404 106088 110406
rect 106144 110404 106168 110406
rect 106224 110404 106230 110406
rect 105922 110395 106230 110404
rect 106658 109916 106966 109925
rect 106658 109914 106664 109916
rect 106720 109914 106744 109916
rect 106800 109914 106824 109916
rect 106880 109914 106904 109916
rect 106960 109914 106966 109916
rect 106720 109862 106722 109914
rect 106902 109862 106904 109914
rect 106658 109860 106664 109862
rect 106720 109860 106744 109862
rect 106800 109860 106824 109862
rect 106880 109860 106904 109862
rect 106960 109860 106966 109862
rect 106658 109851 106966 109860
rect 105922 109372 106230 109381
rect 105922 109370 105928 109372
rect 105984 109370 106008 109372
rect 106064 109370 106088 109372
rect 106144 109370 106168 109372
rect 106224 109370 106230 109372
rect 105984 109318 105986 109370
rect 106166 109318 106168 109370
rect 105922 109316 105928 109318
rect 105984 109316 106008 109318
rect 106064 109316 106088 109318
rect 106144 109316 106168 109318
rect 106224 109316 106230 109318
rect 105922 109307 106230 109316
rect 106658 108828 106966 108837
rect 106658 108826 106664 108828
rect 106720 108826 106744 108828
rect 106800 108826 106824 108828
rect 106880 108826 106904 108828
rect 106960 108826 106966 108828
rect 106720 108774 106722 108826
rect 106902 108774 106904 108826
rect 106658 108772 106664 108774
rect 106720 108772 106744 108774
rect 106800 108772 106824 108774
rect 106880 108772 106904 108774
rect 106960 108772 106966 108774
rect 106658 108763 106966 108772
rect 105922 108284 106230 108293
rect 105922 108282 105928 108284
rect 105984 108282 106008 108284
rect 106064 108282 106088 108284
rect 106144 108282 106168 108284
rect 106224 108282 106230 108284
rect 105984 108230 105986 108282
rect 106166 108230 106168 108282
rect 105922 108228 105928 108230
rect 105984 108228 106008 108230
rect 106064 108228 106088 108230
rect 106144 108228 106168 108230
rect 106224 108228 106230 108230
rect 105922 108219 106230 108228
rect 106658 107740 106966 107749
rect 106658 107738 106664 107740
rect 106720 107738 106744 107740
rect 106800 107738 106824 107740
rect 106880 107738 106904 107740
rect 106960 107738 106966 107740
rect 106720 107686 106722 107738
rect 106902 107686 106904 107738
rect 106658 107684 106664 107686
rect 106720 107684 106744 107686
rect 106800 107684 106824 107686
rect 106880 107684 106904 107686
rect 106960 107684 106966 107686
rect 106658 107675 106966 107684
rect 105922 107196 106230 107205
rect 105922 107194 105928 107196
rect 105984 107194 106008 107196
rect 106064 107194 106088 107196
rect 106144 107194 106168 107196
rect 106224 107194 106230 107196
rect 105984 107142 105986 107194
rect 106166 107142 106168 107194
rect 105922 107140 105928 107142
rect 105984 107140 106008 107142
rect 106064 107140 106088 107142
rect 106144 107140 106168 107142
rect 106224 107140 106230 107142
rect 105922 107131 106230 107140
rect 106658 106652 106966 106661
rect 106658 106650 106664 106652
rect 106720 106650 106744 106652
rect 106800 106650 106824 106652
rect 106880 106650 106904 106652
rect 106960 106650 106966 106652
rect 106720 106598 106722 106650
rect 106902 106598 106904 106650
rect 106658 106596 106664 106598
rect 106720 106596 106744 106598
rect 106800 106596 106824 106598
rect 106880 106596 106904 106598
rect 106960 106596 106966 106598
rect 106658 106587 106966 106596
rect 105922 106108 106230 106117
rect 105922 106106 105928 106108
rect 105984 106106 106008 106108
rect 106064 106106 106088 106108
rect 106144 106106 106168 106108
rect 106224 106106 106230 106108
rect 105984 106054 105986 106106
rect 106166 106054 106168 106106
rect 105922 106052 105928 106054
rect 105984 106052 106008 106054
rect 106064 106052 106088 106054
rect 106144 106052 106168 106054
rect 106224 106052 106230 106054
rect 105922 106043 106230 106052
rect 106658 105564 106966 105573
rect 106658 105562 106664 105564
rect 106720 105562 106744 105564
rect 106800 105562 106824 105564
rect 106880 105562 106904 105564
rect 106960 105562 106966 105564
rect 106720 105510 106722 105562
rect 106902 105510 106904 105562
rect 106658 105508 106664 105510
rect 106720 105508 106744 105510
rect 106800 105508 106824 105510
rect 106880 105508 106904 105510
rect 106960 105508 106966 105510
rect 106658 105499 106966 105508
rect 105922 105020 106230 105029
rect 105922 105018 105928 105020
rect 105984 105018 106008 105020
rect 106064 105018 106088 105020
rect 106144 105018 106168 105020
rect 106224 105018 106230 105020
rect 105984 104966 105986 105018
rect 106166 104966 106168 105018
rect 105922 104964 105928 104966
rect 105984 104964 106008 104966
rect 106064 104964 106088 104966
rect 106144 104964 106168 104966
rect 106224 104964 106230 104966
rect 105922 104955 106230 104964
rect 106658 104476 106966 104485
rect 106658 104474 106664 104476
rect 106720 104474 106744 104476
rect 106800 104474 106824 104476
rect 106880 104474 106904 104476
rect 106960 104474 106966 104476
rect 106720 104422 106722 104474
rect 106902 104422 106904 104474
rect 106658 104420 106664 104422
rect 106720 104420 106744 104422
rect 106800 104420 106824 104422
rect 106880 104420 106904 104422
rect 106960 104420 106966 104422
rect 106658 104411 106966 104420
rect 105922 103932 106230 103941
rect 105922 103930 105928 103932
rect 105984 103930 106008 103932
rect 106064 103930 106088 103932
rect 106144 103930 106168 103932
rect 106224 103930 106230 103932
rect 105984 103878 105986 103930
rect 106166 103878 106168 103930
rect 105922 103876 105928 103878
rect 105984 103876 106008 103878
rect 106064 103876 106088 103878
rect 106144 103876 106168 103878
rect 106224 103876 106230 103878
rect 105922 103867 106230 103876
rect 106658 103388 106966 103397
rect 106658 103386 106664 103388
rect 106720 103386 106744 103388
rect 106800 103386 106824 103388
rect 106880 103386 106904 103388
rect 106960 103386 106966 103388
rect 106720 103334 106722 103386
rect 106902 103334 106904 103386
rect 106658 103332 106664 103334
rect 106720 103332 106744 103334
rect 106800 103332 106824 103334
rect 106880 103332 106904 103334
rect 106960 103332 106966 103334
rect 106658 103323 106966 103332
rect 105922 102844 106230 102853
rect 105922 102842 105928 102844
rect 105984 102842 106008 102844
rect 106064 102842 106088 102844
rect 106144 102842 106168 102844
rect 106224 102842 106230 102844
rect 105984 102790 105986 102842
rect 106166 102790 106168 102842
rect 105922 102788 105928 102790
rect 105984 102788 106008 102790
rect 106064 102788 106088 102790
rect 106144 102788 106168 102790
rect 106224 102788 106230 102790
rect 105922 102779 106230 102788
rect 106658 102300 106966 102309
rect 106658 102298 106664 102300
rect 106720 102298 106744 102300
rect 106800 102298 106824 102300
rect 106880 102298 106904 102300
rect 106960 102298 106966 102300
rect 106720 102246 106722 102298
rect 106902 102246 106904 102298
rect 106658 102244 106664 102246
rect 106720 102244 106744 102246
rect 106800 102244 106824 102246
rect 106880 102244 106904 102246
rect 106960 102244 106966 102246
rect 106658 102235 106966 102244
rect 105922 101756 106230 101765
rect 105922 101754 105928 101756
rect 105984 101754 106008 101756
rect 106064 101754 106088 101756
rect 106144 101754 106168 101756
rect 106224 101754 106230 101756
rect 105984 101702 105986 101754
rect 106166 101702 106168 101754
rect 105922 101700 105928 101702
rect 105984 101700 106008 101702
rect 106064 101700 106088 101702
rect 106144 101700 106168 101702
rect 106224 101700 106230 101702
rect 105922 101691 106230 101700
rect 106658 101212 106966 101221
rect 106658 101210 106664 101212
rect 106720 101210 106744 101212
rect 106800 101210 106824 101212
rect 106880 101210 106904 101212
rect 106960 101210 106966 101212
rect 106720 101158 106722 101210
rect 106902 101158 106904 101210
rect 106658 101156 106664 101158
rect 106720 101156 106744 101158
rect 106800 101156 106824 101158
rect 106880 101156 106904 101158
rect 106960 101156 106966 101158
rect 106658 101147 106966 101156
rect 105922 100668 106230 100677
rect 105922 100666 105928 100668
rect 105984 100666 106008 100668
rect 106064 100666 106088 100668
rect 106144 100666 106168 100668
rect 106224 100666 106230 100668
rect 105984 100614 105986 100666
rect 106166 100614 106168 100666
rect 105922 100612 105928 100614
rect 105984 100612 106008 100614
rect 106064 100612 106088 100614
rect 106144 100612 106168 100614
rect 106224 100612 106230 100614
rect 105922 100603 106230 100612
rect 106658 100124 106966 100133
rect 106658 100122 106664 100124
rect 106720 100122 106744 100124
rect 106800 100122 106824 100124
rect 106880 100122 106904 100124
rect 106960 100122 106966 100124
rect 106720 100070 106722 100122
rect 106902 100070 106904 100122
rect 106658 100068 106664 100070
rect 106720 100068 106744 100070
rect 106800 100068 106824 100070
rect 106880 100068 106904 100070
rect 106960 100068 106966 100070
rect 106658 100059 106966 100068
rect 105922 99580 106230 99589
rect 105922 99578 105928 99580
rect 105984 99578 106008 99580
rect 106064 99578 106088 99580
rect 106144 99578 106168 99580
rect 106224 99578 106230 99580
rect 105984 99526 105986 99578
rect 106166 99526 106168 99578
rect 105922 99524 105928 99526
rect 105984 99524 106008 99526
rect 106064 99524 106088 99526
rect 106144 99524 106168 99526
rect 106224 99524 106230 99526
rect 105922 99515 106230 99524
rect 106658 99036 106966 99045
rect 106658 99034 106664 99036
rect 106720 99034 106744 99036
rect 106800 99034 106824 99036
rect 106880 99034 106904 99036
rect 106960 99034 106966 99036
rect 106720 98982 106722 99034
rect 106902 98982 106904 99034
rect 106658 98980 106664 98982
rect 106720 98980 106744 98982
rect 106800 98980 106824 98982
rect 106880 98980 106904 98982
rect 106960 98980 106966 98982
rect 106658 98971 106966 98980
rect 105922 98492 106230 98501
rect 105922 98490 105928 98492
rect 105984 98490 106008 98492
rect 106064 98490 106088 98492
rect 106144 98490 106168 98492
rect 106224 98490 106230 98492
rect 105984 98438 105986 98490
rect 106166 98438 106168 98490
rect 105922 98436 105928 98438
rect 105984 98436 106008 98438
rect 106064 98436 106088 98438
rect 106144 98436 106168 98438
rect 106224 98436 106230 98438
rect 105922 98427 106230 98436
rect 106658 97948 106966 97957
rect 106658 97946 106664 97948
rect 106720 97946 106744 97948
rect 106800 97946 106824 97948
rect 106880 97946 106904 97948
rect 106960 97946 106966 97948
rect 106720 97894 106722 97946
rect 106902 97894 106904 97946
rect 106658 97892 106664 97894
rect 106720 97892 106744 97894
rect 106800 97892 106824 97894
rect 106880 97892 106904 97894
rect 106960 97892 106966 97894
rect 106658 97883 106966 97892
rect 105922 97404 106230 97413
rect 105922 97402 105928 97404
rect 105984 97402 106008 97404
rect 106064 97402 106088 97404
rect 106144 97402 106168 97404
rect 106224 97402 106230 97404
rect 105984 97350 105986 97402
rect 106166 97350 106168 97402
rect 105922 97348 105928 97350
rect 105984 97348 106008 97350
rect 106064 97348 106088 97350
rect 106144 97348 106168 97350
rect 106224 97348 106230 97350
rect 105922 97339 106230 97348
rect 106658 96860 106966 96869
rect 106658 96858 106664 96860
rect 106720 96858 106744 96860
rect 106800 96858 106824 96860
rect 106880 96858 106904 96860
rect 106960 96858 106966 96860
rect 106720 96806 106722 96858
rect 106902 96806 106904 96858
rect 106658 96804 106664 96806
rect 106720 96804 106744 96806
rect 106800 96804 106824 96806
rect 106880 96804 106904 96806
rect 106960 96804 106966 96806
rect 106658 96795 106966 96804
rect 105922 96316 106230 96325
rect 105922 96314 105928 96316
rect 105984 96314 106008 96316
rect 106064 96314 106088 96316
rect 106144 96314 106168 96316
rect 106224 96314 106230 96316
rect 105984 96262 105986 96314
rect 106166 96262 106168 96314
rect 105922 96260 105928 96262
rect 105984 96260 106008 96262
rect 106064 96260 106088 96262
rect 106144 96260 106168 96262
rect 106224 96260 106230 96262
rect 105922 96251 106230 96260
rect 106658 95772 106966 95781
rect 106658 95770 106664 95772
rect 106720 95770 106744 95772
rect 106800 95770 106824 95772
rect 106880 95770 106904 95772
rect 106960 95770 106966 95772
rect 106720 95718 106722 95770
rect 106902 95718 106904 95770
rect 106658 95716 106664 95718
rect 106720 95716 106744 95718
rect 106800 95716 106824 95718
rect 106880 95716 106904 95718
rect 106960 95716 106966 95718
rect 106658 95707 106966 95716
rect 105922 95228 106230 95237
rect 105922 95226 105928 95228
rect 105984 95226 106008 95228
rect 106064 95226 106088 95228
rect 106144 95226 106168 95228
rect 106224 95226 106230 95228
rect 105984 95174 105986 95226
rect 106166 95174 106168 95226
rect 105922 95172 105928 95174
rect 105984 95172 106008 95174
rect 106064 95172 106088 95174
rect 106144 95172 106168 95174
rect 106224 95172 106230 95174
rect 105922 95163 106230 95172
rect 106658 94684 106966 94693
rect 106658 94682 106664 94684
rect 106720 94682 106744 94684
rect 106800 94682 106824 94684
rect 106880 94682 106904 94684
rect 106960 94682 106966 94684
rect 106720 94630 106722 94682
rect 106902 94630 106904 94682
rect 106658 94628 106664 94630
rect 106720 94628 106744 94630
rect 106800 94628 106824 94630
rect 106880 94628 106904 94630
rect 106960 94628 106966 94630
rect 106658 94619 106966 94628
rect 105922 94140 106230 94149
rect 105922 94138 105928 94140
rect 105984 94138 106008 94140
rect 106064 94138 106088 94140
rect 106144 94138 106168 94140
rect 106224 94138 106230 94140
rect 105984 94086 105986 94138
rect 106166 94086 106168 94138
rect 105922 94084 105928 94086
rect 105984 94084 106008 94086
rect 106064 94084 106088 94086
rect 106144 94084 106168 94086
rect 106224 94084 106230 94086
rect 105922 94075 106230 94084
rect 106658 93596 106966 93605
rect 106658 93594 106664 93596
rect 106720 93594 106744 93596
rect 106800 93594 106824 93596
rect 106880 93594 106904 93596
rect 106960 93594 106966 93596
rect 106720 93542 106722 93594
rect 106902 93542 106904 93594
rect 106658 93540 106664 93542
rect 106720 93540 106744 93542
rect 106800 93540 106824 93542
rect 106880 93540 106904 93542
rect 106960 93540 106966 93542
rect 106658 93531 106966 93540
rect 105922 93052 106230 93061
rect 105922 93050 105928 93052
rect 105984 93050 106008 93052
rect 106064 93050 106088 93052
rect 106144 93050 106168 93052
rect 106224 93050 106230 93052
rect 105984 92998 105986 93050
rect 106166 92998 106168 93050
rect 105922 92996 105928 92998
rect 105984 92996 106008 92998
rect 106064 92996 106088 92998
rect 106144 92996 106168 92998
rect 106224 92996 106230 92998
rect 105922 92987 106230 92996
rect 106658 92508 106966 92517
rect 106658 92506 106664 92508
rect 106720 92506 106744 92508
rect 106800 92506 106824 92508
rect 106880 92506 106904 92508
rect 106960 92506 106966 92508
rect 106720 92454 106722 92506
rect 106902 92454 106904 92506
rect 106658 92452 106664 92454
rect 106720 92452 106744 92454
rect 106800 92452 106824 92454
rect 106880 92452 106904 92454
rect 106960 92452 106966 92454
rect 106658 92443 106966 92452
rect 105922 91964 106230 91973
rect 105922 91962 105928 91964
rect 105984 91962 106008 91964
rect 106064 91962 106088 91964
rect 106144 91962 106168 91964
rect 106224 91962 106230 91964
rect 105984 91910 105986 91962
rect 106166 91910 106168 91962
rect 105922 91908 105928 91910
rect 105984 91908 106008 91910
rect 106064 91908 106088 91910
rect 106144 91908 106168 91910
rect 106224 91908 106230 91910
rect 105922 91899 106230 91908
rect 106658 91420 106966 91429
rect 106658 91418 106664 91420
rect 106720 91418 106744 91420
rect 106800 91418 106824 91420
rect 106880 91418 106904 91420
rect 106960 91418 106966 91420
rect 106720 91366 106722 91418
rect 106902 91366 106904 91418
rect 106658 91364 106664 91366
rect 106720 91364 106744 91366
rect 106800 91364 106824 91366
rect 106880 91364 106904 91366
rect 106960 91364 106966 91366
rect 106658 91355 106966 91364
rect 105922 90876 106230 90885
rect 105922 90874 105928 90876
rect 105984 90874 106008 90876
rect 106064 90874 106088 90876
rect 106144 90874 106168 90876
rect 106224 90874 106230 90876
rect 105984 90822 105986 90874
rect 106166 90822 106168 90874
rect 105922 90820 105928 90822
rect 105984 90820 106008 90822
rect 106064 90820 106088 90822
rect 106144 90820 106168 90822
rect 106224 90820 106230 90822
rect 105922 90811 106230 90820
rect 106658 90332 106966 90341
rect 106658 90330 106664 90332
rect 106720 90330 106744 90332
rect 106800 90330 106824 90332
rect 106880 90330 106904 90332
rect 106960 90330 106966 90332
rect 106720 90278 106722 90330
rect 106902 90278 106904 90330
rect 106658 90276 106664 90278
rect 106720 90276 106744 90278
rect 106800 90276 106824 90278
rect 106880 90276 106904 90278
rect 106960 90276 106966 90278
rect 106658 90267 106966 90276
rect 105922 89788 106230 89797
rect 105922 89786 105928 89788
rect 105984 89786 106008 89788
rect 106064 89786 106088 89788
rect 106144 89786 106168 89788
rect 106224 89786 106230 89788
rect 105984 89734 105986 89786
rect 106166 89734 106168 89786
rect 105922 89732 105928 89734
rect 105984 89732 106008 89734
rect 106064 89732 106088 89734
rect 106144 89732 106168 89734
rect 106224 89732 106230 89734
rect 105922 89723 106230 89732
rect 106658 89244 106966 89253
rect 106658 89242 106664 89244
rect 106720 89242 106744 89244
rect 106800 89242 106824 89244
rect 106880 89242 106904 89244
rect 106960 89242 106966 89244
rect 106720 89190 106722 89242
rect 106902 89190 106904 89242
rect 106658 89188 106664 89190
rect 106720 89188 106744 89190
rect 106800 89188 106824 89190
rect 106880 89188 106904 89190
rect 106960 89188 106966 89190
rect 106658 89179 106966 89188
rect 105922 88700 106230 88709
rect 105922 88698 105928 88700
rect 105984 88698 106008 88700
rect 106064 88698 106088 88700
rect 106144 88698 106168 88700
rect 106224 88698 106230 88700
rect 105984 88646 105986 88698
rect 106166 88646 106168 88698
rect 105922 88644 105928 88646
rect 105984 88644 106008 88646
rect 106064 88644 106088 88646
rect 106144 88644 106168 88646
rect 106224 88644 106230 88646
rect 105922 88635 106230 88644
rect 106658 88156 106966 88165
rect 106658 88154 106664 88156
rect 106720 88154 106744 88156
rect 106800 88154 106824 88156
rect 106880 88154 106904 88156
rect 106960 88154 106966 88156
rect 106720 88102 106722 88154
rect 106902 88102 106904 88154
rect 106658 88100 106664 88102
rect 106720 88100 106744 88102
rect 106800 88100 106824 88102
rect 106880 88100 106904 88102
rect 106960 88100 106966 88102
rect 106658 88091 106966 88100
rect 105922 87612 106230 87621
rect 105922 87610 105928 87612
rect 105984 87610 106008 87612
rect 106064 87610 106088 87612
rect 106144 87610 106168 87612
rect 106224 87610 106230 87612
rect 105984 87558 105986 87610
rect 106166 87558 106168 87610
rect 105922 87556 105928 87558
rect 105984 87556 106008 87558
rect 106064 87556 106088 87558
rect 106144 87556 106168 87558
rect 106224 87556 106230 87558
rect 105922 87547 106230 87556
rect 106658 87068 106966 87077
rect 106658 87066 106664 87068
rect 106720 87066 106744 87068
rect 106800 87066 106824 87068
rect 106880 87066 106904 87068
rect 106960 87066 106966 87068
rect 106720 87014 106722 87066
rect 106902 87014 106904 87066
rect 106658 87012 106664 87014
rect 106720 87012 106744 87014
rect 106800 87012 106824 87014
rect 106880 87012 106904 87014
rect 106960 87012 106966 87014
rect 106658 87003 106966 87012
rect 105922 86524 106230 86533
rect 105922 86522 105928 86524
rect 105984 86522 106008 86524
rect 106064 86522 106088 86524
rect 106144 86522 106168 86524
rect 106224 86522 106230 86524
rect 105984 86470 105986 86522
rect 106166 86470 106168 86522
rect 105922 86468 105928 86470
rect 105984 86468 106008 86470
rect 106064 86468 106088 86470
rect 106144 86468 106168 86470
rect 106224 86468 106230 86470
rect 105922 86459 106230 86468
rect 104716 86420 104768 86426
rect 104716 86362 104768 86368
rect 104808 86148 104860 86154
rect 104808 86090 104860 86096
rect 104716 85740 104768 85746
rect 104716 85682 104768 85688
rect 104440 85332 104492 85338
rect 104440 85274 104492 85280
rect 104728 85134 104756 85682
rect 104820 85678 104848 86090
rect 106658 85980 106966 85989
rect 106658 85978 106664 85980
rect 106720 85978 106744 85980
rect 106800 85978 106824 85980
rect 106880 85978 106904 85980
rect 106960 85978 106966 85980
rect 106720 85926 106722 85978
rect 106902 85926 106904 85978
rect 106658 85924 106664 85926
rect 106720 85924 106744 85926
rect 106800 85924 106824 85926
rect 106880 85924 106904 85926
rect 106960 85924 106966 85926
rect 106658 85915 106966 85924
rect 104808 85672 104860 85678
rect 104808 85614 104860 85620
rect 104716 85128 104768 85134
rect 104622 85096 104678 85105
rect 104716 85070 104768 85076
rect 104622 85031 104678 85040
rect 104164 80300 104216 80306
rect 104164 80242 104216 80248
rect 104072 79144 104124 79150
rect 104072 79086 104124 79092
rect 103888 79008 103940 79014
rect 103888 78950 103940 78956
rect 103900 78470 103928 78950
rect 104084 78538 104112 79086
rect 104072 78532 104124 78538
rect 104072 78474 104124 78480
rect 103888 78464 103940 78470
rect 103888 78406 103940 78412
rect 103900 75914 103928 78406
rect 103808 75886 103928 75914
rect 103704 70032 103756 70038
rect 103704 69974 103756 69980
rect 103612 69896 103664 69902
rect 103612 69838 103664 69844
rect 103520 69692 103572 69698
rect 103520 69634 103572 69640
rect 103808 68898 103836 75886
rect 104084 74534 104112 78474
rect 103992 74506 104112 74534
rect 103992 70394 104020 74506
rect 103624 68870 103836 68898
rect 103900 70366 104020 70394
rect 103624 67726 103652 68870
rect 103900 68762 103928 70366
rect 103716 68734 103928 68762
rect 103716 68678 103744 68734
rect 103704 68672 103756 68678
rect 103704 68614 103756 68620
rect 103796 68264 103848 68270
rect 103796 68206 103848 68212
rect 103704 68128 103756 68134
rect 103704 68070 103756 68076
rect 103612 67720 103664 67726
rect 103612 67662 103664 67668
rect 103060 67108 103112 67114
rect 103060 67050 103112 67056
rect 102322 66736 102378 66745
rect 102322 66671 102378 66680
rect 101772 66632 101824 66638
rect 101772 66574 101824 66580
rect 101864 66632 101916 66638
rect 102140 66632 102192 66638
rect 101864 66574 101916 66580
rect 102060 66580 102140 66586
rect 102060 66574 102192 66580
rect 101956 66564 102008 66570
rect 101956 66506 102008 66512
rect 102060 66558 102180 66574
rect 99748 66496 99800 66502
rect 99748 66438 99800 66444
rect 99760 66230 99788 66438
rect 99748 66224 99800 66230
rect 99748 66166 99800 66172
rect 100208 66156 100260 66162
rect 100208 66098 100260 66104
rect 99564 66020 99616 66026
rect 99564 65962 99616 65968
rect 100220 65958 100248 66098
rect 96804 65952 96856 65958
rect 96804 65894 96856 65900
rect 98368 65952 98420 65958
rect 98368 65894 98420 65900
rect 100208 65952 100260 65958
rect 100208 65894 100260 65900
rect 100576 65952 100628 65958
rect 100576 65894 100628 65900
rect 96712 65544 96764 65550
rect 96712 65486 96764 65492
rect 98380 65346 98408 65894
rect 100588 65618 100616 65894
rect 100576 65612 100628 65618
rect 100576 65554 100628 65560
rect 98368 65340 98420 65346
rect 98368 65282 98420 65288
rect 71870 63880 71926 63889
rect 71870 63815 71926 63824
rect 96158 63880 96214 63889
rect 96158 63815 96214 63824
rect 101968 23866 101996 66506
rect 102060 66162 102088 66558
rect 102140 66224 102192 66230
rect 102140 66166 102192 66172
rect 102048 66156 102100 66162
rect 102048 66098 102100 66104
rect 102152 35894 102180 66166
rect 103428 65340 103480 65346
rect 103428 65282 103480 65288
rect 102784 64184 102836 64190
rect 102784 64126 102836 64132
rect 102796 44946 102824 64126
rect 103440 59634 103468 65282
rect 103428 59628 103480 59634
rect 103428 59570 103480 59576
rect 102784 44940 102836 44946
rect 102784 44882 102836 44888
rect 103716 44334 103744 68070
rect 103808 67726 103836 68206
rect 104176 68134 104204 80242
rect 104532 80096 104584 80102
rect 104532 80038 104584 80044
rect 104440 78668 104492 78674
rect 104440 78610 104492 78616
rect 104256 78600 104308 78606
rect 104256 78542 104308 78548
rect 104268 76090 104296 78542
rect 104452 78266 104480 78610
rect 104440 78260 104492 78266
rect 104440 78202 104492 78208
rect 104440 78124 104492 78130
rect 104440 78066 104492 78072
rect 104452 77382 104480 78066
rect 104440 77376 104492 77382
rect 104440 77318 104492 77324
rect 104452 77058 104480 77318
rect 104360 77030 104480 77058
rect 104256 76084 104308 76090
rect 104256 76026 104308 76032
rect 104268 75342 104296 76026
rect 104256 75336 104308 75342
rect 104256 75278 104308 75284
rect 104164 68128 104216 68134
rect 104164 68070 104216 68076
rect 103796 67720 103848 67726
rect 103796 67662 103848 67668
rect 104360 67153 104388 77030
rect 104544 76022 104572 80038
rect 104636 78810 104664 85031
rect 104624 78804 104676 78810
rect 104624 78746 104676 78752
rect 104728 78470 104756 85070
rect 104820 78538 104848 85614
rect 105820 85604 105872 85610
rect 105820 85546 105872 85552
rect 105176 79144 105228 79150
rect 105176 79086 105228 79092
rect 105188 78606 105216 79086
rect 105176 78600 105228 78606
rect 105176 78542 105228 78548
rect 104808 78532 104860 78538
rect 104808 78474 104860 78480
rect 104716 78464 104768 78470
rect 104716 78406 104768 78412
rect 105544 78464 105596 78470
rect 105544 78406 105596 78412
rect 105556 78266 105584 78406
rect 104624 78260 104676 78266
rect 104624 78202 104676 78208
rect 105544 78260 105596 78266
rect 105544 78202 105596 78208
rect 104532 76016 104584 76022
rect 104532 75958 104584 75964
rect 104530 69864 104586 69873
rect 104530 69799 104586 69808
rect 104346 67144 104402 67153
rect 104346 67079 104402 67088
rect 104256 66836 104308 66842
rect 104256 66778 104308 66784
rect 103796 65952 103848 65958
rect 103796 65894 103848 65900
rect 103808 57526 103836 65894
rect 103888 65748 103940 65754
rect 103888 65690 103940 65696
rect 103796 57520 103848 57526
rect 103796 57462 103848 57468
rect 103796 55412 103848 55418
rect 103796 55354 103848 55360
rect 103704 44328 103756 44334
rect 103704 44270 103756 44276
rect 102152 35866 102364 35894
rect 102336 25097 102364 35866
rect 102600 25152 102652 25158
rect 102598 25120 102600 25129
rect 102652 25120 102654 25129
rect 102322 25088 102378 25097
rect 102598 25055 102654 25064
rect 102322 25023 102378 25032
rect 101956 23860 102008 23866
rect 101956 23802 102008 23808
rect 101968 23374 101996 23802
rect 102046 23388 102102 23397
rect 101968 23346 102046 23374
rect 102046 23323 102102 23332
rect 90732 10056 90784 10062
rect 90732 9998 90784 10004
rect 9586 9888 9642 9897
rect 4874 9820 5182 9829
rect 9586 9823 9642 9832
rect 16118 9888 16174 9897
rect 16118 9823 16174 9832
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 16132 7546 16160 9823
rect 90744 9761 90772 9998
rect 103808 9994 103836 55354
rect 103900 54874 103928 65690
rect 104164 65612 104216 65618
rect 104164 65554 104216 65560
rect 103980 60104 104032 60110
rect 103980 60046 104032 60052
rect 103992 59809 104020 60046
rect 103978 59800 104034 59809
rect 103978 59735 104034 59744
rect 103980 59560 104032 59566
rect 103980 59502 104032 59508
rect 103888 54868 103940 54874
rect 103888 54810 103940 54816
rect 103992 51542 104020 59502
rect 104176 56914 104204 65554
rect 104268 57594 104296 66778
rect 104360 58614 104388 67079
rect 104440 65204 104492 65210
rect 104440 65146 104492 65152
rect 104452 59770 104480 65146
rect 104544 60734 104572 69799
rect 104636 66774 104664 78202
rect 105636 77920 105688 77926
rect 105636 77862 105688 77868
rect 105648 77518 105676 77862
rect 105636 77512 105688 77518
rect 105636 77454 105688 77460
rect 105832 75886 105860 85546
rect 105922 85436 106230 85445
rect 105922 85434 105928 85436
rect 105984 85434 106008 85436
rect 106064 85434 106088 85436
rect 106144 85434 106168 85436
rect 106224 85434 106230 85436
rect 105984 85382 105986 85434
rect 106166 85382 106168 85434
rect 105922 85380 105928 85382
rect 105984 85380 106008 85382
rect 106064 85380 106088 85382
rect 106144 85380 106168 85382
rect 106224 85380 106230 85382
rect 105922 85371 106230 85380
rect 106658 84892 106966 84901
rect 106658 84890 106664 84892
rect 106720 84890 106744 84892
rect 106800 84890 106824 84892
rect 106880 84890 106904 84892
rect 106960 84890 106966 84892
rect 106720 84838 106722 84890
rect 106902 84838 106904 84890
rect 106658 84836 106664 84838
rect 106720 84836 106744 84838
rect 106800 84836 106824 84838
rect 106880 84836 106904 84838
rect 106960 84836 106966 84838
rect 106658 84827 106966 84836
rect 105922 84348 106230 84357
rect 105922 84346 105928 84348
rect 105984 84346 106008 84348
rect 106064 84346 106088 84348
rect 106144 84346 106168 84348
rect 106224 84346 106230 84348
rect 105984 84294 105986 84346
rect 106166 84294 106168 84346
rect 105922 84292 105928 84294
rect 105984 84292 106008 84294
rect 106064 84292 106088 84294
rect 106144 84292 106168 84294
rect 106224 84292 106230 84294
rect 105922 84283 106230 84292
rect 106658 83804 106966 83813
rect 106658 83802 106664 83804
rect 106720 83802 106744 83804
rect 106800 83802 106824 83804
rect 106880 83802 106904 83804
rect 106960 83802 106966 83804
rect 106720 83750 106722 83802
rect 106902 83750 106904 83802
rect 106658 83748 106664 83750
rect 106720 83748 106744 83750
rect 106800 83748 106824 83750
rect 106880 83748 106904 83750
rect 106960 83748 106966 83750
rect 106658 83739 106966 83748
rect 105922 83260 106230 83269
rect 105922 83258 105928 83260
rect 105984 83258 106008 83260
rect 106064 83258 106088 83260
rect 106144 83258 106168 83260
rect 106224 83258 106230 83260
rect 105984 83206 105986 83258
rect 106166 83206 106168 83258
rect 105922 83204 105928 83206
rect 105984 83204 106008 83206
rect 106064 83204 106088 83206
rect 106144 83204 106168 83206
rect 106224 83204 106230 83206
rect 105922 83195 106230 83204
rect 106658 82716 106966 82725
rect 106658 82714 106664 82716
rect 106720 82714 106744 82716
rect 106800 82714 106824 82716
rect 106880 82714 106904 82716
rect 106960 82714 106966 82716
rect 106720 82662 106722 82714
rect 106902 82662 106904 82714
rect 106658 82660 106664 82662
rect 106720 82660 106744 82662
rect 106800 82660 106824 82662
rect 106880 82660 106904 82662
rect 106960 82660 106966 82662
rect 106658 82651 106966 82660
rect 105922 82172 106230 82181
rect 105922 82170 105928 82172
rect 105984 82170 106008 82172
rect 106064 82170 106088 82172
rect 106144 82170 106168 82172
rect 106224 82170 106230 82172
rect 105984 82118 105986 82170
rect 106166 82118 106168 82170
rect 105922 82116 105928 82118
rect 105984 82116 106008 82118
rect 106064 82116 106088 82118
rect 106144 82116 106168 82118
rect 106224 82116 106230 82118
rect 105922 82107 106230 82116
rect 106658 81628 106966 81637
rect 106658 81626 106664 81628
rect 106720 81626 106744 81628
rect 106800 81626 106824 81628
rect 106880 81626 106904 81628
rect 106960 81626 106966 81628
rect 106720 81574 106722 81626
rect 106902 81574 106904 81626
rect 106658 81572 106664 81574
rect 106720 81572 106744 81574
rect 106800 81572 106824 81574
rect 106880 81572 106904 81574
rect 106960 81572 106966 81574
rect 106658 81563 106966 81572
rect 105922 81084 106230 81093
rect 105922 81082 105928 81084
rect 105984 81082 106008 81084
rect 106064 81082 106088 81084
rect 106144 81082 106168 81084
rect 106224 81082 106230 81084
rect 105984 81030 105986 81082
rect 106166 81030 106168 81082
rect 105922 81028 105928 81030
rect 105984 81028 106008 81030
rect 106064 81028 106088 81030
rect 106144 81028 106168 81030
rect 106224 81028 106230 81030
rect 105922 81019 106230 81028
rect 106658 80540 106966 80549
rect 106658 80538 106664 80540
rect 106720 80538 106744 80540
rect 106800 80538 106824 80540
rect 106880 80538 106904 80540
rect 106960 80538 106966 80540
rect 106720 80486 106722 80538
rect 106902 80486 106904 80538
rect 106658 80484 106664 80486
rect 106720 80484 106744 80486
rect 106800 80484 106824 80486
rect 106880 80484 106904 80486
rect 106960 80484 106966 80486
rect 106658 80475 106966 80484
rect 105922 79996 106230 80005
rect 105922 79994 105928 79996
rect 105984 79994 106008 79996
rect 106064 79994 106088 79996
rect 106144 79994 106168 79996
rect 106224 79994 106230 79996
rect 105984 79942 105986 79994
rect 106166 79942 106168 79994
rect 105922 79940 105928 79942
rect 105984 79940 106008 79942
rect 106064 79940 106088 79942
rect 106144 79940 106168 79942
rect 106224 79940 106230 79942
rect 105922 79931 106230 79940
rect 106658 79452 106966 79461
rect 106658 79450 106664 79452
rect 106720 79450 106744 79452
rect 106800 79450 106824 79452
rect 106880 79450 106904 79452
rect 106960 79450 106966 79452
rect 106720 79398 106722 79450
rect 106902 79398 106904 79450
rect 106658 79396 106664 79398
rect 106720 79396 106744 79398
rect 106800 79396 106824 79398
rect 106880 79396 106904 79398
rect 106960 79396 106966 79398
rect 106658 79387 106966 79396
rect 105922 78908 106230 78917
rect 105922 78906 105928 78908
rect 105984 78906 106008 78908
rect 106064 78906 106088 78908
rect 106144 78906 106168 78908
rect 106224 78906 106230 78908
rect 105984 78854 105986 78906
rect 106166 78854 106168 78906
rect 105922 78852 105928 78854
rect 105984 78852 106008 78854
rect 106064 78852 106088 78854
rect 106144 78852 106168 78854
rect 106224 78852 106230 78854
rect 105922 78843 106230 78852
rect 106658 78364 106966 78373
rect 106658 78362 106664 78364
rect 106720 78362 106744 78364
rect 106800 78362 106824 78364
rect 106880 78362 106904 78364
rect 106960 78362 106966 78364
rect 106720 78310 106722 78362
rect 106902 78310 106904 78362
rect 106658 78308 106664 78310
rect 106720 78308 106744 78310
rect 106800 78308 106824 78310
rect 106880 78308 106904 78310
rect 106960 78308 106966 78310
rect 106658 78299 106966 78308
rect 106280 77920 106332 77926
rect 106280 77862 106332 77868
rect 105922 77820 106230 77829
rect 105922 77818 105928 77820
rect 105984 77818 106008 77820
rect 106064 77818 106088 77820
rect 106144 77818 106168 77820
rect 106224 77818 106230 77820
rect 105984 77766 105986 77818
rect 106166 77766 106168 77818
rect 105922 77764 105928 77766
rect 105984 77764 106008 77766
rect 106064 77764 106088 77766
rect 106144 77764 106168 77766
rect 106224 77764 106230 77766
rect 105922 77755 106230 77764
rect 105922 76732 106230 76741
rect 105922 76730 105928 76732
rect 105984 76730 106008 76732
rect 106064 76730 106088 76732
rect 106144 76730 106168 76732
rect 106224 76730 106230 76732
rect 105984 76678 105986 76730
rect 106166 76678 106168 76730
rect 105922 76676 105928 76678
rect 105984 76676 106008 76678
rect 106064 76676 106088 76678
rect 106144 76676 106168 76678
rect 106224 76676 106230 76678
rect 105922 76667 106230 76676
rect 106292 76090 106320 77862
rect 106658 77276 106966 77285
rect 106658 77274 106664 77276
rect 106720 77274 106744 77276
rect 106800 77274 106824 77276
rect 106880 77274 106904 77276
rect 106960 77274 106966 77276
rect 106720 77222 106722 77274
rect 106902 77222 106904 77274
rect 106658 77220 106664 77222
rect 106720 77220 106744 77222
rect 106800 77220 106824 77222
rect 106880 77220 106904 77222
rect 106960 77220 106966 77222
rect 106658 77211 106966 77220
rect 106658 76188 106966 76197
rect 106658 76186 106664 76188
rect 106720 76186 106744 76188
rect 106800 76186 106824 76188
rect 106880 76186 106904 76188
rect 106960 76186 106966 76188
rect 106720 76134 106722 76186
rect 106902 76134 106904 76186
rect 106658 76132 106664 76134
rect 106720 76132 106744 76134
rect 106800 76132 106824 76134
rect 106880 76132 106904 76134
rect 106960 76132 106966 76134
rect 106658 76123 106966 76132
rect 106280 76084 106332 76090
rect 106280 76026 106332 76032
rect 105820 75880 105872 75886
rect 105820 75822 105872 75828
rect 105922 75644 106230 75653
rect 105922 75642 105928 75644
rect 105984 75642 106008 75644
rect 106064 75642 106088 75644
rect 106144 75642 106168 75644
rect 106224 75642 106230 75644
rect 105984 75590 105986 75642
rect 106166 75590 106168 75642
rect 105922 75588 105928 75590
rect 105984 75588 106008 75590
rect 106064 75588 106088 75590
rect 106144 75588 106168 75590
rect 106224 75588 106230 75590
rect 105922 75579 106230 75588
rect 106658 75100 106966 75109
rect 106658 75098 106664 75100
rect 106720 75098 106744 75100
rect 106800 75098 106824 75100
rect 106880 75098 106904 75100
rect 106960 75098 106966 75100
rect 106720 75046 106722 75098
rect 106902 75046 106904 75098
rect 106658 75044 106664 75046
rect 106720 75044 106744 75046
rect 106800 75044 106824 75046
rect 106880 75044 106904 75046
rect 106960 75044 106966 75046
rect 106658 75035 106966 75044
rect 105922 74556 106230 74565
rect 105922 74554 105928 74556
rect 105984 74554 106008 74556
rect 106064 74554 106088 74556
rect 106144 74554 106168 74556
rect 106224 74554 106230 74556
rect 105984 74502 105986 74554
rect 106166 74502 106168 74554
rect 105922 74500 105928 74502
rect 105984 74500 106008 74502
rect 106064 74500 106088 74502
rect 106144 74500 106168 74502
rect 106224 74500 106230 74502
rect 105922 74491 106230 74500
rect 106658 74012 106966 74021
rect 106658 74010 106664 74012
rect 106720 74010 106744 74012
rect 106800 74010 106824 74012
rect 106880 74010 106904 74012
rect 106960 74010 106966 74012
rect 106720 73958 106722 74010
rect 106902 73958 106904 74010
rect 106658 73956 106664 73958
rect 106720 73956 106744 73958
rect 106800 73956 106824 73958
rect 106880 73956 106904 73958
rect 106960 73956 106966 73958
rect 106658 73947 106966 73956
rect 105922 73468 106230 73477
rect 105922 73466 105928 73468
rect 105984 73466 106008 73468
rect 106064 73466 106088 73468
rect 106144 73466 106168 73468
rect 106224 73466 106230 73468
rect 105984 73414 105986 73466
rect 106166 73414 106168 73466
rect 105922 73412 105928 73414
rect 105984 73412 106008 73414
rect 106064 73412 106088 73414
rect 106144 73412 106168 73414
rect 106224 73412 106230 73414
rect 105922 73403 106230 73412
rect 106658 72924 106966 72933
rect 106658 72922 106664 72924
rect 106720 72922 106744 72924
rect 106800 72922 106824 72924
rect 106880 72922 106904 72924
rect 106960 72922 106966 72924
rect 106720 72870 106722 72922
rect 106902 72870 106904 72922
rect 106658 72868 106664 72870
rect 106720 72868 106744 72870
rect 106800 72868 106824 72870
rect 106880 72868 106904 72870
rect 106960 72868 106966 72870
rect 106658 72859 106966 72868
rect 105922 72380 106230 72389
rect 105922 72378 105928 72380
rect 105984 72378 106008 72380
rect 106064 72378 106088 72380
rect 106144 72378 106168 72380
rect 106224 72378 106230 72380
rect 105984 72326 105986 72378
rect 106166 72326 106168 72378
rect 105922 72324 105928 72326
rect 105984 72324 106008 72326
rect 106064 72324 106088 72326
rect 106144 72324 106168 72326
rect 106224 72324 106230 72326
rect 105922 72315 106230 72324
rect 106658 71836 106966 71845
rect 106658 71834 106664 71836
rect 106720 71834 106744 71836
rect 106800 71834 106824 71836
rect 106880 71834 106904 71836
rect 106960 71834 106966 71836
rect 106720 71782 106722 71834
rect 106902 71782 106904 71834
rect 106658 71780 106664 71782
rect 106720 71780 106744 71782
rect 106800 71780 106824 71782
rect 106880 71780 106904 71782
rect 106960 71780 106966 71782
rect 106658 71771 106966 71780
rect 105922 71292 106230 71301
rect 105922 71290 105928 71292
rect 105984 71290 106008 71292
rect 106064 71290 106088 71292
rect 106144 71290 106168 71292
rect 106224 71290 106230 71292
rect 105984 71238 105986 71290
rect 106166 71238 106168 71290
rect 105922 71236 105928 71238
rect 105984 71236 106008 71238
rect 106064 71236 106088 71238
rect 106144 71236 106168 71238
rect 106224 71236 106230 71238
rect 105922 71227 106230 71236
rect 106658 70748 106966 70757
rect 106658 70746 106664 70748
rect 106720 70746 106744 70748
rect 106800 70746 106824 70748
rect 106880 70746 106904 70748
rect 106960 70746 106966 70748
rect 106720 70694 106722 70746
rect 106902 70694 106904 70746
rect 106658 70692 106664 70694
rect 106720 70692 106744 70694
rect 106800 70692 106824 70694
rect 106880 70692 106904 70694
rect 106960 70692 106966 70694
rect 106658 70683 106966 70692
rect 105922 70204 106230 70213
rect 105922 70202 105928 70204
rect 105984 70202 106008 70204
rect 106064 70202 106088 70204
rect 106144 70202 106168 70204
rect 106224 70202 106230 70204
rect 105984 70150 105986 70202
rect 106166 70150 106168 70202
rect 105922 70148 105928 70150
rect 105984 70148 106008 70150
rect 106064 70148 106088 70150
rect 106144 70148 106168 70150
rect 106224 70148 106230 70150
rect 105922 70139 106230 70148
rect 107568 69760 107620 69766
rect 107568 69702 107620 69708
rect 108488 69760 108540 69766
rect 108488 69702 108540 69708
rect 106658 69660 106966 69669
rect 106658 69658 106664 69660
rect 106720 69658 106744 69660
rect 106800 69658 106824 69660
rect 106880 69658 106904 69660
rect 106960 69658 106966 69660
rect 106720 69606 106722 69658
rect 106902 69606 106904 69658
rect 106658 69604 106664 69606
rect 106720 69604 106744 69606
rect 106800 69604 106824 69606
rect 106880 69604 106904 69606
rect 106960 69604 106966 69606
rect 106658 69595 106966 69604
rect 105922 69116 106230 69125
rect 105922 69114 105928 69116
rect 105984 69114 106008 69116
rect 106064 69114 106088 69116
rect 106144 69114 106168 69116
rect 106224 69114 106230 69116
rect 105984 69062 105986 69114
rect 106166 69062 106168 69114
rect 105922 69060 105928 69062
rect 105984 69060 106008 69062
rect 106064 69060 106088 69062
rect 106144 69060 106168 69062
rect 106224 69060 106230 69062
rect 105922 69051 106230 69060
rect 106658 68572 106966 68581
rect 106658 68570 106664 68572
rect 106720 68570 106744 68572
rect 106800 68570 106824 68572
rect 106880 68570 106904 68572
rect 106960 68570 106966 68572
rect 106720 68518 106722 68570
rect 106902 68518 106904 68570
rect 106658 68516 106664 68518
rect 106720 68516 106744 68518
rect 106800 68516 106824 68518
rect 106880 68516 106904 68518
rect 106960 68516 106966 68518
rect 106658 68507 106966 68516
rect 105922 68028 106230 68037
rect 105922 68026 105928 68028
rect 105984 68026 106008 68028
rect 106064 68026 106088 68028
rect 106144 68026 106168 68028
rect 106224 68026 106230 68028
rect 105984 67974 105986 68026
rect 106166 67974 106168 68026
rect 105922 67972 105928 67974
rect 105984 67972 106008 67974
rect 106064 67972 106088 67974
rect 106144 67972 106168 67974
rect 106224 67972 106230 67974
rect 105922 67963 106230 67972
rect 106658 67484 106966 67493
rect 106658 67482 106664 67484
rect 106720 67482 106744 67484
rect 106800 67482 106824 67484
rect 106880 67482 106904 67484
rect 106960 67482 106966 67484
rect 106720 67430 106722 67482
rect 106902 67430 106904 67482
rect 106658 67428 106664 67430
rect 106720 67428 106744 67430
rect 106800 67428 106824 67430
rect 106880 67428 106904 67430
rect 106960 67428 106966 67430
rect 106658 67419 106966 67428
rect 106188 67040 106240 67046
rect 106188 66982 106240 66988
rect 104624 66768 104676 66774
rect 104624 66710 104676 66716
rect 106200 66609 106228 66982
rect 106186 66600 106242 66609
rect 106186 66535 106242 66544
rect 104808 66496 104860 66502
rect 104808 66438 104860 66444
rect 104544 60706 104664 60734
rect 104440 59764 104492 59770
rect 104440 59706 104492 59712
rect 104348 58608 104400 58614
rect 104348 58550 104400 58556
rect 104360 58138 104388 58550
rect 104348 58132 104400 58138
rect 104348 58074 104400 58080
rect 104256 57588 104308 57594
rect 104256 57530 104308 57536
rect 104532 57588 104584 57594
rect 104532 57530 104584 57536
rect 104164 56908 104216 56914
rect 104164 56850 104216 56856
rect 104440 56908 104492 56914
rect 104440 56850 104492 56856
rect 104176 56506 104204 56850
rect 104256 56840 104308 56846
rect 104256 56782 104308 56788
rect 104164 56500 104216 56506
rect 104164 56442 104216 56448
rect 103980 51536 104032 51542
rect 103980 51478 104032 51484
rect 104268 49910 104296 56782
rect 104348 56704 104400 56710
rect 104348 56646 104400 56652
rect 104360 56370 104388 56646
rect 104348 56364 104400 56370
rect 104348 56306 104400 56312
rect 104256 49904 104308 49910
rect 104256 49846 104308 49852
rect 104268 49434 104296 49846
rect 104360 49842 104388 56306
rect 104452 54806 104480 56850
rect 104544 56710 104572 57530
rect 104532 56704 104584 56710
rect 104532 56646 104584 56652
rect 104544 55350 104572 56646
rect 104636 56438 104664 60706
rect 104716 57520 104768 57526
rect 104716 57462 104768 57468
rect 104728 56914 104756 57462
rect 104820 56914 104848 66438
rect 106658 66396 106966 66405
rect 106658 66394 106664 66396
rect 106720 66394 106744 66396
rect 106800 66394 106824 66396
rect 106880 66394 106904 66396
rect 106960 66394 106966 66396
rect 106720 66342 106722 66394
rect 106902 66342 106904 66394
rect 106658 66340 106664 66342
rect 106720 66340 106744 66342
rect 106800 66340 106824 66342
rect 106880 66340 106904 66342
rect 106960 66340 106966 66342
rect 106658 66331 106966 66340
rect 105922 65852 106230 65861
rect 105922 65850 105928 65852
rect 105984 65850 106008 65852
rect 106064 65850 106088 65852
rect 106144 65850 106168 65852
rect 106224 65850 106230 65852
rect 105984 65798 105986 65850
rect 106166 65798 106168 65850
rect 105922 65796 105928 65798
rect 105984 65796 106008 65798
rect 106064 65796 106088 65798
rect 106144 65796 106168 65798
rect 106224 65796 106230 65798
rect 105922 65787 106230 65796
rect 107580 65482 107608 69702
rect 108500 69465 108528 69702
rect 108486 69456 108542 69465
rect 108486 69391 108542 69400
rect 108486 68776 108542 68785
rect 108486 68711 108542 68720
rect 108500 68678 108528 68711
rect 108488 68672 108540 68678
rect 108488 68614 108540 68620
rect 108488 68128 108540 68134
rect 108486 68096 108488 68105
rect 108540 68096 108542 68105
rect 108486 68031 108542 68040
rect 108488 67856 108540 67862
rect 108488 67798 108540 67804
rect 108500 67425 108528 67798
rect 108486 67416 108542 67425
rect 108486 67351 108542 67360
rect 108488 67040 108540 67046
rect 108488 66982 108540 66988
rect 108500 66745 108528 66982
rect 108486 66736 108542 66745
rect 108486 66671 108542 66680
rect 108304 66156 108356 66162
rect 108304 66098 108356 66104
rect 108316 65686 108344 66098
rect 108486 66056 108542 66065
rect 108486 65991 108488 66000
rect 108540 65991 108542 66000
rect 108488 65962 108540 65968
rect 108304 65680 108356 65686
rect 108304 65622 108356 65628
rect 107568 65476 107620 65482
rect 107568 65418 107620 65424
rect 104992 65408 105044 65414
rect 108488 65408 108540 65414
rect 104992 65350 105044 65356
rect 108486 65376 108488 65385
rect 108540 65376 108542 65385
rect 105004 57050 105032 65350
rect 106658 65308 106966 65317
rect 108486 65311 108542 65320
rect 106658 65306 106664 65308
rect 106720 65306 106744 65308
rect 106800 65306 106824 65308
rect 106880 65306 106904 65308
rect 106960 65306 106966 65308
rect 106720 65254 106722 65306
rect 106902 65254 106904 65306
rect 106658 65252 106664 65254
rect 106720 65252 106744 65254
rect 106800 65252 106824 65254
rect 106880 65252 106904 65254
rect 106960 65252 106966 65254
rect 106658 65243 106966 65252
rect 108488 64932 108540 64938
rect 108488 64874 108540 64880
rect 105922 64764 106230 64773
rect 105922 64762 105928 64764
rect 105984 64762 106008 64764
rect 106064 64762 106088 64764
rect 106144 64762 106168 64764
rect 106224 64762 106230 64764
rect 105984 64710 105986 64762
rect 106166 64710 106168 64762
rect 105922 64708 105928 64710
rect 105984 64708 106008 64710
rect 106064 64708 106088 64710
rect 106144 64708 106168 64710
rect 106224 64708 106230 64710
rect 105922 64699 106230 64708
rect 108500 64705 108528 64874
rect 108486 64696 108542 64705
rect 108486 64631 108542 64640
rect 108488 64320 108540 64326
rect 108488 64262 108540 64268
rect 106658 64220 106966 64229
rect 106658 64218 106664 64220
rect 106720 64218 106744 64220
rect 106800 64218 106824 64220
rect 106880 64218 106904 64220
rect 106960 64218 106966 64220
rect 106720 64166 106722 64218
rect 106902 64166 106904 64218
rect 106658 64164 106664 64166
rect 106720 64164 106744 64166
rect 106800 64164 106824 64166
rect 106880 64164 106904 64166
rect 106960 64164 106966 64166
rect 106658 64155 106966 64164
rect 108500 64025 108528 64262
rect 108486 64016 108542 64025
rect 108486 63951 108542 63960
rect 105634 63880 105690 63889
rect 105634 63815 105690 63824
rect 105648 58682 105676 63815
rect 105922 63676 106230 63685
rect 105922 63674 105928 63676
rect 105984 63674 106008 63676
rect 106064 63674 106088 63676
rect 106144 63674 106168 63676
rect 106224 63674 106230 63676
rect 105984 63622 105986 63674
rect 106166 63622 106168 63674
rect 105922 63620 105928 63622
rect 105984 63620 106008 63622
rect 106064 63620 106088 63622
rect 106144 63620 106168 63622
rect 106224 63620 106230 63622
rect 105922 63611 106230 63620
rect 106658 63132 106966 63141
rect 106658 63130 106664 63132
rect 106720 63130 106744 63132
rect 106800 63130 106824 63132
rect 106880 63130 106904 63132
rect 106960 63130 106966 63132
rect 106720 63078 106722 63130
rect 106902 63078 106904 63130
rect 106658 63076 106664 63078
rect 106720 63076 106744 63078
rect 106800 63076 106824 63078
rect 106880 63076 106904 63078
rect 106960 63076 106966 63078
rect 106658 63067 106966 63076
rect 105922 62588 106230 62597
rect 105922 62586 105928 62588
rect 105984 62586 106008 62588
rect 106064 62586 106088 62588
rect 106144 62586 106168 62588
rect 106224 62586 106230 62588
rect 105984 62534 105986 62586
rect 106166 62534 106168 62586
rect 105922 62532 105928 62534
rect 105984 62532 106008 62534
rect 106064 62532 106088 62534
rect 106144 62532 106168 62534
rect 106224 62532 106230 62534
rect 105922 62523 106230 62532
rect 106658 62044 106966 62053
rect 106658 62042 106664 62044
rect 106720 62042 106744 62044
rect 106800 62042 106824 62044
rect 106880 62042 106904 62044
rect 106960 62042 106966 62044
rect 106720 61990 106722 62042
rect 106902 61990 106904 62042
rect 106658 61988 106664 61990
rect 106720 61988 106744 61990
rect 106800 61988 106824 61990
rect 106880 61988 106904 61990
rect 106960 61988 106966 61990
rect 106658 61979 106966 61988
rect 105922 61500 106230 61509
rect 105922 61498 105928 61500
rect 105984 61498 106008 61500
rect 106064 61498 106088 61500
rect 106144 61498 106168 61500
rect 106224 61498 106230 61500
rect 105984 61446 105986 61498
rect 106166 61446 106168 61498
rect 105922 61444 105928 61446
rect 105984 61444 106008 61446
rect 106064 61444 106088 61446
rect 106144 61444 106168 61446
rect 106224 61444 106230 61446
rect 105922 61435 106230 61444
rect 106658 60956 106966 60965
rect 106658 60954 106664 60956
rect 106720 60954 106744 60956
rect 106800 60954 106824 60956
rect 106880 60954 106904 60956
rect 106960 60954 106966 60956
rect 106720 60902 106722 60954
rect 106902 60902 106904 60954
rect 106658 60900 106664 60902
rect 106720 60900 106744 60902
rect 106800 60900 106824 60902
rect 106880 60900 106904 60902
rect 106960 60900 106966 60902
rect 106658 60891 106966 60900
rect 105922 60412 106230 60421
rect 105922 60410 105928 60412
rect 105984 60410 106008 60412
rect 106064 60410 106088 60412
rect 106144 60410 106168 60412
rect 106224 60410 106230 60412
rect 105984 60358 105986 60410
rect 106166 60358 106168 60410
rect 105922 60356 105928 60358
rect 105984 60356 106008 60358
rect 106064 60356 106088 60358
rect 106144 60356 106168 60358
rect 106224 60356 106230 60358
rect 105922 60347 106230 60356
rect 106658 59868 106966 59877
rect 106658 59866 106664 59868
rect 106720 59866 106744 59868
rect 106800 59866 106824 59868
rect 106880 59866 106904 59868
rect 106960 59866 106966 59868
rect 106720 59814 106722 59866
rect 106902 59814 106904 59866
rect 106658 59812 106664 59814
rect 106720 59812 106744 59814
rect 106800 59812 106824 59814
rect 106880 59812 106904 59814
rect 106960 59812 106966 59814
rect 106658 59803 106966 59812
rect 105922 59324 106230 59333
rect 105922 59322 105928 59324
rect 105984 59322 106008 59324
rect 106064 59322 106088 59324
rect 106144 59322 106168 59324
rect 106224 59322 106230 59324
rect 105984 59270 105986 59322
rect 106166 59270 106168 59322
rect 105922 59268 105928 59270
rect 105984 59268 106008 59270
rect 106064 59268 106088 59270
rect 106144 59268 106168 59270
rect 106224 59268 106230 59270
rect 105922 59259 106230 59268
rect 106658 58780 106966 58789
rect 106658 58778 106664 58780
rect 106720 58778 106744 58780
rect 106800 58778 106824 58780
rect 106880 58778 106904 58780
rect 106960 58778 106966 58780
rect 106720 58726 106722 58778
rect 106902 58726 106904 58778
rect 106658 58724 106664 58726
rect 106720 58724 106744 58726
rect 106800 58724 106824 58726
rect 106880 58724 106904 58726
rect 106960 58724 106966 58726
rect 106658 58715 106966 58724
rect 105636 58676 105688 58682
rect 105636 58618 105688 58624
rect 105820 58676 105872 58682
rect 105820 58618 105872 58624
rect 104992 57044 105044 57050
rect 104992 56986 105044 56992
rect 104716 56908 104768 56914
rect 104716 56850 104768 56856
rect 104808 56908 104860 56914
rect 104808 56850 104860 56856
rect 104716 56500 104768 56506
rect 104716 56442 104768 56448
rect 104624 56432 104676 56438
rect 104624 56374 104676 56380
rect 104532 55344 104584 55350
rect 104532 55286 104584 55292
rect 104440 54800 104492 54806
rect 104440 54742 104492 54748
rect 104452 54330 104480 54742
rect 104544 54670 104572 55286
rect 104728 55214 104756 56442
rect 104636 55186 104756 55214
rect 104532 54664 104584 54670
rect 104532 54606 104584 54612
rect 104544 54330 104572 54606
rect 104636 54534 104664 55186
rect 104624 54528 104676 54534
rect 104624 54470 104676 54476
rect 104716 54528 104768 54534
rect 104716 54470 104768 54476
rect 104440 54324 104492 54330
rect 104440 54266 104492 54272
rect 104532 54324 104584 54330
rect 104532 54266 104584 54272
rect 104452 51338 104480 54266
rect 104544 52154 104572 54266
rect 104532 52148 104584 52154
rect 104532 52090 104584 52096
rect 104544 51610 104572 52090
rect 104532 51604 104584 51610
rect 104532 51546 104584 51552
rect 104636 51490 104664 54470
rect 104544 51462 104664 51490
rect 104440 51332 104492 51338
rect 104440 51274 104492 51280
rect 104452 51066 104480 51274
rect 104544 51270 104572 51462
rect 104624 51400 104676 51406
rect 104624 51342 104676 51348
rect 104532 51264 104584 51270
rect 104532 51206 104584 51212
rect 104544 51066 104572 51206
rect 104440 51060 104492 51066
rect 104440 51002 104492 51008
rect 104532 51060 104584 51066
rect 104532 51002 104584 51008
rect 104348 49836 104400 49842
rect 104348 49778 104400 49784
rect 104256 49428 104308 49434
rect 104256 49370 104308 49376
rect 104360 46170 104388 49778
rect 104348 46164 104400 46170
rect 104348 46106 104400 46112
rect 104256 45960 104308 45966
rect 104256 45902 104308 45908
rect 104268 42226 104296 45902
rect 104636 45422 104664 51342
rect 104728 49978 104756 54470
rect 105360 51264 105412 51270
rect 105360 51206 105412 51212
rect 104716 49972 104768 49978
rect 104716 49914 104768 49920
rect 104808 49768 104860 49774
rect 104808 49710 104860 49716
rect 104624 45416 104676 45422
rect 104624 45358 104676 45364
rect 104716 44192 104768 44198
rect 104716 44134 104768 44140
rect 104256 42220 104308 42226
rect 104256 42162 104308 42168
rect 104268 38010 104296 42162
rect 104348 38888 104400 38894
rect 104348 38830 104400 38836
rect 104256 38004 104308 38010
rect 104256 37946 104308 37952
rect 104268 37262 104296 37946
rect 104256 37256 104308 37262
rect 104256 37198 104308 37204
rect 104360 22778 104388 38830
rect 104728 37874 104756 44134
rect 104716 37868 104768 37874
rect 104716 37810 104768 37816
rect 104716 37324 104768 37330
rect 104716 37266 104768 37272
rect 104348 22772 104400 22778
rect 104348 22714 104400 22720
rect 104360 22273 104388 22714
rect 104346 22264 104402 22273
rect 104346 22199 104402 22208
rect 104728 10062 104756 37266
rect 104716 10056 104768 10062
rect 104716 9998 104768 10004
rect 90824 9988 90876 9994
rect 90824 9930 90876 9936
rect 103796 9988 103848 9994
rect 103796 9930 103848 9936
rect 90836 9897 90864 9930
rect 104820 9897 104848 49710
rect 105084 45484 105136 45490
rect 105084 45426 105136 45432
rect 105096 42362 105124 45426
rect 105176 45280 105228 45286
rect 105176 45222 105228 45228
rect 105084 42356 105136 42362
rect 105084 42298 105136 42304
rect 105188 37806 105216 45222
rect 105372 38894 105400 51206
rect 105360 38888 105412 38894
rect 105360 38830 105412 38836
rect 105832 38010 105860 58618
rect 105922 58236 106230 58245
rect 105922 58234 105928 58236
rect 105984 58234 106008 58236
rect 106064 58234 106088 58236
rect 106144 58234 106168 58236
rect 106224 58234 106230 58236
rect 105984 58182 105986 58234
rect 106166 58182 106168 58234
rect 105922 58180 105928 58182
rect 105984 58180 106008 58182
rect 106064 58180 106088 58182
rect 106144 58180 106168 58182
rect 106224 58180 106230 58182
rect 105922 58171 106230 58180
rect 106658 57692 106966 57701
rect 106658 57690 106664 57692
rect 106720 57690 106744 57692
rect 106800 57690 106824 57692
rect 106880 57690 106904 57692
rect 106960 57690 106966 57692
rect 106720 57638 106722 57690
rect 106902 57638 106904 57690
rect 106658 57636 106664 57638
rect 106720 57636 106744 57638
rect 106800 57636 106824 57638
rect 106880 57636 106904 57638
rect 106960 57636 106966 57638
rect 106658 57627 106966 57636
rect 105922 57148 106230 57157
rect 105922 57146 105928 57148
rect 105984 57146 106008 57148
rect 106064 57146 106088 57148
rect 106144 57146 106168 57148
rect 106224 57146 106230 57148
rect 105984 57094 105986 57146
rect 106166 57094 106168 57146
rect 105922 57092 105928 57094
rect 105984 57092 106008 57094
rect 106064 57092 106088 57094
rect 106144 57092 106168 57094
rect 106224 57092 106230 57094
rect 105922 57083 106230 57092
rect 106658 56604 106966 56613
rect 106658 56602 106664 56604
rect 106720 56602 106744 56604
rect 106800 56602 106824 56604
rect 106880 56602 106904 56604
rect 106960 56602 106966 56604
rect 106720 56550 106722 56602
rect 106902 56550 106904 56602
rect 106658 56548 106664 56550
rect 106720 56548 106744 56550
rect 106800 56548 106824 56550
rect 106880 56548 106904 56550
rect 106960 56548 106966 56550
rect 106658 56539 106966 56548
rect 105922 56060 106230 56069
rect 105922 56058 105928 56060
rect 105984 56058 106008 56060
rect 106064 56058 106088 56060
rect 106144 56058 106168 56060
rect 106224 56058 106230 56060
rect 105984 56006 105986 56058
rect 106166 56006 106168 56058
rect 105922 56004 105928 56006
rect 105984 56004 106008 56006
rect 106064 56004 106088 56006
rect 106144 56004 106168 56006
rect 106224 56004 106230 56006
rect 105922 55995 106230 56004
rect 106658 55516 106966 55525
rect 106658 55514 106664 55516
rect 106720 55514 106744 55516
rect 106800 55514 106824 55516
rect 106880 55514 106904 55516
rect 106960 55514 106966 55516
rect 106720 55462 106722 55514
rect 106902 55462 106904 55514
rect 106658 55460 106664 55462
rect 106720 55460 106744 55462
rect 106800 55460 106824 55462
rect 106880 55460 106904 55462
rect 106960 55460 106966 55462
rect 106658 55451 106966 55460
rect 105922 54972 106230 54981
rect 105922 54970 105928 54972
rect 105984 54970 106008 54972
rect 106064 54970 106088 54972
rect 106144 54970 106168 54972
rect 106224 54970 106230 54972
rect 105984 54918 105986 54970
rect 106166 54918 106168 54970
rect 105922 54916 105928 54918
rect 105984 54916 106008 54918
rect 106064 54916 106088 54918
rect 106144 54916 106168 54918
rect 106224 54916 106230 54918
rect 105922 54907 106230 54916
rect 106658 54428 106966 54437
rect 106658 54426 106664 54428
rect 106720 54426 106744 54428
rect 106800 54426 106824 54428
rect 106880 54426 106904 54428
rect 106960 54426 106966 54428
rect 106720 54374 106722 54426
rect 106902 54374 106904 54426
rect 106658 54372 106664 54374
rect 106720 54372 106744 54374
rect 106800 54372 106824 54374
rect 106880 54372 106904 54374
rect 106960 54372 106966 54374
rect 106658 54363 106966 54372
rect 105922 53884 106230 53893
rect 105922 53882 105928 53884
rect 105984 53882 106008 53884
rect 106064 53882 106088 53884
rect 106144 53882 106168 53884
rect 106224 53882 106230 53884
rect 105984 53830 105986 53882
rect 106166 53830 106168 53882
rect 105922 53828 105928 53830
rect 105984 53828 106008 53830
rect 106064 53828 106088 53830
rect 106144 53828 106168 53830
rect 106224 53828 106230 53830
rect 105922 53819 106230 53828
rect 106658 53340 106966 53349
rect 106658 53338 106664 53340
rect 106720 53338 106744 53340
rect 106800 53338 106824 53340
rect 106880 53338 106904 53340
rect 106960 53338 106966 53340
rect 106720 53286 106722 53338
rect 106902 53286 106904 53338
rect 106658 53284 106664 53286
rect 106720 53284 106744 53286
rect 106800 53284 106824 53286
rect 106880 53284 106904 53286
rect 106960 53284 106966 53286
rect 106658 53275 106966 53284
rect 105922 52796 106230 52805
rect 105922 52794 105928 52796
rect 105984 52794 106008 52796
rect 106064 52794 106088 52796
rect 106144 52794 106168 52796
rect 106224 52794 106230 52796
rect 105984 52742 105986 52794
rect 106166 52742 106168 52794
rect 105922 52740 105928 52742
rect 105984 52740 106008 52742
rect 106064 52740 106088 52742
rect 106144 52740 106168 52742
rect 106224 52740 106230 52742
rect 105922 52731 106230 52740
rect 106658 52252 106966 52261
rect 106658 52250 106664 52252
rect 106720 52250 106744 52252
rect 106800 52250 106824 52252
rect 106880 52250 106904 52252
rect 106960 52250 106966 52252
rect 106720 52198 106722 52250
rect 106902 52198 106904 52250
rect 106658 52196 106664 52198
rect 106720 52196 106744 52198
rect 106800 52196 106824 52198
rect 106880 52196 106904 52198
rect 106960 52196 106966 52198
rect 106658 52187 106966 52196
rect 105922 51708 106230 51717
rect 105922 51706 105928 51708
rect 105984 51706 106008 51708
rect 106064 51706 106088 51708
rect 106144 51706 106168 51708
rect 106224 51706 106230 51708
rect 105984 51654 105986 51706
rect 106166 51654 106168 51706
rect 105922 51652 105928 51654
rect 105984 51652 106008 51654
rect 106064 51652 106088 51654
rect 106144 51652 106168 51654
rect 106224 51652 106230 51654
rect 105922 51643 106230 51652
rect 108488 51400 108540 51406
rect 108488 51342 108540 51348
rect 108304 51264 108356 51270
rect 108304 51206 108356 51212
rect 106658 51164 106966 51173
rect 106658 51162 106664 51164
rect 106720 51162 106744 51164
rect 106800 51162 106824 51164
rect 106880 51162 106904 51164
rect 106960 51162 106966 51164
rect 106720 51110 106722 51162
rect 106902 51110 106904 51162
rect 106658 51108 106664 51110
rect 106720 51108 106744 51110
rect 106800 51108 106824 51110
rect 106880 51108 106904 51110
rect 106960 51108 106966 51110
rect 106658 51099 106966 51108
rect 105922 50620 106230 50629
rect 105922 50618 105928 50620
rect 105984 50618 106008 50620
rect 106064 50618 106088 50620
rect 106144 50618 106168 50620
rect 106224 50618 106230 50620
rect 105984 50566 105986 50618
rect 106166 50566 106168 50618
rect 105922 50564 105928 50566
rect 105984 50564 106008 50566
rect 106064 50564 106088 50566
rect 106144 50564 106168 50566
rect 106224 50564 106230 50566
rect 105922 50555 106230 50564
rect 106658 50076 106966 50085
rect 106658 50074 106664 50076
rect 106720 50074 106744 50076
rect 106800 50074 106824 50076
rect 106880 50074 106904 50076
rect 106960 50074 106966 50076
rect 106720 50022 106722 50074
rect 106902 50022 106904 50074
rect 106658 50020 106664 50022
rect 106720 50020 106744 50022
rect 106800 50020 106824 50022
rect 106880 50020 106904 50022
rect 106960 50020 106966 50022
rect 106658 50011 106966 50020
rect 105922 49532 106230 49541
rect 105922 49530 105928 49532
rect 105984 49530 106008 49532
rect 106064 49530 106088 49532
rect 106144 49530 106168 49532
rect 106224 49530 106230 49532
rect 105984 49478 105986 49530
rect 106166 49478 106168 49530
rect 105922 49476 105928 49478
rect 105984 49476 106008 49478
rect 106064 49476 106088 49478
rect 106144 49476 106168 49478
rect 106224 49476 106230 49478
rect 105922 49467 106230 49476
rect 106658 48988 106966 48997
rect 106658 48986 106664 48988
rect 106720 48986 106744 48988
rect 106800 48986 106824 48988
rect 106880 48986 106904 48988
rect 106960 48986 106966 48988
rect 106720 48934 106722 48986
rect 106902 48934 106904 48986
rect 106658 48932 106664 48934
rect 106720 48932 106744 48934
rect 106800 48932 106824 48934
rect 106880 48932 106904 48934
rect 106960 48932 106966 48934
rect 106658 48923 106966 48932
rect 105922 48444 106230 48453
rect 105922 48442 105928 48444
rect 105984 48442 106008 48444
rect 106064 48442 106088 48444
rect 106144 48442 106168 48444
rect 106224 48442 106230 48444
rect 105984 48390 105986 48442
rect 106166 48390 106168 48442
rect 105922 48388 105928 48390
rect 105984 48388 106008 48390
rect 106064 48388 106088 48390
rect 106144 48388 106168 48390
rect 106224 48388 106230 48390
rect 105922 48379 106230 48388
rect 106658 47900 106966 47909
rect 106658 47898 106664 47900
rect 106720 47898 106744 47900
rect 106800 47898 106824 47900
rect 106880 47898 106904 47900
rect 106960 47898 106966 47900
rect 106720 47846 106722 47898
rect 106902 47846 106904 47898
rect 106658 47844 106664 47846
rect 106720 47844 106744 47846
rect 106800 47844 106824 47846
rect 106880 47844 106904 47846
rect 106960 47844 106966 47846
rect 106658 47835 106966 47844
rect 105922 47356 106230 47365
rect 105922 47354 105928 47356
rect 105984 47354 106008 47356
rect 106064 47354 106088 47356
rect 106144 47354 106168 47356
rect 106224 47354 106230 47356
rect 105984 47302 105986 47354
rect 106166 47302 106168 47354
rect 105922 47300 105928 47302
rect 105984 47300 106008 47302
rect 106064 47300 106088 47302
rect 106144 47300 106168 47302
rect 106224 47300 106230 47302
rect 105922 47291 106230 47300
rect 106658 46812 106966 46821
rect 106658 46810 106664 46812
rect 106720 46810 106744 46812
rect 106800 46810 106824 46812
rect 106880 46810 106904 46812
rect 106960 46810 106966 46812
rect 106720 46758 106722 46810
rect 106902 46758 106904 46810
rect 106658 46756 106664 46758
rect 106720 46756 106744 46758
rect 106800 46756 106824 46758
rect 106880 46756 106904 46758
rect 106960 46756 106966 46758
rect 106658 46747 106966 46756
rect 105922 46268 106230 46277
rect 105922 46266 105928 46268
rect 105984 46266 106008 46268
rect 106064 46266 106088 46268
rect 106144 46266 106168 46268
rect 106224 46266 106230 46268
rect 105984 46214 105986 46266
rect 106166 46214 106168 46266
rect 105922 46212 105928 46214
rect 105984 46212 106008 46214
rect 106064 46212 106088 46214
rect 106144 46212 106168 46214
rect 106224 46212 106230 46214
rect 105922 46203 106230 46212
rect 106658 45724 106966 45733
rect 106658 45722 106664 45724
rect 106720 45722 106744 45724
rect 106800 45722 106824 45724
rect 106880 45722 106904 45724
rect 106960 45722 106966 45724
rect 106720 45670 106722 45722
rect 106902 45670 106904 45722
rect 106658 45668 106664 45670
rect 106720 45668 106744 45670
rect 106800 45668 106824 45670
rect 106880 45668 106904 45670
rect 106960 45668 106966 45670
rect 106658 45659 106966 45668
rect 105922 45180 106230 45189
rect 105922 45178 105928 45180
rect 105984 45178 106008 45180
rect 106064 45178 106088 45180
rect 106144 45178 106168 45180
rect 106224 45178 106230 45180
rect 105984 45126 105986 45178
rect 106166 45126 106168 45178
rect 105922 45124 105928 45126
rect 105984 45124 106008 45126
rect 106064 45124 106088 45126
rect 106144 45124 106168 45126
rect 106224 45124 106230 45126
rect 105922 45115 106230 45124
rect 108316 44878 108344 51206
rect 108500 51105 108528 51342
rect 108486 51096 108542 51105
rect 108486 51031 108542 51040
rect 108304 44872 108356 44878
rect 108304 44814 108356 44820
rect 106658 44636 106966 44645
rect 106658 44634 106664 44636
rect 106720 44634 106744 44636
rect 106800 44634 106824 44636
rect 106880 44634 106904 44636
rect 106960 44634 106966 44636
rect 106720 44582 106722 44634
rect 106902 44582 106904 44634
rect 106658 44580 106664 44582
rect 106720 44580 106744 44582
rect 106800 44580 106824 44582
rect 106880 44580 106904 44582
rect 106960 44580 106966 44582
rect 106658 44571 106966 44580
rect 105922 44092 106230 44101
rect 105922 44090 105928 44092
rect 105984 44090 106008 44092
rect 106064 44090 106088 44092
rect 106144 44090 106168 44092
rect 106224 44090 106230 44092
rect 105984 44038 105986 44090
rect 106166 44038 106168 44090
rect 105922 44036 105928 44038
rect 105984 44036 106008 44038
rect 106064 44036 106088 44038
rect 106144 44036 106168 44038
rect 106224 44036 106230 44038
rect 105922 44027 106230 44036
rect 106658 43548 106966 43557
rect 106658 43546 106664 43548
rect 106720 43546 106744 43548
rect 106800 43546 106824 43548
rect 106880 43546 106904 43548
rect 106960 43546 106966 43548
rect 106720 43494 106722 43546
rect 106902 43494 106904 43546
rect 106658 43492 106664 43494
rect 106720 43492 106744 43494
rect 106800 43492 106824 43494
rect 106880 43492 106904 43494
rect 106960 43492 106966 43494
rect 106658 43483 106966 43492
rect 105922 43004 106230 43013
rect 105922 43002 105928 43004
rect 105984 43002 106008 43004
rect 106064 43002 106088 43004
rect 106144 43002 106168 43004
rect 106224 43002 106230 43004
rect 105984 42950 105986 43002
rect 106166 42950 106168 43002
rect 105922 42948 105928 42950
rect 105984 42948 106008 42950
rect 106064 42948 106088 42950
rect 106144 42948 106168 42950
rect 106224 42948 106230 42950
rect 105922 42939 106230 42948
rect 106658 42460 106966 42469
rect 106658 42458 106664 42460
rect 106720 42458 106744 42460
rect 106800 42458 106824 42460
rect 106880 42458 106904 42460
rect 106960 42458 106966 42460
rect 106720 42406 106722 42458
rect 106902 42406 106904 42458
rect 106658 42404 106664 42406
rect 106720 42404 106744 42406
rect 106800 42404 106824 42406
rect 106880 42404 106904 42406
rect 106960 42404 106966 42406
rect 106658 42395 106966 42404
rect 105922 41916 106230 41925
rect 105922 41914 105928 41916
rect 105984 41914 106008 41916
rect 106064 41914 106088 41916
rect 106144 41914 106168 41916
rect 106224 41914 106230 41916
rect 105984 41862 105986 41914
rect 106166 41862 106168 41914
rect 105922 41860 105928 41862
rect 105984 41860 106008 41862
rect 106064 41860 106088 41862
rect 106144 41860 106168 41862
rect 106224 41860 106230 41862
rect 105922 41851 106230 41860
rect 106658 41372 106966 41381
rect 106658 41370 106664 41372
rect 106720 41370 106744 41372
rect 106800 41370 106824 41372
rect 106880 41370 106904 41372
rect 106960 41370 106966 41372
rect 106720 41318 106722 41370
rect 106902 41318 106904 41370
rect 106658 41316 106664 41318
rect 106720 41316 106744 41318
rect 106800 41316 106824 41318
rect 106880 41316 106904 41318
rect 106960 41316 106966 41318
rect 106658 41307 106966 41316
rect 105922 40828 106230 40837
rect 105922 40826 105928 40828
rect 105984 40826 106008 40828
rect 106064 40826 106088 40828
rect 106144 40826 106168 40828
rect 106224 40826 106230 40828
rect 105984 40774 105986 40826
rect 106166 40774 106168 40826
rect 105922 40772 105928 40774
rect 105984 40772 106008 40774
rect 106064 40772 106088 40774
rect 106144 40772 106168 40774
rect 106224 40772 106230 40774
rect 105922 40763 106230 40772
rect 106658 40284 106966 40293
rect 106658 40282 106664 40284
rect 106720 40282 106744 40284
rect 106800 40282 106824 40284
rect 106880 40282 106904 40284
rect 106960 40282 106966 40284
rect 106720 40230 106722 40282
rect 106902 40230 106904 40282
rect 106658 40228 106664 40230
rect 106720 40228 106744 40230
rect 106800 40228 106824 40230
rect 106880 40228 106904 40230
rect 106960 40228 106966 40230
rect 106658 40219 106966 40228
rect 105922 39740 106230 39749
rect 105922 39738 105928 39740
rect 105984 39738 106008 39740
rect 106064 39738 106088 39740
rect 106144 39738 106168 39740
rect 106224 39738 106230 39740
rect 105984 39686 105986 39738
rect 106166 39686 106168 39738
rect 105922 39684 105928 39686
rect 105984 39684 106008 39686
rect 106064 39684 106088 39686
rect 106144 39684 106168 39686
rect 106224 39684 106230 39686
rect 105922 39675 106230 39684
rect 106658 39196 106966 39205
rect 106658 39194 106664 39196
rect 106720 39194 106744 39196
rect 106800 39194 106824 39196
rect 106880 39194 106904 39196
rect 106960 39194 106966 39196
rect 106720 39142 106722 39194
rect 106902 39142 106904 39194
rect 106658 39140 106664 39142
rect 106720 39140 106744 39142
rect 106800 39140 106824 39142
rect 106880 39140 106904 39142
rect 106960 39140 106966 39142
rect 106658 39131 106966 39140
rect 105922 38652 106230 38661
rect 105922 38650 105928 38652
rect 105984 38650 106008 38652
rect 106064 38650 106088 38652
rect 106144 38650 106168 38652
rect 106224 38650 106230 38652
rect 105984 38598 105986 38650
rect 106166 38598 106168 38650
rect 105922 38596 105928 38598
rect 105984 38596 106008 38598
rect 106064 38596 106088 38598
rect 106144 38596 106168 38598
rect 106224 38596 106230 38598
rect 105922 38587 106230 38596
rect 106658 38108 106966 38117
rect 106658 38106 106664 38108
rect 106720 38106 106744 38108
rect 106800 38106 106824 38108
rect 106880 38106 106904 38108
rect 106960 38106 106966 38108
rect 106720 38054 106722 38106
rect 106902 38054 106904 38106
rect 106658 38052 106664 38054
rect 106720 38052 106744 38054
rect 106800 38052 106824 38054
rect 106880 38052 106904 38054
rect 106960 38052 106966 38054
rect 106658 38043 106966 38052
rect 105820 38004 105872 38010
rect 105820 37946 105872 37952
rect 105176 37800 105228 37806
rect 105176 37742 105228 37748
rect 105922 37564 106230 37573
rect 105922 37562 105928 37564
rect 105984 37562 106008 37564
rect 106064 37562 106088 37564
rect 106144 37562 106168 37564
rect 106224 37562 106230 37564
rect 105984 37510 105986 37562
rect 106166 37510 106168 37562
rect 105922 37508 105928 37510
rect 105984 37508 106008 37510
rect 106064 37508 106088 37510
rect 106144 37508 106168 37510
rect 106224 37508 106230 37510
rect 105922 37499 106230 37508
rect 106658 37020 106966 37029
rect 106658 37018 106664 37020
rect 106720 37018 106744 37020
rect 106800 37018 106824 37020
rect 106880 37018 106904 37020
rect 106960 37018 106966 37020
rect 106720 36966 106722 37018
rect 106902 36966 106904 37018
rect 106658 36964 106664 36966
rect 106720 36964 106744 36966
rect 106800 36964 106824 36966
rect 106880 36964 106904 36966
rect 106960 36964 106966 36966
rect 106658 36955 106966 36964
rect 105922 36476 106230 36485
rect 105922 36474 105928 36476
rect 105984 36474 106008 36476
rect 106064 36474 106088 36476
rect 106144 36474 106168 36476
rect 106224 36474 106230 36476
rect 105984 36422 105986 36474
rect 106166 36422 106168 36474
rect 105922 36420 105928 36422
rect 105984 36420 106008 36422
rect 106064 36420 106088 36422
rect 106144 36420 106168 36422
rect 106224 36420 106230 36422
rect 105922 36411 106230 36420
rect 106658 35932 106966 35941
rect 106658 35930 106664 35932
rect 106720 35930 106744 35932
rect 106800 35930 106824 35932
rect 106880 35930 106904 35932
rect 106960 35930 106966 35932
rect 106720 35878 106722 35930
rect 106902 35878 106904 35930
rect 106658 35876 106664 35878
rect 106720 35876 106744 35878
rect 106800 35876 106824 35878
rect 106880 35876 106904 35878
rect 106960 35876 106966 35878
rect 106658 35867 106966 35876
rect 105922 35388 106230 35397
rect 105922 35386 105928 35388
rect 105984 35386 106008 35388
rect 106064 35386 106088 35388
rect 106144 35386 106168 35388
rect 106224 35386 106230 35388
rect 105984 35334 105986 35386
rect 106166 35334 106168 35386
rect 105922 35332 105928 35334
rect 105984 35332 106008 35334
rect 106064 35332 106088 35334
rect 106144 35332 106168 35334
rect 106224 35332 106230 35334
rect 105922 35323 106230 35332
rect 106658 34844 106966 34853
rect 106658 34842 106664 34844
rect 106720 34842 106744 34844
rect 106800 34842 106824 34844
rect 106880 34842 106904 34844
rect 106960 34842 106966 34844
rect 106720 34790 106722 34842
rect 106902 34790 106904 34842
rect 106658 34788 106664 34790
rect 106720 34788 106744 34790
rect 106800 34788 106824 34790
rect 106880 34788 106904 34790
rect 106960 34788 106966 34790
rect 106658 34779 106966 34788
rect 105922 34300 106230 34309
rect 105922 34298 105928 34300
rect 105984 34298 106008 34300
rect 106064 34298 106088 34300
rect 106144 34298 106168 34300
rect 106224 34298 106230 34300
rect 105984 34246 105986 34298
rect 106166 34246 106168 34298
rect 105922 34244 105928 34246
rect 105984 34244 106008 34246
rect 106064 34244 106088 34246
rect 106144 34244 106168 34246
rect 106224 34244 106230 34246
rect 105922 34235 106230 34244
rect 106658 33756 106966 33765
rect 106658 33754 106664 33756
rect 106720 33754 106744 33756
rect 106800 33754 106824 33756
rect 106880 33754 106904 33756
rect 106960 33754 106966 33756
rect 106720 33702 106722 33754
rect 106902 33702 106904 33754
rect 106658 33700 106664 33702
rect 106720 33700 106744 33702
rect 106800 33700 106824 33702
rect 106880 33700 106904 33702
rect 106960 33700 106966 33702
rect 106658 33691 106966 33700
rect 105922 33212 106230 33221
rect 105922 33210 105928 33212
rect 105984 33210 106008 33212
rect 106064 33210 106088 33212
rect 106144 33210 106168 33212
rect 106224 33210 106230 33212
rect 105984 33158 105986 33210
rect 106166 33158 106168 33210
rect 105922 33156 105928 33158
rect 105984 33156 106008 33158
rect 106064 33156 106088 33158
rect 106144 33156 106168 33158
rect 106224 33156 106230 33158
rect 105922 33147 106230 33156
rect 106658 32668 106966 32677
rect 106658 32666 106664 32668
rect 106720 32666 106744 32668
rect 106800 32666 106824 32668
rect 106880 32666 106904 32668
rect 106960 32666 106966 32668
rect 106720 32614 106722 32666
rect 106902 32614 106904 32666
rect 106658 32612 106664 32614
rect 106720 32612 106744 32614
rect 106800 32612 106824 32614
rect 106880 32612 106904 32614
rect 106960 32612 106966 32614
rect 106658 32603 106966 32612
rect 105922 32124 106230 32133
rect 105922 32122 105928 32124
rect 105984 32122 106008 32124
rect 106064 32122 106088 32124
rect 106144 32122 106168 32124
rect 106224 32122 106230 32124
rect 105984 32070 105986 32122
rect 106166 32070 106168 32122
rect 105922 32068 105928 32070
rect 105984 32068 106008 32070
rect 106064 32068 106088 32070
rect 106144 32068 106168 32070
rect 106224 32068 106230 32070
rect 105922 32059 106230 32068
rect 106658 31580 106966 31589
rect 106658 31578 106664 31580
rect 106720 31578 106744 31580
rect 106800 31578 106824 31580
rect 106880 31578 106904 31580
rect 106960 31578 106966 31580
rect 106720 31526 106722 31578
rect 106902 31526 106904 31578
rect 106658 31524 106664 31526
rect 106720 31524 106744 31526
rect 106800 31524 106824 31526
rect 106880 31524 106904 31526
rect 106960 31524 106966 31526
rect 106658 31515 106966 31524
rect 105922 31036 106230 31045
rect 105922 31034 105928 31036
rect 105984 31034 106008 31036
rect 106064 31034 106088 31036
rect 106144 31034 106168 31036
rect 106224 31034 106230 31036
rect 105984 30982 105986 31034
rect 106166 30982 106168 31034
rect 105922 30980 105928 30982
rect 105984 30980 106008 30982
rect 106064 30980 106088 30982
rect 106144 30980 106168 30982
rect 106224 30980 106230 30982
rect 105922 30971 106230 30980
rect 106658 30492 106966 30501
rect 106658 30490 106664 30492
rect 106720 30490 106744 30492
rect 106800 30490 106824 30492
rect 106880 30490 106904 30492
rect 106960 30490 106966 30492
rect 106720 30438 106722 30490
rect 106902 30438 106904 30490
rect 106658 30436 106664 30438
rect 106720 30436 106744 30438
rect 106800 30436 106824 30438
rect 106880 30436 106904 30438
rect 106960 30436 106966 30438
rect 106658 30427 106966 30436
rect 105922 29948 106230 29957
rect 105922 29946 105928 29948
rect 105984 29946 106008 29948
rect 106064 29946 106088 29948
rect 106144 29946 106168 29948
rect 106224 29946 106230 29948
rect 105984 29894 105986 29946
rect 106166 29894 106168 29946
rect 105922 29892 105928 29894
rect 105984 29892 106008 29894
rect 106064 29892 106088 29894
rect 106144 29892 106168 29894
rect 106224 29892 106230 29894
rect 105922 29883 106230 29892
rect 106658 29404 106966 29413
rect 106658 29402 106664 29404
rect 106720 29402 106744 29404
rect 106800 29402 106824 29404
rect 106880 29402 106904 29404
rect 106960 29402 106966 29404
rect 106720 29350 106722 29402
rect 106902 29350 106904 29402
rect 106658 29348 106664 29350
rect 106720 29348 106744 29350
rect 106800 29348 106824 29350
rect 106880 29348 106904 29350
rect 106960 29348 106966 29350
rect 106658 29339 106966 29348
rect 105922 28860 106230 28869
rect 105922 28858 105928 28860
rect 105984 28858 106008 28860
rect 106064 28858 106088 28860
rect 106144 28858 106168 28860
rect 106224 28858 106230 28860
rect 105984 28806 105986 28858
rect 106166 28806 106168 28858
rect 105922 28804 105928 28806
rect 105984 28804 106008 28806
rect 106064 28804 106088 28806
rect 106144 28804 106168 28806
rect 106224 28804 106230 28806
rect 105922 28795 106230 28804
rect 106658 28316 106966 28325
rect 106658 28314 106664 28316
rect 106720 28314 106744 28316
rect 106800 28314 106824 28316
rect 106880 28314 106904 28316
rect 106960 28314 106966 28316
rect 106720 28262 106722 28314
rect 106902 28262 106904 28314
rect 106658 28260 106664 28262
rect 106720 28260 106744 28262
rect 106800 28260 106824 28262
rect 106880 28260 106904 28262
rect 106960 28260 106966 28262
rect 106658 28251 106966 28260
rect 105922 27772 106230 27781
rect 105922 27770 105928 27772
rect 105984 27770 106008 27772
rect 106064 27770 106088 27772
rect 106144 27770 106168 27772
rect 106224 27770 106230 27772
rect 105984 27718 105986 27770
rect 106166 27718 106168 27770
rect 105922 27716 105928 27718
rect 105984 27716 106008 27718
rect 106064 27716 106088 27718
rect 106144 27716 106168 27718
rect 106224 27716 106230 27718
rect 105922 27707 106230 27716
rect 106658 27228 106966 27237
rect 106658 27226 106664 27228
rect 106720 27226 106744 27228
rect 106800 27226 106824 27228
rect 106880 27226 106904 27228
rect 106960 27226 106966 27228
rect 106720 27174 106722 27226
rect 106902 27174 106904 27226
rect 106658 27172 106664 27174
rect 106720 27172 106744 27174
rect 106800 27172 106824 27174
rect 106880 27172 106904 27174
rect 106960 27172 106966 27174
rect 106658 27163 106966 27172
rect 105922 26684 106230 26693
rect 105922 26682 105928 26684
rect 105984 26682 106008 26684
rect 106064 26682 106088 26684
rect 106144 26682 106168 26684
rect 106224 26682 106230 26684
rect 105984 26630 105986 26682
rect 106166 26630 106168 26682
rect 105922 26628 105928 26630
rect 105984 26628 106008 26630
rect 106064 26628 106088 26630
rect 106144 26628 106168 26630
rect 106224 26628 106230 26630
rect 105922 26619 106230 26628
rect 106658 26140 106966 26149
rect 106658 26138 106664 26140
rect 106720 26138 106744 26140
rect 106800 26138 106824 26140
rect 106880 26138 106904 26140
rect 106960 26138 106966 26140
rect 106720 26086 106722 26138
rect 106902 26086 106904 26138
rect 106658 26084 106664 26086
rect 106720 26084 106744 26086
rect 106800 26084 106824 26086
rect 106880 26084 106904 26086
rect 106960 26084 106966 26086
rect 106658 26075 106966 26084
rect 105922 25596 106230 25605
rect 105922 25594 105928 25596
rect 105984 25594 106008 25596
rect 106064 25594 106088 25596
rect 106144 25594 106168 25596
rect 106224 25594 106230 25596
rect 105984 25542 105986 25594
rect 106166 25542 106168 25594
rect 105922 25540 105928 25542
rect 105984 25540 106008 25542
rect 106064 25540 106088 25542
rect 106144 25540 106168 25542
rect 106224 25540 106230 25542
rect 105922 25531 106230 25540
rect 106658 25052 106966 25061
rect 106658 25050 106664 25052
rect 106720 25050 106744 25052
rect 106800 25050 106824 25052
rect 106880 25050 106904 25052
rect 106960 25050 106966 25052
rect 106720 24998 106722 25050
rect 106902 24998 106904 25050
rect 106658 24996 106664 24998
rect 106720 24996 106744 24998
rect 106800 24996 106824 24998
rect 106880 24996 106904 24998
rect 106960 24996 106966 24998
rect 106658 24987 106966 24996
rect 105922 24508 106230 24517
rect 105922 24506 105928 24508
rect 105984 24506 106008 24508
rect 106064 24506 106088 24508
rect 106144 24506 106168 24508
rect 106224 24506 106230 24508
rect 105984 24454 105986 24506
rect 106166 24454 106168 24506
rect 105922 24452 105928 24454
rect 105984 24452 106008 24454
rect 106064 24452 106088 24454
rect 106144 24452 106168 24454
rect 106224 24452 106230 24454
rect 105922 24443 106230 24452
rect 106658 23964 106966 23973
rect 106658 23962 106664 23964
rect 106720 23962 106744 23964
rect 106800 23962 106824 23964
rect 106880 23962 106904 23964
rect 106960 23962 106966 23964
rect 106720 23910 106722 23962
rect 106902 23910 106904 23962
rect 106658 23908 106664 23910
rect 106720 23908 106744 23910
rect 106800 23908 106824 23910
rect 106880 23908 106904 23910
rect 106960 23908 106966 23910
rect 106658 23899 106966 23908
rect 105922 23420 106230 23429
rect 105922 23418 105928 23420
rect 105984 23418 106008 23420
rect 106064 23418 106088 23420
rect 106144 23418 106168 23420
rect 106224 23418 106230 23420
rect 105984 23366 105986 23418
rect 106166 23366 106168 23418
rect 105922 23364 105928 23366
rect 105984 23364 106008 23366
rect 106064 23364 106088 23366
rect 106144 23364 106168 23366
rect 106224 23364 106230 23366
rect 105922 23355 106230 23364
rect 106658 22876 106966 22885
rect 106658 22874 106664 22876
rect 106720 22874 106744 22876
rect 106800 22874 106824 22876
rect 106880 22874 106904 22876
rect 106960 22874 106966 22876
rect 106720 22822 106722 22874
rect 106902 22822 106904 22874
rect 106658 22820 106664 22822
rect 106720 22820 106744 22822
rect 106800 22820 106824 22822
rect 106880 22820 106904 22822
rect 106960 22820 106966 22822
rect 106658 22811 106966 22820
rect 105922 22332 106230 22341
rect 105922 22330 105928 22332
rect 105984 22330 106008 22332
rect 106064 22330 106088 22332
rect 106144 22330 106168 22332
rect 106224 22330 106230 22332
rect 105984 22278 105986 22330
rect 106166 22278 106168 22330
rect 105922 22276 105928 22278
rect 105984 22276 106008 22278
rect 106064 22276 106088 22278
rect 106144 22276 106168 22278
rect 106224 22276 106230 22278
rect 105922 22267 106230 22276
rect 106658 21788 106966 21797
rect 106658 21786 106664 21788
rect 106720 21786 106744 21788
rect 106800 21786 106824 21788
rect 106880 21786 106904 21788
rect 106960 21786 106966 21788
rect 106720 21734 106722 21786
rect 106902 21734 106904 21786
rect 106658 21732 106664 21734
rect 106720 21732 106744 21734
rect 106800 21732 106824 21734
rect 106880 21732 106904 21734
rect 106960 21732 106966 21734
rect 106658 21723 106966 21732
rect 105922 21244 106230 21253
rect 105922 21242 105928 21244
rect 105984 21242 106008 21244
rect 106064 21242 106088 21244
rect 106144 21242 106168 21244
rect 106224 21242 106230 21244
rect 105984 21190 105986 21242
rect 106166 21190 106168 21242
rect 105922 21188 105928 21190
rect 105984 21188 106008 21190
rect 106064 21188 106088 21190
rect 106144 21188 106168 21190
rect 106224 21188 106230 21190
rect 105922 21179 106230 21188
rect 106658 20700 106966 20709
rect 106658 20698 106664 20700
rect 106720 20698 106744 20700
rect 106800 20698 106824 20700
rect 106880 20698 106904 20700
rect 106960 20698 106966 20700
rect 106720 20646 106722 20698
rect 106902 20646 106904 20698
rect 106658 20644 106664 20646
rect 106720 20644 106744 20646
rect 106800 20644 106824 20646
rect 106880 20644 106904 20646
rect 106960 20644 106966 20646
rect 106658 20635 106966 20644
rect 105922 20156 106230 20165
rect 105922 20154 105928 20156
rect 105984 20154 106008 20156
rect 106064 20154 106088 20156
rect 106144 20154 106168 20156
rect 106224 20154 106230 20156
rect 105984 20102 105986 20154
rect 106166 20102 106168 20154
rect 105922 20100 105928 20102
rect 105984 20100 106008 20102
rect 106064 20100 106088 20102
rect 106144 20100 106168 20102
rect 106224 20100 106230 20102
rect 105922 20091 106230 20100
rect 106658 19612 106966 19621
rect 106658 19610 106664 19612
rect 106720 19610 106744 19612
rect 106800 19610 106824 19612
rect 106880 19610 106904 19612
rect 106960 19610 106966 19612
rect 106720 19558 106722 19610
rect 106902 19558 106904 19610
rect 106658 19556 106664 19558
rect 106720 19556 106744 19558
rect 106800 19556 106824 19558
rect 106880 19556 106904 19558
rect 106960 19556 106966 19558
rect 106658 19547 106966 19556
rect 105922 19068 106230 19077
rect 105922 19066 105928 19068
rect 105984 19066 106008 19068
rect 106064 19066 106088 19068
rect 106144 19066 106168 19068
rect 106224 19066 106230 19068
rect 105984 19014 105986 19066
rect 106166 19014 106168 19066
rect 105922 19012 105928 19014
rect 105984 19012 106008 19014
rect 106064 19012 106088 19014
rect 106144 19012 106168 19014
rect 106224 19012 106230 19014
rect 105922 19003 106230 19012
rect 106658 18524 106966 18533
rect 106658 18522 106664 18524
rect 106720 18522 106744 18524
rect 106800 18522 106824 18524
rect 106880 18522 106904 18524
rect 106960 18522 106966 18524
rect 106720 18470 106722 18522
rect 106902 18470 106904 18522
rect 106658 18468 106664 18470
rect 106720 18468 106744 18470
rect 106800 18468 106824 18470
rect 106880 18468 106904 18470
rect 106960 18468 106966 18470
rect 106658 18459 106966 18468
rect 105922 17980 106230 17989
rect 105922 17978 105928 17980
rect 105984 17978 106008 17980
rect 106064 17978 106088 17980
rect 106144 17978 106168 17980
rect 106224 17978 106230 17980
rect 105984 17926 105986 17978
rect 106166 17926 106168 17978
rect 105922 17924 105928 17926
rect 105984 17924 106008 17926
rect 106064 17924 106088 17926
rect 106144 17924 106168 17926
rect 106224 17924 106230 17926
rect 105922 17915 106230 17924
rect 106658 17436 106966 17445
rect 106658 17434 106664 17436
rect 106720 17434 106744 17436
rect 106800 17434 106824 17436
rect 106880 17434 106904 17436
rect 106960 17434 106966 17436
rect 106720 17382 106722 17434
rect 106902 17382 106904 17434
rect 106658 17380 106664 17382
rect 106720 17380 106744 17382
rect 106800 17380 106824 17382
rect 106880 17380 106904 17382
rect 106960 17380 106966 17382
rect 106658 17371 106966 17380
rect 105922 16892 106230 16901
rect 105922 16890 105928 16892
rect 105984 16890 106008 16892
rect 106064 16890 106088 16892
rect 106144 16890 106168 16892
rect 106224 16890 106230 16892
rect 105984 16838 105986 16890
rect 106166 16838 106168 16890
rect 105922 16836 105928 16838
rect 105984 16836 106008 16838
rect 106064 16836 106088 16838
rect 106144 16836 106168 16838
rect 106224 16836 106230 16838
rect 105922 16827 106230 16836
rect 106658 16348 106966 16357
rect 106658 16346 106664 16348
rect 106720 16346 106744 16348
rect 106800 16346 106824 16348
rect 106880 16346 106904 16348
rect 106960 16346 106966 16348
rect 106720 16294 106722 16346
rect 106902 16294 106904 16346
rect 106658 16292 106664 16294
rect 106720 16292 106744 16294
rect 106800 16292 106824 16294
rect 106880 16292 106904 16294
rect 106960 16292 106966 16294
rect 106658 16283 106966 16292
rect 105922 15804 106230 15813
rect 105922 15802 105928 15804
rect 105984 15802 106008 15804
rect 106064 15802 106088 15804
rect 106144 15802 106168 15804
rect 106224 15802 106230 15804
rect 105984 15750 105986 15802
rect 106166 15750 106168 15802
rect 105922 15748 105928 15750
rect 105984 15748 106008 15750
rect 106064 15748 106088 15750
rect 106144 15748 106168 15750
rect 106224 15748 106230 15750
rect 105922 15739 106230 15748
rect 106658 15260 106966 15269
rect 106658 15258 106664 15260
rect 106720 15258 106744 15260
rect 106800 15258 106824 15260
rect 106880 15258 106904 15260
rect 106960 15258 106966 15260
rect 106720 15206 106722 15258
rect 106902 15206 106904 15258
rect 106658 15204 106664 15206
rect 106720 15204 106744 15206
rect 106800 15204 106824 15206
rect 106880 15204 106904 15206
rect 106960 15204 106966 15206
rect 106658 15195 106966 15204
rect 105922 14716 106230 14725
rect 105922 14714 105928 14716
rect 105984 14714 106008 14716
rect 106064 14714 106088 14716
rect 106144 14714 106168 14716
rect 106224 14714 106230 14716
rect 105984 14662 105986 14714
rect 106166 14662 106168 14714
rect 105922 14660 105928 14662
rect 105984 14660 106008 14662
rect 106064 14660 106088 14662
rect 106144 14660 106168 14662
rect 106224 14660 106230 14662
rect 105922 14651 106230 14660
rect 106658 14172 106966 14181
rect 106658 14170 106664 14172
rect 106720 14170 106744 14172
rect 106800 14170 106824 14172
rect 106880 14170 106904 14172
rect 106960 14170 106966 14172
rect 106720 14118 106722 14170
rect 106902 14118 106904 14170
rect 106658 14116 106664 14118
rect 106720 14116 106744 14118
rect 106800 14116 106824 14118
rect 106880 14116 106904 14118
rect 106960 14116 106966 14118
rect 106658 14107 106966 14116
rect 105922 13628 106230 13637
rect 105922 13626 105928 13628
rect 105984 13626 106008 13628
rect 106064 13626 106088 13628
rect 106144 13626 106168 13628
rect 106224 13626 106230 13628
rect 105984 13574 105986 13626
rect 106166 13574 106168 13626
rect 105922 13572 105928 13574
rect 105984 13572 106008 13574
rect 106064 13572 106088 13574
rect 106144 13572 106168 13574
rect 106224 13572 106230 13574
rect 105922 13563 106230 13572
rect 106658 13084 106966 13093
rect 106658 13082 106664 13084
rect 106720 13082 106744 13084
rect 106800 13082 106824 13084
rect 106880 13082 106904 13084
rect 106960 13082 106966 13084
rect 106720 13030 106722 13082
rect 106902 13030 106904 13082
rect 106658 13028 106664 13030
rect 106720 13028 106744 13030
rect 106800 13028 106824 13030
rect 106880 13028 106904 13030
rect 106960 13028 106966 13030
rect 106658 13019 106966 13028
rect 105922 12540 106230 12549
rect 105922 12538 105928 12540
rect 105984 12538 106008 12540
rect 106064 12538 106088 12540
rect 106144 12538 106168 12540
rect 106224 12538 106230 12540
rect 105984 12486 105986 12538
rect 106166 12486 106168 12538
rect 105922 12484 105928 12486
rect 105984 12484 106008 12486
rect 106064 12484 106088 12486
rect 106144 12484 106168 12486
rect 106224 12484 106230 12486
rect 105922 12475 106230 12484
rect 106658 11996 106966 12005
rect 106658 11994 106664 11996
rect 106720 11994 106744 11996
rect 106800 11994 106824 11996
rect 106880 11994 106904 11996
rect 106960 11994 106966 11996
rect 106720 11942 106722 11994
rect 106902 11942 106904 11994
rect 106658 11940 106664 11942
rect 106720 11940 106744 11942
rect 106800 11940 106824 11942
rect 106880 11940 106904 11942
rect 106960 11940 106966 11942
rect 106658 11931 106966 11940
rect 105922 11452 106230 11461
rect 105922 11450 105928 11452
rect 105984 11450 106008 11452
rect 106064 11450 106088 11452
rect 106144 11450 106168 11452
rect 106224 11450 106230 11452
rect 105984 11398 105986 11450
rect 106166 11398 106168 11450
rect 105922 11396 105928 11398
rect 105984 11396 106008 11398
rect 106064 11396 106088 11398
rect 106144 11396 106168 11398
rect 106224 11396 106230 11398
rect 105922 11387 106230 11396
rect 106658 10908 106966 10917
rect 106658 10906 106664 10908
rect 106720 10906 106744 10908
rect 106800 10906 106824 10908
rect 106880 10906 106904 10908
rect 106960 10906 106966 10908
rect 106720 10854 106722 10906
rect 106902 10854 106904 10906
rect 106658 10852 106664 10854
rect 106720 10852 106744 10854
rect 106800 10852 106824 10854
rect 106880 10852 106904 10854
rect 106960 10852 106966 10854
rect 106658 10843 106966 10852
rect 105922 10364 106230 10373
rect 105922 10362 105928 10364
rect 105984 10362 106008 10364
rect 106064 10362 106088 10364
rect 106144 10362 106168 10364
rect 106224 10362 106230 10364
rect 105984 10310 105986 10362
rect 106166 10310 106168 10362
rect 105922 10308 105928 10310
rect 105984 10308 106008 10310
rect 106064 10308 106088 10310
rect 106144 10308 106168 10310
rect 106224 10308 106230 10310
rect 105922 10299 106230 10308
rect 90822 9888 90878 9897
rect 90822 9823 90878 9832
rect 104806 9888 104862 9897
rect 104806 9823 104862 9832
rect 106658 9820 106966 9829
rect 106658 9818 106664 9820
rect 106720 9818 106744 9820
rect 106800 9818 106824 9820
rect 106880 9818 106904 9820
rect 106960 9818 106966 9820
rect 106720 9766 106722 9818
rect 106902 9766 106904 9818
rect 106658 9764 106664 9766
rect 106720 9764 106744 9766
rect 106800 9764 106824 9766
rect 106880 9764 106904 9766
rect 106960 9764 106966 9766
rect 90730 9752 90786 9761
rect 106658 9755 106966 9764
rect 90730 9687 90786 9696
rect 23478 8256 23534 8265
rect 23478 8191 23534 8200
rect 24766 8256 24822 8265
rect 24766 8191 24822 8200
rect 25870 8256 25926 8265
rect 25870 8191 25926 8200
rect 27158 8256 27214 8265
rect 27158 8191 27214 8200
rect 28446 8256 28502 8265
rect 28446 8191 28502 8200
rect 29274 8256 29330 8265
rect 29274 8191 29330 8200
rect 30562 8256 30618 8265
rect 30562 8191 30618 8200
rect 31666 8256 31722 8265
rect 31666 8191 31722 8200
rect 32954 8256 33010 8265
rect 32954 8191 33010 8200
rect 34242 8256 34298 8265
rect 34242 8191 34298 8200
rect 35438 8256 35494 8265
rect 35438 8191 35494 8200
rect 36358 8256 36414 8265
rect 36358 8191 36414 8200
rect 37462 8256 37518 8265
rect 37462 8191 37518 8200
rect 38750 8256 38806 8265
rect 38750 8191 38806 8200
rect 41326 8256 41382 8265
rect 41326 8191 41382 8200
rect 42154 8256 42210 8265
rect 42154 8191 42210 8200
rect 43442 8256 43498 8265
rect 43442 8191 43498 8200
rect 90638 8256 90694 8265
rect 90638 8191 90694 8200
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 23492 2650 23520 8191
rect 24780 2650 24808 8191
rect 25884 2650 25912 8191
rect 27172 2650 27200 8191
rect 28460 2650 28488 8191
rect 29288 2650 29316 8191
rect 30576 2650 30604 8191
rect 31680 2650 31708 8191
rect 32968 2650 32996 8191
rect 34256 2650 34284 8191
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35452 2650 35480 8191
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 36372 2650 36400 8191
rect 37476 2650 37504 8191
rect 38764 2650 38792 8191
rect 39946 4584 40002 4593
rect 39946 4519 40002 4528
rect 39960 2650 39988 4519
rect 41340 2650 41368 8191
rect 42168 2650 42196 8191
rect 43456 2650 43484 8191
rect 66314 7644 66622 7653
rect 66314 7642 66320 7644
rect 66376 7642 66400 7644
rect 66456 7642 66480 7644
rect 66536 7642 66560 7644
rect 66616 7642 66622 7644
rect 66376 7590 66378 7642
rect 66558 7590 66560 7642
rect 66314 7588 66320 7590
rect 66376 7588 66400 7590
rect 66456 7588 66480 7590
rect 66536 7588 66560 7590
rect 66616 7588 66622 7590
rect 66314 7579 66622 7588
rect 90652 7546 90680 8191
rect 90744 7546 90772 9687
rect 105922 9276 106230 9285
rect 105922 9274 105928 9276
rect 105984 9274 106008 9276
rect 106064 9274 106088 9276
rect 106144 9274 106168 9276
rect 106224 9274 106230 9276
rect 105984 9222 105986 9274
rect 106166 9222 106168 9274
rect 105922 9220 105928 9222
rect 105984 9220 106008 9222
rect 106064 9220 106088 9222
rect 106144 9220 106168 9222
rect 106224 9220 106230 9222
rect 105922 9211 106230 9220
rect 106658 8732 106966 8741
rect 106658 8730 106664 8732
rect 106720 8730 106744 8732
rect 106800 8730 106824 8732
rect 106880 8730 106904 8732
rect 106960 8730 106966 8732
rect 106720 8678 106722 8730
rect 106902 8678 106904 8730
rect 106658 8676 106664 8678
rect 106720 8676 106744 8678
rect 106800 8676 106824 8678
rect 106880 8676 106904 8678
rect 106960 8676 106966 8678
rect 106658 8667 106966 8676
rect 91006 8256 91062 8265
rect 91006 8191 91062 8200
rect 91020 7546 91048 8191
rect 105922 8188 106230 8197
rect 105922 8186 105928 8188
rect 105984 8186 106008 8188
rect 106064 8186 106088 8188
rect 106144 8186 106168 8188
rect 106224 8186 106230 8188
rect 105984 8134 105986 8186
rect 106166 8134 106168 8186
rect 105922 8132 105928 8134
rect 105984 8132 106008 8134
rect 106064 8132 106088 8134
rect 106144 8132 106168 8134
rect 106224 8132 106230 8134
rect 105922 8123 106230 8132
rect 97034 7644 97342 7653
rect 97034 7642 97040 7644
rect 97096 7642 97120 7644
rect 97176 7642 97200 7644
rect 97256 7642 97280 7644
rect 97336 7642 97342 7644
rect 97096 7590 97098 7642
rect 97278 7590 97280 7642
rect 97034 7588 97040 7590
rect 97096 7588 97120 7590
rect 97176 7588 97200 7590
rect 97256 7588 97280 7590
rect 97336 7588 97342 7590
rect 97034 7579 97342 7588
rect 106658 7644 106966 7653
rect 106658 7642 106664 7644
rect 106720 7642 106744 7644
rect 106800 7642 106824 7644
rect 106880 7642 106904 7644
rect 106960 7642 106966 7644
rect 106720 7590 106722 7642
rect 106902 7590 106904 7642
rect 106658 7588 106664 7590
rect 106720 7588 106744 7590
rect 106800 7588 106824 7590
rect 106880 7588 106904 7590
rect 106960 7588 106966 7590
rect 106658 7579 106966 7588
rect 90640 7540 90692 7546
rect 90640 7482 90692 7488
rect 90732 7540 90784 7546
rect 90732 7482 90784 7488
rect 91008 7540 91060 7546
rect 91008 7482 91060 7488
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 96374 7100 96682 7109
rect 96374 7098 96380 7100
rect 96436 7098 96460 7100
rect 96516 7098 96540 7100
rect 96596 7098 96620 7100
rect 96676 7098 96682 7100
rect 96436 7046 96438 7098
rect 96618 7046 96620 7098
rect 96374 7044 96380 7046
rect 96436 7044 96460 7046
rect 96516 7044 96540 7046
rect 96596 7044 96620 7046
rect 96676 7044 96682 7046
rect 96374 7035 96682 7044
rect 105922 7100 106230 7109
rect 105922 7098 105928 7100
rect 105984 7098 106008 7100
rect 106064 7098 106088 7100
rect 106144 7098 106168 7100
rect 106224 7098 106230 7100
rect 105984 7046 105986 7098
rect 106166 7046 106168 7098
rect 105922 7044 105928 7046
rect 105984 7044 106008 7046
rect 106064 7044 106088 7046
rect 106144 7044 106168 7046
rect 106224 7044 106230 7046
rect 105922 7035 106230 7044
rect 66314 6556 66622 6565
rect 66314 6554 66320 6556
rect 66376 6554 66400 6556
rect 66456 6554 66480 6556
rect 66536 6554 66560 6556
rect 66616 6554 66622 6556
rect 66376 6502 66378 6554
rect 66558 6502 66560 6554
rect 66314 6500 66320 6502
rect 66376 6500 66400 6502
rect 66456 6500 66480 6502
rect 66536 6500 66560 6502
rect 66616 6500 66622 6502
rect 66314 6491 66622 6500
rect 97034 6556 97342 6565
rect 97034 6554 97040 6556
rect 97096 6554 97120 6556
rect 97176 6554 97200 6556
rect 97256 6554 97280 6556
rect 97336 6554 97342 6556
rect 97096 6502 97098 6554
rect 97278 6502 97280 6554
rect 97034 6500 97040 6502
rect 97096 6500 97120 6502
rect 97176 6500 97200 6502
rect 97256 6500 97280 6502
rect 97336 6500 97342 6502
rect 97034 6491 97342 6500
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 96374 6012 96682 6021
rect 96374 6010 96380 6012
rect 96436 6010 96460 6012
rect 96516 6010 96540 6012
rect 96596 6010 96620 6012
rect 96676 6010 96682 6012
rect 96436 5958 96438 6010
rect 96618 5958 96620 6010
rect 96374 5956 96380 5958
rect 96436 5956 96460 5958
rect 96516 5956 96540 5958
rect 96596 5956 96620 5958
rect 96676 5956 96682 5958
rect 96374 5947 96682 5956
rect 66314 5468 66622 5477
rect 66314 5466 66320 5468
rect 66376 5466 66400 5468
rect 66456 5466 66480 5468
rect 66536 5466 66560 5468
rect 66616 5466 66622 5468
rect 66376 5414 66378 5466
rect 66558 5414 66560 5466
rect 66314 5412 66320 5414
rect 66376 5412 66400 5414
rect 66456 5412 66480 5414
rect 66536 5412 66560 5414
rect 66616 5412 66622 5414
rect 66314 5403 66622 5412
rect 97034 5468 97342 5477
rect 97034 5466 97040 5468
rect 97096 5466 97120 5468
rect 97176 5466 97200 5468
rect 97256 5466 97280 5468
rect 97336 5466 97342 5468
rect 97096 5414 97098 5466
rect 97278 5414 97280 5466
rect 97034 5412 97040 5414
rect 97096 5412 97120 5414
rect 97176 5412 97200 5414
rect 97256 5412 97280 5414
rect 97336 5412 97342 5414
rect 97034 5403 97342 5412
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 96374 4924 96682 4933
rect 96374 4922 96380 4924
rect 96436 4922 96460 4924
rect 96516 4922 96540 4924
rect 96596 4922 96620 4924
rect 96676 4922 96682 4924
rect 96436 4870 96438 4922
rect 96618 4870 96620 4922
rect 96374 4868 96380 4870
rect 96436 4868 96460 4870
rect 96516 4868 96540 4870
rect 96596 4868 96620 4870
rect 96676 4868 96682 4870
rect 96374 4859 96682 4868
rect 66314 4380 66622 4389
rect 66314 4378 66320 4380
rect 66376 4378 66400 4380
rect 66456 4378 66480 4380
rect 66536 4378 66560 4380
rect 66616 4378 66622 4380
rect 66376 4326 66378 4378
rect 66558 4326 66560 4378
rect 66314 4324 66320 4326
rect 66376 4324 66400 4326
rect 66456 4324 66480 4326
rect 66536 4324 66560 4326
rect 66616 4324 66622 4326
rect 66314 4315 66622 4324
rect 97034 4380 97342 4389
rect 97034 4378 97040 4380
rect 97096 4378 97120 4380
rect 97176 4378 97200 4380
rect 97256 4378 97280 4380
rect 97336 4378 97342 4380
rect 97096 4326 97098 4378
rect 97278 4326 97280 4378
rect 97034 4324 97040 4326
rect 97096 4324 97120 4326
rect 97176 4324 97200 4326
rect 97256 4324 97280 4326
rect 97336 4324 97342 4326
rect 97034 4315 97342 4324
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 96374 3836 96682 3845
rect 96374 3834 96380 3836
rect 96436 3834 96460 3836
rect 96516 3834 96540 3836
rect 96596 3834 96620 3836
rect 96676 3834 96682 3836
rect 96436 3782 96438 3834
rect 96618 3782 96620 3834
rect 96374 3780 96380 3782
rect 96436 3780 96460 3782
rect 96516 3780 96540 3782
rect 96596 3780 96620 3782
rect 96676 3780 96682 3782
rect 96374 3771 96682 3780
rect 66314 3292 66622 3301
rect 66314 3290 66320 3292
rect 66376 3290 66400 3292
rect 66456 3290 66480 3292
rect 66536 3290 66560 3292
rect 66616 3290 66622 3292
rect 66376 3238 66378 3290
rect 66558 3238 66560 3290
rect 66314 3236 66320 3238
rect 66376 3236 66400 3238
rect 66456 3236 66480 3238
rect 66536 3236 66560 3238
rect 66616 3236 66622 3238
rect 66314 3227 66622 3236
rect 97034 3292 97342 3301
rect 97034 3290 97040 3292
rect 97096 3290 97120 3292
rect 97176 3290 97200 3292
rect 97256 3290 97280 3292
rect 97336 3290 97342 3292
rect 97096 3238 97098 3290
rect 97278 3238 97280 3290
rect 97034 3236 97040 3238
rect 97096 3236 97120 3238
rect 97176 3236 97200 3238
rect 97256 3236 97280 3238
rect 97336 3236 97342 3238
rect 97034 3227 97342 3236
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 96374 2748 96682 2757
rect 96374 2746 96380 2748
rect 96436 2746 96460 2748
rect 96516 2746 96540 2748
rect 96596 2746 96620 2748
rect 96676 2746 96682 2748
rect 96436 2694 96438 2746
rect 96618 2694 96620 2746
rect 96374 2692 96380 2694
rect 96436 2692 96460 2694
rect 96516 2692 96540 2694
rect 96596 2692 96620 2694
rect 96676 2692 96682 2694
rect 96374 2683 96682 2692
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 25872 2644 25924 2650
rect 25872 2586 25924 2592
rect 27160 2644 27212 2650
rect 27160 2586 27212 2592
rect 28448 2644 28500 2650
rect 28448 2586 28500 2592
rect 29276 2644 29328 2650
rect 29276 2586 29328 2592
rect 30564 2644 30616 2650
rect 30564 2586 30616 2592
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 32956 2644 33008 2650
rect 32956 2586 33008 2592
rect 34244 2644 34296 2650
rect 34244 2586 34296 2592
rect 35440 2644 35492 2650
rect 35440 2586 35492 2592
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 38752 2644 38804 2650
rect 38752 2586 38804 2592
rect 39948 2644 40000 2650
rect 39948 2586 40000 2592
rect 41328 2644 41380 2650
rect 41328 2586 41380 2592
rect 42156 2644 42208 2650
rect 42156 2586 42208 2592
rect 43444 2644 43496 2650
rect 43444 2586 43496 2592
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 28356 2304 28408 2310
rect 28356 2246 28408 2252
rect 29000 2304 29052 2310
rect 29000 2246 29052 2252
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 39948 2304 40000 2310
rect 39948 2246 40000 2252
rect 41236 2304 41288 2310
rect 41236 2246 41288 2252
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 43168 2304 43220 2310
rect 43168 2246 43220 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 23216 800 23244 2246
rect 24504 800 24532 2246
rect 25792 800 25820 2246
rect 27080 800 27108 2246
rect 28368 800 28396 2246
rect 29012 800 29040 2246
rect 30300 800 30328 2246
rect 31588 800 31616 2246
rect 32876 800 32904 2246
rect 34164 800 34192 2246
rect 35452 800 35480 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 36096 800 36124 2246
rect 37384 800 37412 2246
rect 38672 800 38700 2246
rect 39960 800 39988 2246
rect 41248 800 41276 2246
rect 41892 800 41920 2246
rect 43180 800 43208 2246
rect 66314 2204 66622 2213
rect 66314 2202 66320 2204
rect 66376 2202 66400 2204
rect 66456 2202 66480 2204
rect 66536 2202 66560 2204
rect 66616 2202 66622 2204
rect 66376 2150 66378 2202
rect 66558 2150 66560 2202
rect 66314 2148 66320 2150
rect 66376 2148 66400 2150
rect 66456 2148 66480 2150
rect 66536 2148 66560 2150
rect 66616 2148 66622 2150
rect 66314 2139 66622 2148
rect 97034 2204 97342 2213
rect 97034 2202 97040 2204
rect 97096 2202 97120 2204
rect 97176 2202 97200 2204
rect 97256 2202 97280 2204
rect 97336 2202 97342 2204
rect 97096 2150 97098 2202
rect 97278 2150 97280 2202
rect 97034 2148 97040 2150
rect 97096 2148 97120 2150
rect 97176 2148 97200 2150
rect 97256 2148 97280 2150
rect 97336 2148 97342 2150
rect 97034 2139 97342 2148
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 30286 0 30342 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 43166 0 43222 800
<< via2 >>
rect 4880 127322 4936 127324
rect 4960 127322 5016 127324
rect 5040 127322 5096 127324
rect 5120 127322 5176 127324
rect 4880 127270 4926 127322
rect 4926 127270 4936 127322
rect 4960 127270 4990 127322
rect 4990 127270 5002 127322
rect 5002 127270 5016 127322
rect 5040 127270 5054 127322
rect 5054 127270 5066 127322
rect 5066 127270 5096 127322
rect 5120 127270 5130 127322
rect 5130 127270 5176 127322
rect 4880 127268 4936 127270
rect 4960 127268 5016 127270
rect 5040 127268 5096 127270
rect 5120 127268 5176 127270
rect 35600 127322 35656 127324
rect 35680 127322 35736 127324
rect 35760 127322 35816 127324
rect 35840 127322 35896 127324
rect 35600 127270 35646 127322
rect 35646 127270 35656 127322
rect 35680 127270 35710 127322
rect 35710 127270 35722 127322
rect 35722 127270 35736 127322
rect 35760 127270 35774 127322
rect 35774 127270 35786 127322
rect 35786 127270 35816 127322
rect 35840 127270 35850 127322
rect 35850 127270 35896 127322
rect 35600 127268 35656 127270
rect 35680 127268 35736 127270
rect 35760 127268 35816 127270
rect 35840 127268 35896 127270
rect 66320 127322 66376 127324
rect 66400 127322 66456 127324
rect 66480 127322 66536 127324
rect 66560 127322 66616 127324
rect 66320 127270 66366 127322
rect 66366 127270 66376 127322
rect 66400 127270 66430 127322
rect 66430 127270 66442 127322
rect 66442 127270 66456 127322
rect 66480 127270 66494 127322
rect 66494 127270 66506 127322
rect 66506 127270 66536 127322
rect 66560 127270 66570 127322
rect 66570 127270 66616 127322
rect 66320 127268 66376 127270
rect 66400 127268 66456 127270
rect 66480 127268 66536 127270
rect 66560 127268 66616 127270
rect 97040 127322 97096 127324
rect 97120 127322 97176 127324
rect 97200 127322 97256 127324
rect 97280 127322 97336 127324
rect 97040 127270 97086 127322
rect 97086 127270 97096 127322
rect 97120 127270 97150 127322
rect 97150 127270 97162 127322
rect 97162 127270 97176 127322
rect 97200 127270 97214 127322
rect 97214 127270 97226 127322
rect 97226 127270 97256 127322
rect 97280 127270 97290 127322
rect 97290 127270 97336 127322
rect 97040 127268 97096 127270
rect 97120 127268 97176 127270
rect 97200 127268 97256 127270
rect 97280 127268 97336 127270
rect 4220 126778 4276 126780
rect 4300 126778 4356 126780
rect 4380 126778 4436 126780
rect 4460 126778 4516 126780
rect 4220 126726 4266 126778
rect 4266 126726 4276 126778
rect 4300 126726 4330 126778
rect 4330 126726 4342 126778
rect 4342 126726 4356 126778
rect 4380 126726 4394 126778
rect 4394 126726 4406 126778
rect 4406 126726 4436 126778
rect 4460 126726 4470 126778
rect 4470 126726 4516 126778
rect 4220 126724 4276 126726
rect 4300 126724 4356 126726
rect 4380 126724 4436 126726
rect 4460 126724 4516 126726
rect 34940 126778 34996 126780
rect 35020 126778 35076 126780
rect 35100 126778 35156 126780
rect 35180 126778 35236 126780
rect 34940 126726 34986 126778
rect 34986 126726 34996 126778
rect 35020 126726 35050 126778
rect 35050 126726 35062 126778
rect 35062 126726 35076 126778
rect 35100 126726 35114 126778
rect 35114 126726 35126 126778
rect 35126 126726 35156 126778
rect 35180 126726 35190 126778
rect 35190 126726 35236 126778
rect 34940 126724 34996 126726
rect 35020 126724 35076 126726
rect 35100 126724 35156 126726
rect 35180 126724 35236 126726
rect 65660 126778 65716 126780
rect 65740 126778 65796 126780
rect 65820 126778 65876 126780
rect 65900 126778 65956 126780
rect 65660 126726 65706 126778
rect 65706 126726 65716 126778
rect 65740 126726 65770 126778
rect 65770 126726 65782 126778
rect 65782 126726 65796 126778
rect 65820 126726 65834 126778
rect 65834 126726 65846 126778
rect 65846 126726 65876 126778
rect 65900 126726 65910 126778
rect 65910 126726 65956 126778
rect 65660 126724 65716 126726
rect 65740 126724 65796 126726
rect 65820 126724 65876 126726
rect 65900 126724 65956 126726
rect 96380 126778 96436 126780
rect 96460 126778 96516 126780
rect 96540 126778 96596 126780
rect 96620 126778 96676 126780
rect 96380 126726 96426 126778
rect 96426 126726 96436 126778
rect 96460 126726 96490 126778
rect 96490 126726 96502 126778
rect 96502 126726 96516 126778
rect 96540 126726 96554 126778
rect 96554 126726 96566 126778
rect 96566 126726 96596 126778
rect 96620 126726 96630 126778
rect 96630 126726 96676 126778
rect 96380 126724 96436 126726
rect 96460 126724 96516 126726
rect 96540 126724 96596 126726
rect 96620 126724 96676 126726
rect 4880 126234 4936 126236
rect 4960 126234 5016 126236
rect 5040 126234 5096 126236
rect 5120 126234 5176 126236
rect 4880 126182 4926 126234
rect 4926 126182 4936 126234
rect 4960 126182 4990 126234
rect 4990 126182 5002 126234
rect 5002 126182 5016 126234
rect 5040 126182 5054 126234
rect 5054 126182 5066 126234
rect 5066 126182 5096 126234
rect 5120 126182 5130 126234
rect 5130 126182 5176 126234
rect 4880 126180 4936 126182
rect 4960 126180 5016 126182
rect 5040 126180 5096 126182
rect 5120 126180 5176 126182
rect 35600 126234 35656 126236
rect 35680 126234 35736 126236
rect 35760 126234 35816 126236
rect 35840 126234 35896 126236
rect 35600 126182 35646 126234
rect 35646 126182 35656 126234
rect 35680 126182 35710 126234
rect 35710 126182 35722 126234
rect 35722 126182 35736 126234
rect 35760 126182 35774 126234
rect 35774 126182 35786 126234
rect 35786 126182 35816 126234
rect 35840 126182 35850 126234
rect 35850 126182 35896 126234
rect 35600 126180 35656 126182
rect 35680 126180 35736 126182
rect 35760 126180 35816 126182
rect 35840 126180 35896 126182
rect 4220 125690 4276 125692
rect 4300 125690 4356 125692
rect 4380 125690 4436 125692
rect 4460 125690 4516 125692
rect 4220 125638 4266 125690
rect 4266 125638 4276 125690
rect 4300 125638 4330 125690
rect 4330 125638 4342 125690
rect 4342 125638 4356 125690
rect 4380 125638 4394 125690
rect 4394 125638 4406 125690
rect 4406 125638 4436 125690
rect 4460 125638 4470 125690
rect 4470 125638 4516 125690
rect 4220 125636 4276 125638
rect 4300 125636 4356 125638
rect 4380 125636 4436 125638
rect 4460 125636 4516 125638
rect 4880 125146 4936 125148
rect 4960 125146 5016 125148
rect 5040 125146 5096 125148
rect 5120 125146 5176 125148
rect 4880 125094 4926 125146
rect 4926 125094 4936 125146
rect 4960 125094 4990 125146
rect 4990 125094 5002 125146
rect 5002 125094 5016 125146
rect 5040 125094 5054 125146
rect 5054 125094 5066 125146
rect 5066 125094 5096 125146
rect 5120 125094 5130 125146
rect 5130 125094 5176 125146
rect 4880 125092 4936 125094
rect 4960 125092 5016 125094
rect 5040 125092 5096 125094
rect 5120 125092 5176 125094
rect 4220 124602 4276 124604
rect 4300 124602 4356 124604
rect 4380 124602 4436 124604
rect 4460 124602 4516 124604
rect 4220 124550 4266 124602
rect 4266 124550 4276 124602
rect 4300 124550 4330 124602
rect 4330 124550 4342 124602
rect 4342 124550 4356 124602
rect 4380 124550 4394 124602
rect 4394 124550 4406 124602
rect 4406 124550 4436 124602
rect 4460 124550 4470 124602
rect 4470 124550 4516 124602
rect 4220 124548 4276 124550
rect 4300 124548 4356 124550
rect 4380 124548 4436 124550
rect 4460 124548 4516 124550
rect 4880 124058 4936 124060
rect 4960 124058 5016 124060
rect 5040 124058 5096 124060
rect 5120 124058 5176 124060
rect 4880 124006 4926 124058
rect 4926 124006 4936 124058
rect 4960 124006 4990 124058
rect 4990 124006 5002 124058
rect 5002 124006 5016 124058
rect 5040 124006 5054 124058
rect 5054 124006 5066 124058
rect 5066 124006 5096 124058
rect 5120 124006 5130 124058
rect 5130 124006 5176 124058
rect 4880 124004 4936 124006
rect 4960 124004 5016 124006
rect 5040 124004 5096 124006
rect 5120 124004 5176 124006
rect 4220 123514 4276 123516
rect 4300 123514 4356 123516
rect 4380 123514 4436 123516
rect 4460 123514 4516 123516
rect 4220 123462 4266 123514
rect 4266 123462 4276 123514
rect 4300 123462 4330 123514
rect 4330 123462 4342 123514
rect 4342 123462 4356 123514
rect 4380 123462 4394 123514
rect 4394 123462 4406 123514
rect 4406 123462 4436 123514
rect 4460 123462 4470 123514
rect 4470 123462 4516 123514
rect 4220 123460 4276 123462
rect 4300 123460 4356 123462
rect 4380 123460 4436 123462
rect 4460 123460 4516 123462
rect 4880 122970 4936 122972
rect 4960 122970 5016 122972
rect 5040 122970 5096 122972
rect 5120 122970 5176 122972
rect 4880 122918 4926 122970
rect 4926 122918 4936 122970
rect 4960 122918 4990 122970
rect 4990 122918 5002 122970
rect 5002 122918 5016 122970
rect 5040 122918 5054 122970
rect 5054 122918 5066 122970
rect 5066 122918 5096 122970
rect 5120 122918 5130 122970
rect 5130 122918 5176 122970
rect 4880 122916 4936 122918
rect 4960 122916 5016 122918
rect 5040 122916 5096 122918
rect 5120 122916 5176 122918
rect 4220 122426 4276 122428
rect 4300 122426 4356 122428
rect 4380 122426 4436 122428
rect 4460 122426 4516 122428
rect 4220 122374 4266 122426
rect 4266 122374 4276 122426
rect 4300 122374 4330 122426
rect 4330 122374 4342 122426
rect 4342 122374 4356 122426
rect 4380 122374 4394 122426
rect 4394 122374 4406 122426
rect 4406 122374 4436 122426
rect 4460 122374 4470 122426
rect 4470 122374 4516 122426
rect 4220 122372 4276 122374
rect 4300 122372 4356 122374
rect 4380 122372 4436 122374
rect 4460 122372 4516 122374
rect 4880 121882 4936 121884
rect 4960 121882 5016 121884
rect 5040 121882 5096 121884
rect 5120 121882 5176 121884
rect 4880 121830 4926 121882
rect 4926 121830 4936 121882
rect 4960 121830 4990 121882
rect 4990 121830 5002 121882
rect 5002 121830 5016 121882
rect 5040 121830 5054 121882
rect 5054 121830 5066 121882
rect 5066 121830 5096 121882
rect 5120 121830 5130 121882
rect 5130 121830 5176 121882
rect 4880 121828 4936 121830
rect 4960 121828 5016 121830
rect 5040 121828 5096 121830
rect 5120 121828 5176 121830
rect 4220 121338 4276 121340
rect 4300 121338 4356 121340
rect 4380 121338 4436 121340
rect 4460 121338 4516 121340
rect 4220 121286 4266 121338
rect 4266 121286 4276 121338
rect 4300 121286 4330 121338
rect 4330 121286 4342 121338
rect 4342 121286 4356 121338
rect 4380 121286 4394 121338
rect 4394 121286 4406 121338
rect 4406 121286 4436 121338
rect 4460 121286 4470 121338
rect 4470 121286 4516 121338
rect 4220 121284 4276 121286
rect 4300 121284 4356 121286
rect 4380 121284 4436 121286
rect 4460 121284 4516 121286
rect 4880 120794 4936 120796
rect 4960 120794 5016 120796
rect 5040 120794 5096 120796
rect 5120 120794 5176 120796
rect 4880 120742 4926 120794
rect 4926 120742 4936 120794
rect 4960 120742 4990 120794
rect 4990 120742 5002 120794
rect 5002 120742 5016 120794
rect 5040 120742 5054 120794
rect 5054 120742 5066 120794
rect 5066 120742 5096 120794
rect 5120 120742 5130 120794
rect 5130 120742 5176 120794
rect 4880 120740 4936 120742
rect 4960 120740 5016 120742
rect 5040 120740 5096 120742
rect 5120 120740 5176 120742
rect 4220 120250 4276 120252
rect 4300 120250 4356 120252
rect 4380 120250 4436 120252
rect 4460 120250 4516 120252
rect 4220 120198 4266 120250
rect 4266 120198 4276 120250
rect 4300 120198 4330 120250
rect 4330 120198 4342 120250
rect 4342 120198 4356 120250
rect 4380 120198 4394 120250
rect 4394 120198 4406 120250
rect 4406 120198 4436 120250
rect 4460 120198 4470 120250
rect 4470 120198 4516 120250
rect 4220 120196 4276 120198
rect 4300 120196 4356 120198
rect 4380 120196 4436 120198
rect 4460 120196 4516 120198
rect 4880 119706 4936 119708
rect 4960 119706 5016 119708
rect 5040 119706 5096 119708
rect 5120 119706 5176 119708
rect 4880 119654 4926 119706
rect 4926 119654 4936 119706
rect 4960 119654 4990 119706
rect 4990 119654 5002 119706
rect 5002 119654 5016 119706
rect 5040 119654 5054 119706
rect 5054 119654 5066 119706
rect 5066 119654 5096 119706
rect 5120 119654 5130 119706
rect 5130 119654 5176 119706
rect 4880 119652 4936 119654
rect 4960 119652 5016 119654
rect 5040 119652 5096 119654
rect 5120 119652 5176 119654
rect 4220 119162 4276 119164
rect 4300 119162 4356 119164
rect 4380 119162 4436 119164
rect 4460 119162 4516 119164
rect 4220 119110 4266 119162
rect 4266 119110 4276 119162
rect 4300 119110 4330 119162
rect 4330 119110 4342 119162
rect 4342 119110 4356 119162
rect 4380 119110 4394 119162
rect 4394 119110 4406 119162
rect 4406 119110 4436 119162
rect 4460 119110 4470 119162
rect 4470 119110 4516 119162
rect 4220 119108 4276 119110
rect 4300 119108 4356 119110
rect 4380 119108 4436 119110
rect 4460 119108 4516 119110
rect 4880 118618 4936 118620
rect 4960 118618 5016 118620
rect 5040 118618 5096 118620
rect 5120 118618 5176 118620
rect 4880 118566 4926 118618
rect 4926 118566 4936 118618
rect 4960 118566 4990 118618
rect 4990 118566 5002 118618
rect 5002 118566 5016 118618
rect 5040 118566 5054 118618
rect 5054 118566 5066 118618
rect 5066 118566 5096 118618
rect 5120 118566 5130 118618
rect 5130 118566 5176 118618
rect 4880 118564 4936 118566
rect 4960 118564 5016 118566
rect 5040 118564 5096 118566
rect 5120 118564 5176 118566
rect 4220 118074 4276 118076
rect 4300 118074 4356 118076
rect 4380 118074 4436 118076
rect 4460 118074 4516 118076
rect 4220 118022 4266 118074
rect 4266 118022 4276 118074
rect 4300 118022 4330 118074
rect 4330 118022 4342 118074
rect 4342 118022 4356 118074
rect 4380 118022 4394 118074
rect 4394 118022 4406 118074
rect 4406 118022 4436 118074
rect 4460 118022 4470 118074
rect 4470 118022 4516 118074
rect 4220 118020 4276 118022
rect 4300 118020 4356 118022
rect 4380 118020 4436 118022
rect 4460 118020 4516 118022
rect 4880 117530 4936 117532
rect 4960 117530 5016 117532
rect 5040 117530 5096 117532
rect 5120 117530 5176 117532
rect 4880 117478 4926 117530
rect 4926 117478 4936 117530
rect 4960 117478 4990 117530
rect 4990 117478 5002 117530
rect 5002 117478 5016 117530
rect 5040 117478 5054 117530
rect 5054 117478 5066 117530
rect 5066 117478 5096 117530
rect 5120 117478 5130 117530
rect 5130 117478 5176 117530
rect 4880 117476 4936 117478
rect 4960 117476 5016 117478
rect 5040 117476 5096 117478
rect 5120 117476 5176 117478
rect 4220 116986 4276 116988
rect 4300 116986 4356 116988
rect 4380 116986 4436 116988
rect 4460 116986 4516 116988
rect 4220 116934 4266 116986
rect 4266 116934 4276 116986
rect 4300 116934 4330 116986
rect 4330 116934 4342 116986
rect 4342 116934 4356 116986
rect 4380 116934 4394 116986
rect 4394 116934 4406 116986
rect 4406 116934 4436 116986
rect 4460 116934 4470 116986
rect 4470 116934 4516 116986
rect 4220 116932 4276 116934
rect 4300 116932 4356 116934
rect 4380 116932 4436 116934
rect 4460 116932 4516 116934
rect 4880 116442 4936 116444
rect 4960 116442 5016 116444
rect 5040 116442 5096 116444
rect 5120 116442 5176 116444
rect 4880 116390 4926 116442
rect 4926 116390 4936 116442
rect 4960 116390 4990 116442
rect 4990 116390 5002 116442
rect 5002 116390 5016 116442
rect 5040 116390 5054 116442
rect 5054 116390 5066 116442
rect 5066 116390 5096 116442
rect 5120 116390 5130 116442
rect 5130 116390 5176 116442
rect 4880 116388 4936 116390
rect 4960 116388 5016 116390
rect 5040 116388 5096 116390
rect 5120 116388 5176 116390
rect 4220 115898 4276 115900
rect 4300 115898 4356 115900
rect 4380 115898 4436 115900
rect 4460 115898 4516 115900
rect 4220 115846 4266 115898
rect 4266 115846 4276 115898
rect 4300 115846 4330 115898
rect 4330 115846 4342 115898
rect 4342 115846 4356 115898
rect 4380 115846 4394 115898
rect 4394 115846 4406 115898
rect 4406 115846 4436 115898
rect 4460 115846 4470 115898
rect 4470 115846 4516 115898
rect 4220 115844 4276 115846
rect 4300 115844 4356 115846
rect 4380 115844 4436 115846
rect 4460 115844 4516 115846
rect 4880 115354 4936 115356
rect 4960 115354 5016 115356
rect 5040 115354 5096 115356
rect 5120 115354 5176 115356
rect 4880 115302 4926 115354
rect 4926 115302 4936 115354
rect 4960 115302 4990 115354
rect 4990 115302 5002 115354
rect 5002 115302 5016 115354
rect 5040 115302 5054 115354
rect 5054 115302 5066 115354
rect 5066 115302 5096 115354
rect 5120 115302 5130 115354
rect 5130 115302 5176 115354
rect 4880 115300 4936 115302
rect 4960 115300 5016 115302
rect 5040 115300 5096 115302
rect 5120 115300 5176 115302
rect 4220 114810 4276 114812
rect 4300 114810 4356 114812
rect 4380 114810 4436 114812
rect 4460 114810 4516 114812
rect 4220 114758 4266 114810
rect 4266 114758 4276 114810
rect 4300 114758 4330 114810
rect 4330 114758 4342 114810
rect 4342 114758 4356 114810
rect 4380 114758 4394 114810
rect 4394 114758 4406 114810
rect 4406 114758 4436 114810
rect 4460 114758 4470 114810
rect 4470 114758 4516 114810
rect 4220 114756 4276 114758
rect 4300 114756 4356 114758
rect 4380 114756 4436 114758
rect 4460 114756 4516 114758
rect 4880 114266 4936 114268
rect 4960 114266 5016 114268
rect 5040 114266 5096 114268
rect 5120 114266 5176 114268
rect 4880 114214 4926 114266
rect 4926 114214 4936 114266
rect 4960 114214 4990 114266
rect 4990 114214 5002 114266
rect 5002 114214 5016 114266
rect 5040 114214 5054 114266
rect 5054 114214 5066 114266
rect 5066 114214 5096 114266
rect 5120 114214 5130 114266
rect 5130 114214 5176 114266
rect 4880 114212 4936 114214
rect 4960 114212 5016 114214
rect 5040 114212 5096 114214
rect 5120 114212 5176 114214
rect 4220 113722 4276 113724
rect 4300 113722 4356 113724
rect 4380 113722 4436 113724
rect 4460 113722 4516 113724
rect 4220 113670 4266 113722
rect 4266 113670 4276 113722
rect 4300 113670 4330 113722
rect 4330 113670 4342 113722
rect 4342 113670 4356 113722
rect 4380 113670 4394 113722
rect 4394 113670 4406 113722
rect 4406 113670 4436 113722
rect 4460 113670 4470 113722
rect 4470 113670 4516 113722
rect 4220 113668 4276 113670
rect 4300 113668 4356 113670
rect 4380 113668 4436 113670
rect 4460 113668 4516 113670
rect 4880 113178 4936 113180
rect 4960 113178 5016 113180
rect 5040 113178 5096 113180
rect 5120 113178 5176 113180
rect 4880 113126 4926 113178
rect 4926 113126 4936 113178
rect 4960 113126 4990 113178
rect 4990 113126 5002 113178
rect 5002 113126 5016 113178
rect 5040 113126 5054 113178
rect 5054 113126 5066 113178
rect 5066 113126 5096 113178
rect 5120 113126 5130 113178
rect 5130 113126 5176 113178
rect 4880 113124 4936 113126
rect 4960 113124 5016 113126
rect 5040 113124 5096 113126
rect 5120 113124 5176 113126
rect 4220 112634 4276 112636
rect 4300 112634 4356 112636
rect 4380 112634 4436 112636
rect 4460 112634 4516 112636
rect 4220 112582 4266 112634
rect 4266 112582 4276 112634
rect 4300 112582 4330 112634
rect 4330 112582 4342 112634
rect 4342 112582 4356 112634
rect 4380 112582 4394 112634
rect 4394 112582 4406 112634
rect 4406 112582 4436 112634
rect 4460 112582 4470 112634
rect 4470 112582 4516 112634
rect 4220 112580 4276 112582
rect 4300 112580 4356 112582
rect 4380 112580 4436 112582
rect 4460 112580 4516 112582
rect 4880 112090 4936 112092
rect 4960 112090 5016 112092
rect 5040 112090 5096 112092
rect 5120 112090 5176 112092
rect 4880 112038 4926 112090
rect 4926 112038 4936 112090
rect 4960 112038 4990 112090
rect 4990 112038 5002 112090
rect 5002 112038 5016 112090
rect 5040 112038 5054 112090
rect 5054 112038 5066 112090
rect 5066 112038 5096 112090
rect 5120 112038 5130 112090
rect 5130 112038 5176 112090
rect 4880 112036 4936 112038
rect 4960 112036 5016 112038
rect 5040 112036 5096 112038
rect 5120 112036 5176 112038
rect 4220 111546 4276 111548
rect 4300 111546 4356 111548
rect 4380 111546 4436 111548
rect 4460 111546 4516 111548
rect 4220 111494 4266 111546
rect 4266 111494 4276 111546
rect 4300 111494 4330 111546
rect 4330 111494 4342 111546
rect 4342 111494 4356 111546
rect 4380 111494 4394 111546
rect 4394 111494 4406 111546
rect 4406 111494 4436 111546
rect 4460 111494 4470 111546
rect 4470 111494 4516 111546
rect 4220 111492 4276 111494
rect 4300 111492 4356 111494
rect 4380 111492 4436 111494
rect 4460 111492 4516 111494
rect 4880 111002 4936 111004
rect 4960 111002 5016 111004
rect 5040 111002 5096 111004
rect 5120 111002 5176 111004
rect 4880 110950 4926 111002
rect 4926 110950 4936 111002
rect 4960 110950 4990 111002
rect 4990 110950 5002 111002
rect 5002 110950 5016 111002
rect 5040 110950 5054 111002
rect 5054 110950 5066 111002
rect 5066 110950 5096 111002
rect 5120 110950 5130 111002
rect 5130 110950 5176 111002
rect 4880 110948 4936 110950
rect 4960 110948 5016 110950
rect 5040 110948 5096 110950
rect 5120 110948 5176 110950
rect 4220 110458 4276 110460
rect 4300 110458 4356 110460
rect 4380 110458 4436 110460
rect 4460 110458 4516 110460
rect 4220 110406 4266 110458
rect 4266 110406 4276 110458
rect 4300 110406 4330 110458
rect 4330 110406 4342 110458
rect 4342 110406 4356 110458
rect 4380 110406 4394 110458
rect 4394 110406 4406 110458
rect 4406 110406 4436 110458
rect 4460 110406 4470 110458
rect 4470 110406 4516 110458
rect 4220 110404 4276 110406
rect 4300 110404 4356 110406
rect 4380 110404 4436 110406
rect 4460 110404 4516 110406
rect 4880 109914 4936 109916
rect 4960 109914 5016 109916
rect 5040 109914 5096 109916
rect 5120 109914 5176 109916
rect 4880 109862 4926 109914
rect 4926 109862 4936 109914
rect 4960 109862 4990 109914
rect 4990 109862 5002 109914
rect 5002 109862 5016 109914
rect 5040 109862 5054 109914
rect 5054 109862 5066 109914
rect 5066 109862 5096 109914
rect 5120 109862 5130 109914
rect 5130 109862 5176 109914
rect 4880 109860 4936 109862
rect 4960 109860 5016 109862
rect 5040 109860 5096 109862
rect 5120 109860 5176 109862
rect 4220 109370 4276 109372
rect 4300 109370 4356 109372
rect 4380 109370 4436 109372
rect 4460 109370 4516 109372
rect 4220 109318 4266 109370
rect 4266 109318 4276 109370
rect 4300 109318 4330 109370
rect 4330 109318 4342 109370
rect 4342 109318 4356 109370
rect 4380 109318 4394 109370
rect 4394 109318 4406 109370
rect 4406 109318 4436 109370
rect 4460 109318 4470 109370
rect 4470 109318 4516 109370
rect 4220 109316 4276 109318
rect 4300 109316 4356 109318
rect 4380 109316 4436 109318
rect 4460 109316 4516 109318
rect 4880 108826 4936 108828
rect 4960 108826 5016 108828
rect 5040 108826 5096 108828
rect 5120 108826 5176 108828
rect 4880 108774 4926 108826
rect 4926 108774 4936 108826
rect 4960 108774 4990 108826
rect 4990 108774 5002 108826
rect 5002 108774 5016 108826
rect 5040 108774 5054 108826
rect 5054 108774 5066 108826
rect 5066 108774 5096 108826
rect 5120 108774 5130 108826
rect 5130 108774 5176 108826
rect 4880 108772 4936 108774
rect 4960 108772 5016 108774
rect 5040 108772 5096 108774
rect 5120 108772 5176 108774
rect 4220 108282 4276 108284
rect 4300 108282 4356 108284
rect 4380 108282 4436 108284
rect 4460 108282 4516 108284
rect 4220 108230 4266 108282
rect 4266 108230 4276 108282
rect 4300 108230 4330 108282
rect 4330 108230 4342 108282
rect 4342 108230 4356 108282
rect 4380 108230 4394 108282
rect 4394 108230 4406 108282
rect 4406 108230 4436 108282
rect 4460 108230 4470 108282
rect 4470 108230 4516 108282
rect 4220 108228 4276 108230
rect 4300 108228 4356 108230
rect 4380 108228 4436 108230
rect 4460 108228 4516 108230
rect 4880 107738 4936 107740
rect 4960 107738 5016 107740
rect 5040 107738 5096 107740
rect 5120 107738 5176 107740
rect 4880 107686 4926 107738
rect 4926 107686 4936 107738
rect 4960 107686 4990 107738
rect 4990 107686 5002 107738
rect 5002 107686 5016 107738
rect 5040 107686 5054 107738
rect 5054 107686 5066 107738
rect 5066 107686 5096 107738
rect 5120 107686 5130 107738
rect 5130 107686 5176 107738
rect 4880 107684 4936 107686
rect 4960 107684 5016 107686
rect 5040 107684 5096 107686
rect 5120 107684 5176 107686
rect 4220 107194 4276 107196
rect 4300 107194 4356 107196
rect 4380 107194 4436 107196
rect 4460 107194 4516 107196
rect 4220 107142 4266 107194
rect 4266 107142 4276 107194
rect 4300 107142 4330 107194
rect 4330 107142 4342 107194
rect 4342 107142 4356 107194
rect 4380 107142 4394 107194
rect 4394 107142 4406 107194
rect 4406 107142 4436 107194
rect 4460 107142 4470 107194
rect 4470 107142 4516 107194
rect 4220 107140 4276 107142
rect 4300 107140 4356 107142
rect 4380 107140 4436 107142
rect 4460 107140 4516 107142
rect 4880 106650 4936 106652
rect 4960 106650 5016 106652
rect 5040 106650 5096 106652
rect 5120 106650 5176 106652
rect 4880 106598 4926 106650
rect 4926 106598 4936 106650
rect 4960 106598 4990 106650
rect 4990 106598 5002 106650
rect 5002 106598 5016 106650
rect 5040 106598 5054 106650
rect 5054 106598 5066 106650
rect 5066 106598 5096 106650
rect 5120 106598 5130 106650
rect 5130 106598 5176 106650
rect 4880 106596 4936 106598
rect 4960 106596 5016 106598
rect 5040 106596 5096 106598
rect 5120 106596 5176 106598
rect 4220 106106 4276 106108
rect 4300 106106 4356 106108
rect 4380 106106 4436 106108
rect 4460 106106 4516 106108
rect 4220 106054 4266 106106
rect 4266 106054 4276 106106
rect 4300 106054 4330 106106
rect 4330 106054 4342 106106
rect 4342 106054 4356 106106
rect 4380 106054 4394 106106
rect 4394 106054 4406 106106
rect 4406 106054 4436 106106
rect 4460 106054 4470 106106
rect 4470 106054 4516 106106
rect 4220 106052 4276 106054
rect 4300 106052 4356 106054
rect 4380 106052 4436 106054
rect 4460 106052 4516 106054
rect 4880 105562 4936 105564
rect 4960 105562 5016 105564
rect 5040 105562 5096 105564
rect 5120 105562 5176 105564
rect 4880 105510 4926 105562
rect 4926 105510 4936 105562
rect 4960 105510 4990 105562
rect 4990 105510 5002 105562
rect 5002 105510 5016 105562
rect 5040 105510 5054 105562
rect 5054 105510 5066 105562
rect 5066 105510 5096 105562
rect 5120 105510 5130 105562
rect 5130 105510 5176 105562
rect 4880 105508 4936 105510
rect 4960 105508 5016 105510
rect 5040 105508 5096 105510
rect 5120 105508 5176 105510
rect 4220 105018 4276 105020
rect 4300 105018 4356 105020
rect 4380 105018 4436 105020
rect 4460 105018 4516 105020
rect 4220 104966 4266 105018
rect 4266 104966 4276 105018
rect 4300 104966 4330 105018
rect 4330 104966 4342 105018
rect 4342 104966 4356 105018
rect 4380 104966 4394 105018
rect 4394 104966 4406 105018
rect 4406 104966 4436 105018
rect 4460 104966 4470 105018
rect 4470 104966 4516 105018
rect 4220 104964 4276 104966
rect 4300 104964 4356 104966
rect 4380 104964 4436 104966
rect 4460 104964 4516 104966
rect 4880 104474 4936 104476
rect 4960 104474 5016 104476
rect 5040 104474 5096 104476
rect 5120 104474 5176 104476
rect 4880 104422 4926 104474
rect 4926 104422 4936 104474
rect 4960 104422 4990 104474
rect 4990 104422 5002 104474
rect 5002 104422 5016 104474
rect 5040 104422 5054 104474
rect 5054 104422 5066 104474
rect 5066 104422 5096 104474
rect 5120 104422 5130 104474
rect 5130 104422 5176 104474
rect 4880 104420 4936 104422
rect 4960 104420 5016 104422
rect 5040 104420 5096 104422
rect 5120 104420 5176 104422
rect 4220 103930 4276 103932
rect 4300 103930 4356 103932
rect 4380 103930 4436 103932
rect 4460 103930 4516 103932
rect 4220 103878 4266 103930
rect 4266 103878 4276 103930
rect 4300 103878 4330 103930
rect 4330 103878 4342 103930
rect 4342 103878 4356 103930
rect 4380 103878 4394 103930
rect 4394 103878 4406 103930
rect 4406 103878 4436 103930
rect 4460 103878 4470 103930
rect 4470 103878 4516 103930
rect 4220 103876 4276 103878
rect 4300 103876 4356 103878
rect 4380 103876 4436 103878
rect 4460 103876 4516 103878
rect 4880 103386 4936 103388
rect 4960 103386 5016 103388
rect 5040 103386 5096 103388
rect 5120 103386 5176 103388
rect 4880 103334 4926 103386
rect 4926 103334 4936 103386
rect 4960 103334 4990 103386
rect 4990 103334 5002 103386
rect 5002 103334 5016 103386
rect 5040 103334 5054 103386
rect 5054 103334 5066 103386
rect 5066 103334 5096 103386
rect 5120 103334 5130 103386
rect 5130 103334 5176 103386
rect 4880 103332 4936 103334
rect 4960 103332 5016 103334
rect 5040 103332 5096 103334
rect 5120 103332 5176 103334
rect 4220 102842 4276 102844
rect 4300 102842 4356 102844
rect 4380 102842 4436 102844
rect 4460 102842 4516 102844
rect 4220 102790 4266 102842
rect 4266 102790 4276 102842
rect 4300 102790 4330 102842
rect 4330 102790 4342 102842
rect 4342 102790 4356 102842
rect 4380 102790 4394 102842
rect 4394 102790 4406 102842
rect 4406 102790 4436 102842
rect 4460 102790 4470 102842
rect 4470 102790 4516 102842
rect 4220 102788 4276 102790
rect 4300 102788 4356 102790
rect 4380 102788 4436 102790
rect 4460 102788 4516 102790
rect 4880 102298 4936 102300
rect 4960 102298 5016 102300
rect 5040 102298 5096 102300
rect 5120 102298 5176 102300
rect 4880 102246 4926 102298
rect 4926 102246 4936 102298
rect 4960 102246 4990 102298
rect 4990 102246 5002 102298
rect 5002 102246 5016 102298
rect 5040 102246 5054 102298
rect 5054 102246 5066 102298
rect 5066 102246 5096 102298
rect 5120 102246 5130 102298
rect 5130 102246 5176 102298
rect 4880 102244 4936 102246
rect 4960 102244 5016 102246
rect 5040 102244 5096 102246
rect 5120 102244 5176 102246
rect 4220 101754 4276 101756
rect 4300 101754 4356 101756
rect 4380 101754 4436 101756
rect 4460 101754 4516 101756
rect 4220 101702 4266 101754
rect 4266 101702 4276 101754
rect 4300 101702 4330 101754
rect 4330 101702 4342 101754
rect 4342 101702 4356 101754
rect 4380 101702 4394 101754
rect 4394 101702 4406 101754
rect 4406 101702 4436 101754
rect 4460 101702 4470 101754
rect 4470 101702 4516 101754
rect 4220 101700 4276 101702
rect 4300 101700 4356 101702
rect 4380 101700 4436 101702
rect 4460 101700 4516 101702
rect 1214 101396 1216 101416
rect 1216 101396 1268 101416
rect 1268 101396 1270 101416
rect 1214 101360 1270 101396
rect 4880 101210 4936 101212
rect 4960 101210 5016 101212
rect 5040 101210 5096 101212
rect 5120 101210 5176 101212
rect 4880 101158 4926 101210
rect 4926 101158 4936 101210
rect 4960 101158 4990 101210
rect 4990 101158 5002 101210
rect 5002 101158 5016 101210
rect 5040 101158 5054 101210
rect 5054 101158 5066 101210
rect 5066 101158 5096 101210
rect 5120 101158 5130 101210
rect 5130 101158 5176 101210
rect 4880 101156 4936 101158
rect 4960 101156 5016 101158
rect 5040 101156 5096 101158
rect 5120 101156 5176 101158
rect 4220 100666 4276 100668
rect 4300 100666 4356 100668
rect 4380 100666 4436 100668
rect 4460 100666 4516 100668
rect 4220 100614 4266 100666
rect 4266 100614 4276 100666
rect 4300 100614 4330 100666
rect 4330 100614 4342 100666
rect 4342 100614 4356 100666
rect 4380 100614 4394 100666
rect 4394 100614 4406 100666
rect 4406 100614 4436 100666
rect 4460 100614 4470 100666
rect 4470 100614 4516 100666
rect 4220 100612 4276 100614
rect 4300 100612 4356 100614
rect 4380 100612 4436 100614
rect 4460 100612 4516 100614
rect 4880 100122 4936 100124
rect 4960 100122 5016 100124
rect 5040 100122 5096 100124
rect 5120 100122 5176 100124
rect 4880 100070 4926 100122
rect 4926 100070 4936 100122
rect 4960 100070 4990 100122
rect 4990 100070 5002 100122
rect 5002 100070 5016 100122
rect 5040 100070 5054 100122
rect 5054 100070 5066 100122
rect 5066 100070 5096 100122
rect 5120 100070 5130 100122
rect 5130 100070 5176 100122
rect 4880 100068 4936 100070
rect 4960 100068 5016 100070
rect 5040 100068 5096 100070
rect 5120 100068 5176 100070
rect 4220 99578 4276 99580
rect 4300 99578 4356 99580
rect 4380 99578 4436 99580
rect 4460 99578 4516 99580
rect 4220 99526 4266 99578
rect 4266 99526 4276 99578
rect 4300 99526 4330 99578
rect 4330 99526 4342 99578
rect 4342 99526 4356 99578
rect 4380 99526 4394 99578
rect 4394 99526 4406 99578
rect 4406 99526 4436 99578
rect 4460 99526 4470 99578
rect 4470 99526 4516 99578
rect 4220 99524 4276 99526
rect 4300 99524 4356 99526
rect 4380 99524 4436 99526
rect 4460 99524 4516 99526
rect 1398 99320 1454 99376
rect 4880 99034 4936 99036
rect 4960 99034 5016 99036
rect 5040 99034 5096 99036
rect 5120 99034 5176 99036
rect 4880 98982 4926 99034
rect 4926 98982 4936 99034
rect 4960 98982 4990 99034
rect 4990 98982 5002 99034
rect 5002 98982 5016 99034
rect 5040 98982 5054 99034
rect 5054 98982 5066 99034
rect 5066 98982 5096 99034
rect 5120 98982 5130 99034
rect 5130 98982 5176 99034
rect 4880 98980 4936 98982
rect 4960 98980 5016 98982
rect 5040 98980 5096 98982
rect 5120 98980 5176 98982
rect 1306 98640 1362 98696
rect 4220 98490 4276 98492
rect 4300 98490 4356 98492
rect 4380 98490 4436 98492
rect 4460 98490 4516 98492
rect 4220 98438 4266 98490
rect 4266 98438 4276 98490
rect 4300 98438 4330 98490
rect 4330 98438 4342 98490
rect 4342 98438 4356 98490
rect 4380 98438 4394 98490
rect 4394 98438 4406 98490
rect 4406 98438 4436 98490
rect 4460 98438 4470 98490
rect 4470 98438 4516 98490
rect 4220 98436 4276 98438
rect 4300 98436 4356 98438
rect 4380 98436 4436 98438
rect 4460 98436 4516 98438
rect 4880 97946 4936 97948
rect 4960 97946 5016 97948
rect 5040 97946 5096 97948
rect 5120 97946 5176 97948
rect 4880 97894 4926 97946
rect 4926 97894 4936 97946
rect 4960 97894 4990 97946
rect 4990 97894 5002 97946
rect 5002 97894 5016 97946
rect 5040 97894 5054 97946
rect 5054 97894 5066 97946
rect 5066 97894 5096 97946
rect 5120 97894 5130 97946
rect 5130 97894 5176 97946
rect 4880 97892 4936 97894
rect 4960 97892 5016 97894
rect 5040 97892 5096 97894
rect 5120 97892 5176 97894
rect 4220 97402 4276 97404
rect 4300 97402 4356 97404
rect 4380 97402 4436 97404
rect 4460 97402 4516 97404
rect 4220 97350 4266 97402
rect 4266 97350 4276 97402
rect 4300 97350 4330 97402
rect 4330 97350 4342 97402
rect 4342 97350 4356 97402
rect 4380 97350 4394 97402
rect 4394 97350 4406 97402
rect 4406 97350 4436 97402
rect 4460 97350 4470 97402
rect 4470 97350 4516 97402
rect 4220 97348 4276 97350
rect 4300 97348 4356 97350
rect 4380 97348 4436 97350
rect 4460 97348 4516 97350
rect 4880 96858 4936 96860
rect 4960 96858 5016 96860
rect 5040 96858 5096 96860
rect 5120 96858 5176 96860
rect 4880 96806 4926 96858
rect 4926 96806 4936 96858
rect 4960 96806 4990 96858
rect 4990 96806 5002 96858
rect 5002 96806 5016 96858
rect 5040 96806 5054 96858
rect 5054 96806 5066 96858
rect 5066 96806 5096 96858
rect 5120 96806 5130 96858
rect 5130 96806 5176 96858
rect 4880 96804 4936 96806
rect 4960 96804 5016 96806
rect 5040 96804 5096 96806
rect 5120 96804 5176 96806
rect 1306 96600 1362 96656
rect 4220 96314 4276 96316
rect 4300 96314 4356 96316
rect 4380 96314 4436 96316
rect 4460 96314 4516 96316
rect 4220 96262 4266 96314
rect 4266 96262 4276 96314
rect 4300 96262 4330 96314
rect 4330 96262 4342 96314
rect 4342 96262 4356 96314
rect 4380 96262 4394 96314
rect 4394 96262 4406 96314
rect 4406 96262 4436 96314
rect 4460 96262 4470 96314
rect 4470 96262 4516 96314
rect 4220 96260 4276 96262
rect 4300 96260 4356 96262
rect 4380 96260 4436 96262
rect 4460 96260 4516 96262
rect 1214 95956 1216 95976
rect 1216 95956 1268 95976
rect 1268 95956 1270 95976
rect 1214 95920 1270 95956
rect 4880 95770 4936 95772
rect 4960 95770 5016 95772
rect 5040 95770 5096 95772
rect 5120 95770 5176 95772
rect 4880 95718 4926 95770
rect 4926 95718 4936 95770
rect 4960 95718 4990 95770
rect 4990 95718 5002 95770
rect 5002 95718 5016 95770
rect 5040 95718 5054 95770
rect 5054 95718 5066 95770
rect 5066 95718 5096 95770
rect 5120 95718 5130 95770
rect 5130 95718 5176 95770
rect 4880 95716 4936 95718
rect 4960 95716 5016 95718
rect 5040 95716 5096 95718
rect 5120 95716 5176 95718
rect 4220 95226 4276 95228
rect 4300 95226 4356 95228
rect 4380 95226 4436 95228
rect 4460 95226 4516 95228
rect 4220 95174 4266 95226
rect 4266 95174 4276 95226
rect 4300 95174 4330 95226
rect 4330 95174 4342 95226
rect 4342 95174 4356 95226
rect 4380 95174 4394 95226
rect 4394 95174 4406 95226
rect 4406 95174 4436 95226
rect 4460 95174 4470 95226
rect 4470 95174 4516 95226
rect 4220 95172 4276 95174
rect 4300 95172 4356 95174
rect 4380 95172 4436 95174
rect 4460 95172 4516 95174
rect 4880 94682 4936 94684
rect 4960 94682 5016 94684
rect 5040 94682 5096 94684
rect 5120 94682 5176 94684
rect 4880 94630 4926 94682
rect 4926 94630 4936 94682
rect 4960 94630 4990 94682
rect 4990 94630 5002 94682
rect 5002 94630 5016 94682
rect 5040 94630 5054 94682
rect 5054 94630 5066 94682
rect 5066 94630 5096 94682
rect 5120 94630 5130 94682
rect 5130 94630 5176 94682
rect 4880 94628 4936 94630
rect 4960 94628 5016 94630
rect 5040 94628 5096 94630
rect 5120 94628 5176 94630
rect 4220 94138 4276 94140
rect 4300 94138 4356 94140
rect 4380 94138 4436 94140
rect 4460 94138 4516 94140
rect 4220 94086 4266 94138
rect 4266 94086 4276 94138
rect 4300 94086 4330 94138
rect 4330 94086 4342 94138
rect 4342 94086 4356 94138
rect 4380 94086 4394 94138
rect 4394 94086 4406 94138
rect 4406 94086 4436 94138
rect 4460 94086 4470 94138
rect 4470 94086 4516 94138
rect 4220 94084 4276 94086
rect 4300 94084 4356 94086
rect 4380 94084 4436 94086
rect 4460 94084 4516 94086
rect 1306 93880 1362 93936
rect 4880 93594 4936 93596
rect 4960 93594 5016 93596
rect 5040 93594 5096 93596
rect 5120 93594 5176 93596
rect 4880 93542 4926 93594
rect 4926 93542 4936 93594
rect 4960 93542 4990 93594
rect 4990 93542 5002 93594
rect 5002 93542 5016 93594
rect 5040 93542 5054 93594
rect 5054 93542 5066 93594
rect 5066 93542 5096 93594
rect 5120 93542 5130 93594
rect 5130 93542 5176 93594
rect 4880 93540 4936 93542
rect 4960 93540 5016 93542
rect 5040 93540 5096 93542
rect 5120 93540 5176 93542
rect 4220 93050 4276 93052
rect 4300 93050 4356 93052
rect 4380 93050 4436 93052
rect 4460 93050 4516 93052
rect 4220 92998 4266 93050
rect 4266 92998 4276 93050
rect 4300 92998 4330 93050
rect 4330 92998 4342 93050
rect 4342 92998 4356 93050
rect 4380 92998 4394 93050
rect 4394 92998 4406 93050
rect 4406 92998 4436 93050
rect 4460 92998 4470 93050
rect 4470 92998 4516 93050
rect 4220 92996 4276 92998
rect 4300 92996 4356 92998
rect 4380 92996 4436 92998
rect 4460 92996 4516 92998
rect 4880 92506 4936 92508
rect 4960 92506 5016 92508
rect 5040 92506 5096 92508
rect 5120 92506 5176 92508
rect 4880 92454 4926 92506
rect 4926 92454 4936 92506
rect 4960 92454 4990 92506
rect 4990 92454 5002 92506
rect 5002 92454 5016 92506
rect 5040 92454 5054 92506
rect 5054 92454 5066 92506
rect 5066 92454 5096 92506
rect 5120 92454 5130 92506
rect 5130 92454 5176 92506
rect 4880 92452 4936 92454
rect 4960 92452 5016 92454
rect 5040 92452 5096 92454
rect 5120 92452 5176 92454
rect 4220 91962 4276 91964
rect 4300 91962 4356 91964
rect 4380 91962 4436 91964
rect 4460 91962 4516 91964
rect 4220 91910 4266 91962
rect 4266 91910 4276 91962
rect 4300 91910 4330 91962
rect 4330 91910 4342 91962
rect 4342 91910 4356 91962
rect 4380 91910 4394 91962
rect 4394 91910 4406 91962
rect 4406 91910 4436 91962
rect 4460 91910 4470 91962
rect 4470 91910 4516 91962
rect 4220 91908 4276 91910
rect 4300 91908 4356 91910
rect 4380 91908 4436 91910
rect 4460 91908 4516 91910
rect 4880 91418 4936 91420
rect 4960 91418 5016 91420
rect 5040 91418 5096 91420
rect 5120 91418 5176 91420
rect 4880 91366 4926 91418
rect 4926 91366 4936 91418
rect 4960 91366 4990 91418
rect 4990 91366 5002 91418
rect 5002 91366 5016 91418
rect 5040 91366 5054 91418
rect 5054 91366 5066 91418
rect 5066 91366 5096 91418
rect 5120 91366 5130 91418
rect 5130 91366 5176 91418
rect 4880 91364 4936 91366
rect 4960 91364 5016 91366
rect 5040 91364 5096 91366
rect 5120 91364 5176 91366
rect 4220 90874 4276 90876
rect 4300 90874 4356 90876
rect 4380 90874 4436 90876
rect 4460 90874 4516 90876
rect 4220 90822 4266 90874
rect 4266 90822 4276 90874
rect 4300 90822 4330 90874
rect 4330 90822 4342 90874
rect 4342 90822 4356 90874
rect 4380 90822 4394 90874
rect 4394 90822 4406 90874
rect 4406 90822 4436 90874
rect 4460 90822 4470 90874
rect 4470 90822 4516 90874
rect 4220 90820 4276 90822
rect 4300 90820 4356 90822
rect 4380 90820 4436 90822
rect 4460 90820 4516 90822
rect 4880 90330 4936 90332
rect 4960 90330 5016 90332
rect 5040 90330 5096 90332
rect 5120 90330 5176 90332
rect 4880 90278 4926 90330
rect 4926 90278 4936 90330
rect 4960 90278 4990 90330
rect 4990 90278 5002 90330
rect 5002 90278 5016 90330
rect 5040 90278 5054 90330
rect 5054 90278 5066 90330
rect 5066 90278 5096 90330
rect 5120 90278 5130 90330
rect 5130 90278 5176 90330
rect 4880 90276 4936 90278
rect 4960 90276 5016 90278
rect 5040 90276 5096 90278
rect 5120 90276 5176 90278
rect 4220 89786 4276 89788
rect 4300 89786 4356 89788
rect 4380 89786 4436 89788
rect 4460 89786 4516 89788
rect 4220 89734 4266 89786
rect 4266 89734 4276 89786
rect 4300 89734 4330 89786
rect 4330 89734 4342 89786
rect 4342 89734 4356 89786
rect 4380 89734 4394 89786
rect 4394 89734 4406 89786
rect 4406 89734 4436 89786
rect 4460 89734 4470 89786
rect 4470 89734 4516 89786
rect 4220 89732 4276 89734
rect 4300 89732 4356 89734
rect 4380 89732 4436 89734
rect 4460 89732 4516 89734
rect 4880 89242 4936 89244
rect 4960 89242 5016 89244
rect 5040 89242 5096 89244
rect 5120 89242 5176 89244
rect 4880 89190 4926 89242
rect 4926 89190 4936 89242
rect 4960 89190 4990 89242
rect 4990 89190 5002 89242
rect 5002 89190 5016 89242
rect 5040 89190 5054 89242
rect 5054 89190 5066 89242
rect 5066 89190 5096 89242
rect 5120 89190 5130 89242
rect 5130 89190 5176 89242
rect 4880 89188 4936 89190
rect 4960 89188 5016 89190
rect 5040 89188 5096 89190
rect 5120 89188 5176 89190
rect 4220 88698 4276 88700
rect 4300 88698 4356 88700
rect 4380 88698 4436 88700
rect 4460 88698 4516 88700
rect 4220 88646 4266 88698
rect 4266 88646 4276 88698
rect 4300 88646 4330 88698
rect 4330 88646 4342 88698
rect 4342 88646 4356 88698
rect 4380 88646 4394 88698
rect 4394 88646 4406 88698
rect 4406 88646 4436 88698
rect 4460 88646 4470 88698
rect 4470 88646 4516 88698
rect 4220 88644 4276 88646
rect 4300 88644 4356 88646
rect 4380 88644 4436 88646
rect 4460 88644 4516 88646
rect 4880 88154 4936 88156
rect 4960 88154 5016 88156
rect 5040 88154 5096 88156
rect 5120 88154 5176 88156
rect 4880 88102 4926 88154
rect 4926 88102 4936 88154
rect 4960 88102 4990 88154
rect 4990 88102 5002 88154
rect 5002 88102 5016 88154
rect 5040 88102 5054 88154
rect 5054 88102 5066 88154
rect 5066 88102 5096 88154
rect 5120 88102 5130 88154
rect 5130 88102 5176 88154
rect 4880 88100 4936 88102
rect 4960 88100 5016 88102
rect 5040 88100 5096 88102
rect 5120 88100 5176 88102
rect 4220 87610 4276 87612
rect 4300 87610 4356 87612
rect 4380 87610 4436 87612
rect 4460 87610 4516 87612
rect 4220 87558 4266 87610
rect 4266 87558 4276 87610
rect 4300 87558 4330 87610
rect 4330 87558 4342 87610
rect 4342 87558 4356 87610
rect 4380 87558 4394 87610
rect 4394 87558 4406 87610
rect 4406 87558 4436 87610
rect 4460 87558 4470 87610
rect 4470 87558 4516 87610
rect 4220 87556 4276 87558
rect 4300 87556 4356 87558
rect 4380 87556 4436 87558
rect 4460 87556 4516 87558
rect 4880 87066 4936 87068
rect 4960 87066 5016 87068
rect 5040 87066 5096 87068
rect 5120 87066 5176 87068
rect 4880 87014 4926 87066
rect 4926 87014 4936 87066
rect 4960 87014 4990 87066
rect 4990 87014 5002 87066
rect 5002 87014 5016 87066
rect 5040 87014 5054 87066
rect 5054 87014 5066 87066
rect 5066 87014 5096 87066
rect 5120 87014 5130 87066
rect 5130 87014 5176 87066
rect 4880 87012 4936 87014
rect 4960 87012 5016 87014
rect 5040 87012 5096 87014
rect 5120 87012 5176 87014
rect 4220 86522 4276 86524
rect 4300 86522 4356 86524
rect 4380 86522 4436 86524
rect 4460 86522 4516 86524
rect 4220 86470 4266 86522
rect 4266 86470 4276 86522
rect 4300 86470 4330 86522
rect 4330 86470 4342 86522
rect 4342 86470 4356 86522
rect 4380 86470 4394 86522
rect 4394 86470 4406 86522
rect 4406 86470 4436 86522
rect 4460 86470 4470 86522
rect 4470 86470 4516 86522
rect 4220 86468 4276 86470
rect 4300 86468 4356 86470
rect 4380 86468 4436 86470
rect 4460 86468 4516 86470
rect 4880 85978 4936 85980
rect 4960 85978 5016 85980
rect 5040 85978 5096 85980
rect 5120 85978 5176 85980
rect 4880 85926 4926 85978
rect 4926 85926 4936 85978
rect 4960 85926 4990 85978
rect 4990 85926 5002 85978
rect 5002 85926 5016 85978
rect 5040 85926 5054 85978
rect 5054 85926 5066 85978
rect 5066 85926 5096 85978
rect 5120 85926 5130 85978
rect 5130 85926 5176 85978
rect 4880 85924 4936 85926
rect 4960 85924 5016 85926
rect 5040 85924 5096 85926
rect 5120 85924 5176 85926
rect 4220 85434 4276 85436
rect 4300 85434 4356 85436
rect 4380 85434 4436 85436
rect 4460 85434 4516 85436
rect 4220 85382 4266 85434
rect 4266 85382 4276 85434
rect 4300 85382 4330 85434
rect 4330 85382 4342 85434
rect 4342 85382 4356 85434
rect 4380 85382 4394 85434
rect 4394 85382 4406 85434
rect 4406 85382 4436 85434
rect 4460 85382 4470 85434
rect 4470 85382 4516 85434
rect 4220 85380 4276 85382
rect 4300 85380 4356 85382
rect 4380 85380 4436 85382
rect 4460 85380 4516 85382
rect 4880 84890 4936 84892
rect 4960 84890 5016 84892
rect 5040 84890 5096 84892
rect 5120 84890 5176 84892
rect 4880 84838 4926 84890
rect 4926 84838 4936 84890
rect 4960 84838 4990 84890
rect 4990 84838 5002 84890
rect 5002 84838 5016 84890
rect 5040 84838 5054 84890
rect 5054 84838 5066 84890
rect 5066 84838 5096 84890
rect 5120 84838 5130 84890
rect 5130 84838 5176 84890
rect 4880 84836 4936 84838
rect 4960 84836 5016 84838
rect 5040 84836 5096 84838
rect 5120 84836 5176 84838
rect 4220 84346 4276 84348
rect 4300 84346 4356 84348
rect 4380 84346 4436 84348
rect 4460 84346 4516 84348
rect 4220 84294 4266 84346
rect 4266 84294 4276 84346
rect 4300 84294 4330 84346
rect 4330 84294 4342 84346
rect 4342 84294 4356 84346
rect 4380 84294 4394 84346
rect 4394 84294 4406 84346
rect 4406 84294 4436 84346
rect 4460 84294 4470 84346
rect 4470 84294 4516 84346
rect 4220 84292 4276 84294
rect 4300 84292 4356 84294
rect 4380 84292 4436 84294
rect 4460 84292 4516 84294
rect 4880 83802 4936 83804
rect 4960 83802 5016 83804
rect 5040 83802 5096 83804
rect 5120 83802 5176 83804
rect 4880 83750 4926 83802
rect 4926 83750 4936 83802
rect 4960 83750 4990 83802
rect 4990 83750 5002 83802
rect 5002 83750 5016 83802
rect 5040 83750 5054 83802
rect 5054 83750 5066 83802
rect 5066 83750 5096 83802
rect 5120 83750 5130 83802
rect 5130 83750 5176 83802
rect 4880 83748 4936 83750
rect 4960 83748 5016 83750
rect 5040 83748 5096 83750
rect 5120 83748 5176 83750
rect 4220 83258 4276 83260
rect 4300 83258 4356 83260
rect 4380 83258 4436 83260
rect 4460 83258 4516 83260
rect 4220 83206 4266 83258
rect 4266 83206 4276 83258
rect 4300 83206 4330 83258
rect 4330 83206 4342 83258
rect 4342 83206 4356 83258
rect 4380 83206 4394 83258
rect 4394 83206 4406 83258
rect 4406 83206 4436 83258
rect 4460 83206 4470 83258
rect 4470 83206 4516 83258
rect 4220 83204 4276 83206
rect 4300 83204 4356 83206
rect 4380 83204 4436 83206
rect 4460 83204 4516 83206
rect 4880 82714 4936 82716
rect 4960 82714 5016 82716
rect 5040 82714 5096 82716
rect 5120 82714 5176 82716
rect 4880 82662 4926 82714
rect 4926 82662 4936 82714
rect 4960 82662 4990 82714
rect 4990 82662 5002 82714
rect 5002 82662 5016 82714
rect 5040 82662 5054 82714
rect 5054 82662 5066 82714
rect 5066 82662 5096 82714
rect 5120 82662 5130 82714
rect 5130 82662 5176 82714
rect 4880 82660 4936 82662
rect 4960 82660 5016 82662
rect 5040 82660 5096 82662
rect 5120 82660 5176 82662
rect 4220 82170 4276 82172
rect 4300 82170 4356 82172
rect 4380 82170 4436 82172
rect 4460 82170 4516 82172
rect 4220 82118 4266 82170
rect 4266 82118 4276 82170
rect 4300 82118 4330 82170
rect 4330 82118 4342 82170
rect 4342 82118 4356 82170
rect 4380 82118 4394 82170
rect 4394 82118 4406 82170
rect 4406 82118 4436 82170
rect 4460 82118 4470 82170
rect 4470 82118 4516 82170
rect 4220 82116 4276 82118
rect 4300 82116 4356 82118
rect 4380 82116 4436 82118
rect 4460 82116 4516 82118
rect 4880 81626 4936 81628
rect 4960 81626 5016 81628
rect 5040 81626 5096 81628
rect 5120 81626 5176 81628
rect 4880 81574 4926 81626
rect 4926 81574 4936 81626
rect 4960 81574 4990 81626
rect 4990 81574 5002 81626
rect 5002 81574 5016 81626
rect 5040 81574 5054 81626
rect 5054 81574 5066 81626
rect 5066 81574 5096 81626
rect 5120 81574 5130 81626
rect 5130 81574 5176 81626
rect 4880 81572 4936 81574
rect 4960 81572 5016 81574
rect 5040 81572 5096 81574
rect 5120 81572 5176 81574
rect 4220 81082 4276 81084
rect 4300 81082 4356 81084
rect 4380 81082 4436 81084
rect 4460 81082 4516 81084
rect 4220 81030 4266 81082
rect 4266 81030 4276 81082
rect 4300 81030 4330 81082
rect 4330 81030 4342 81082
rect 4342 81030 4356 81082
rect 4380 81030 4394 81082
rect 4394 81030 4406 81082
rect 4406 81030 4436 81082
rect 4460 81030 4470 81082
rect 4470 81030 4516 81082
rect 4220 81028 4276 81030
rect 4300 81028 4356 81030
rect 4380 81028 4436 81030
rect 4460 81028 4516 81030
rect 4880 80538 4936 80540
rect 4960 80538 5016 80540
rect 5040 80538 5096 80540
rect 5120 80538 5176 80540
rect 4880 80486 4926 80538
rect 4926 80486 4936 80538
rect 4960 80486 4990 80538
rect 4990 80486 5002 80538
rect 5002 80486 5016 80538
rect 5040 80486 5054 80538
rect 5054 80486 5066 80538
rect 5066 80486 5096 80538
rect 5120 80486 5130 80538
rect 5130 80486 5176 80538
rect 4880 80484 4936 80486
rect 4960 80484 5016 80486
rect 5040 80484 5096 80486
rect 5120 80484 5176 80486
rect 4220 79994 4276 79996
rect 4300 79994 4356 79996
rect 4380 79994 4436 79996
rect 4460 79994 4516 79996
rect 4220 79942 4266 79994
rect 4266 79942 4276 79994
rect 4300 79942 4330 79994
rect 4330 79942 4342 79994
rect 4342 79942 4356 79994
rect 4380 79942 4394 79994
rect 4394 79942 4406 79994
rect 4406 79942 4436 79994
rect 4460 79942 4470 79994
rect 4470 79942 4516 79994
rect 4220 79940 4276 79942
rect 4300 79940 4356 79942
rect 4380 79940 4436 79942
rect 4460 79940 4516 79942
rect 4880 79450 4936 79452
rect 4960 79450 5016 79452
rect 5040 79450 5096 79452
rect 5120 79450 5176 79452
rect 4880 79398 4926 79450
rect 4926 79398 4936 79450
rect 4960 79398 4990 79450
rect 4990 79398 5002 79450
rect 5002 79398 5016 79450
rect 5040 79398 5054 79450
rect 5054 79398 5066 79450
rect 5066 79398 5096 79450
rect 5120 79398 5130 79450
rect 5130 79398 5176 79450
rect 4880 79396 4936 79398
rect 4960 79396 5016 79398
rect 5040 79396 5096 79398
rect 5120 79396 5176 79398
rect 4220 78906 4276 78908
rect 4300 78906 4356 78908
rect 4380 78906 4436 78908
rect 4460 78906 4516 78908
rect 4220 78854 4266 78906
rect 4266 78854 4276 78906
rect 4300 78854 4330 78906
rect 4330 78854 4342 78906
rect 4342 78854 4356 78906
rect 4380 78854 4394 78906
rect 4394 78854 4406 78906
rect 4406 78854 4436 78906
rect 4460 78854 4470 78906
rect 4470 78854 4516 78906
rect 4220 78852 4276 78854
rect 4300 78852 4356 78854
rect 4380 78852 4436 78854
rect 4460 78852 4516 78854
rect 4880 78362 4936 78364
rect 4960 78362 5016 78364
rect 5040 78362 5096 78364
rect 5120 78362 5176 78364
rect 4880 78310 4926 78362
rect 4926 78310 4936 78362
rect 4960 78310 4990 78362
rect 4990 78310 5002 78362
rect 5002 78310 5016 78362
rect 5040 78310 5054 78362
rect 5054 78310 5066 78362
rect 5066 78310 5096 78362
rect 5120 78310 5130 78362
rect 5130 78310 5176 78362
rect 4880 78308 4936 78310
rect 4960 78308 5016 78310
rect 5040 78308 5096 78310
rect 5120 78308 5176 78310
rect 1306 78240 1362 78296
rect 4220 77818 4276 77820
rect 4300 77818 4356 77820
rect 4380 77818 4436 77820
rect 4460 77818 4516 77820
rect 4220 77766 4266 77818
rect 4266 77766 4276 77818
rect 4300 77766 4330 77818
rect 4330 77766 4342 77818
rect 4342 77766 4356 77818
rect 4380 77766 4394 77818
rect 4394 77766 4406 77818
rect 4406 77766 4436 77818
rect 4460 77766 4470 77818
rect 4470 77766 4516 77818
rect 4220 77764 4276 77766
rect 4300 77764 4356 77766
rect 4380 77764 4436 77766
rect 4460 77764 4516 77766
rect 1306 77560 1362 77616
rect 4880 77274 4936 77276
rect 4960 77274 5016 77276
rect 5040 77274 5096 77276
rect 5120 77274 5176 77276
rect 4880 77222 4926 77274
rect 4926 77222 4936 77274
rect 4960 77222 4990 77274
rect 4990 77222 5002 77274
rect 5002 77222 5016 77274
rect 5040 77222 5054 77274
rect 5054 77222 5066 77274
rect 5066 77222 5096 77274
rect 5120 77222 5130 77274
rect 5130 77222 5176 77274
rect 4880 77220 4936 77222
rect 4960 77220 5016 77222
rect 5040 77220 5096 77222
rect 5120 77220 5176 77222
rect 1214 76880 1270 76936
rect 4220 76730 4276 76732
rect 4300 76730 4356 76732
rect 4380 76730 4436 76732
rect 4460 76730 4516 76732
rect 4220 76678 4266 76730
rect 4266 76678 4276 76730
rect 4300 76678 4330 76730
rect 4330 76678 4342 76730
rect 4342 76678 4356 76730
rect 4380 76678 4394 76730
rect 4394 76678 4406 76730
rect 4406 76678 4436 76730
rect 4460 76678 4470 76730
rect 4470 76678 4516 76730
rect 4220 76676 4276 76678
rect 4300 76676 4356 76678
rect 4380 76676 4436 76678
rect 4460 76676 4516 76678
rect 1214 76200 1270 76256
rect 4880 76186 4936 76188
rect 4960 76186 5016 76188
rect 5040 76186 5096 76188
rect 5120 76186 5176 76188
rect 4880 76134 4926 76186
rect 4926 76134 4936 76186
rect 4960 76134 4990 76186
rect 4990 76134 5002 76186
rect 5002 76134 5016 76186
rect 5040 76134 5054 76186
rect 5054 76134 5066 76186
rect 5066 76134 5096 76186
rect 5120 76134 5130 76186
rect 5130 76134 5176 76186
rect 4880 76132 4936 76134
rect 4960 76132 5016 76134
rect 5040 76132 5096 76134
rect 5120 76132 5176 76134
rect 4220 75642 4276 75644
rect 4300 75642 4356 75644
rect 4380 75642 4436 75644
rect 4460 75642 4516 75644
rect 4220 75590 4266 75642
rect 4266 75590 4276 75642
rect 4300 75590 4330 75642
rect 4330 75590 4342 75642
rect 4342 75590 4356 75642
rect 4380 75590 4394 75642
rect 4394 75590 4406 75642
rect 4406 75590 4436 75642
rect 4460 75590 4470 75642
rect 4470 75590 4516 75642
rect 4220 75588 4276 75590
rect 4300 75588 4356 75590
rect 4380 75588 4436 75590
rect 4460 75588 4516 75590
rect 1398 75520 1454 75576
rect 5538 75520 5594 75576
rect 4880 75098 4936 75100
rect 4960 75098 5016 75100
rect 5040 75098 5096 75100
rect 5120 75098 5176 75100
rect 4880 75046 4926 75098
rect 4926 75046 4936 75098
rect 4960 75046 4990 75098
rect 4990 75046 5002 75098
rect 5002 75046 5016 75098
rect 5040 75046 5054 75098
rect 5054 75046 5066 75098
rect 5066 75046 5096 75098
rect 5120 75046 5130 75098
rect 5130 75046 5176 75098
rect 4880 75044 4936 75046
rect 4960 75044 5016 75046
rect 5040 75044 5096 75046
rect 5120 75044 5176 75046
rect 1306 74840 1362 74896
rect 4220 74554 4276 74556
rect 4300 74554 4356 74556
rect 4380 74554 4436 74556
rect 4460 74554 4516 74556
rect 4220 74502 4266 74554
rect 4266 74502 4276 74554
rect 4300 74502 4330 74554
rect 4330 74502 4342 74554
rect 4342 74502 4356 74554
rect 4380 74502 4394 74554
rect 4394 74502 4406 74554
rect 4406 74502 4436 74554
rect 4460 74502 4470 74554
rect 4470 74502 4516 74554
rect 4220 74500 4276 74502
rect 4300 74500 4356 74502
rect 4380 74500 4436 74502
rect 4460 74500 4516 74502
rect 1214 74180 1270 74216
rect 1214 74160 1216 74180
rect 1216 74160 1268 74180
rect 1268 74160 1270 74180
rect 1306 73480 1362 73536
rect 1490 72800 1546 72856
rect 1306 72120 1362 72176
rect 4880 74010 4936 74012
rect 4960 74010 5016 74012
rect 5040 74010 5096 74012
rect 5120 74010 5176 74012
rect 4880 73958 4926 74010
rect 4926 73958 4936 74010
rect 4960 73958 4990 74010
rect 4990 73958 5002 74010
rect 5002 73958 5016 74010
rect 5040 73958 5054 74010
rect 5054 73958 5066 74010
rect 5066 73958 5096 74010
rect 5120 73958 5130 74010
rect 5130 73958 5176 74010
rect 4880 73956 4936 73958
rect 4960 73956 5016 73958
rect 5040 73956 5096 73958
rect 5120 73956 5176 73958
rect 4220 73466 4276 73468
rect 4300 73466 4356 73468
rect 4380 73466 4436 73468
rect 4460 73466 4516 73468
rect 4220 73414 4266 73466
rect 4266 73414 4276 73466
rect 4300 73414 4330 73466
rect 4330 73414 4342 73466
rect 4342 73414 4356 73466
rect 4380 73414 4394 73466
rect 4394 73414 4406 73466
rect 4406 73414 4436 73466
rect 4460 73414 4470 73466
rect 4470 73414 4516 73466
rect 4220 73412 4276 73414
rect 4300 73412 4356 73414
rect 4380 73412 4436 73414
rect 4460 73412 4516 73414
rect 4880 72922 4936 72924
rect 4960 72922 5016 72924
rect 5040 72922 5096 72924
rect 5120 72922 5176 72924
rect 4880 72870 4926 72922
rect 4926 72870 4936 72922
rect 4960 72870 4990 72922
rect 4990 72870 5002 72922
rect 5002 72870 5016 72922
rect 5040 72870 5054 72922
rect 5054 72870 5066 72922
rect 5066 72870 5096 72922
rect 5120 72870 5130 72922
rect 5130 72870 5176 72922
rect 4880 72868 4936 72870
rect 4960 72868 5016 72870
rect 5040 72868 5096 72870
rect 5120 72868 5176 72870
rect 4220 72378 4276 72380
rect 4300 72378 4356 72380
rect 4380 72378 4436 72380
rect 4460 72378 4516 72380
rect 4220 72326 4266 72378
rect 4266 72326 4276 72378
rect 4300 72326 4330 72378
rect 4330 72326 4342 72378
rect 4342 72326 4356 72378
rect 4380 72326 4394 72378
rect 4394 72326 4406 72378
rect 4406 72326 4436 72378
rect 4460 72326 4470 72378
rect 4470 72326 4516 72378
rect 4220 72324 4276 72326
rect 4300 72324 4356 72326
rect 4380 72324 4436 72326
rect 4460 72324 4516 72326
rect 4880 71834 4936 71836
rect 4960 71834 5016 71836
rect 5040 71834 5096 71836
rect 5120 71834 5176 71836
rect 4880 71782 4926 71834
rect 4926 71782 4936 71834
rect 4960 71782 4990 71834
rect 4990 71782 5002 71834
rect 5002 71782 5016 71834
rect 5040 71782 5054 71834
rect 5054 71782 5066 71834
rect 5066 71782 5096 71834
rect 5120 71782 5130 71834
rect 5130 71782 5176 71834
rect 4880 71780 4936 71782
rect 4960 71780 5016 71782
rect 5040 71780 5096 71782
rect 5120 71780 5176 71782
rect 1214 71440 1270 71496
rect 1306 70760 1362 70816
rect 4220 71290 4276 71292
rect 4300 71290 4356 71292
rect 4380 71290 4436 71292
rect 4460 71290 4516 71292
rect 4220 71238 4266 71290
rect 4266 71238 4276 71290
rect 4300 71238 4330 71290
rect 4330 71238 4342 71290
rect 4342 71238 4356 71290
rect 4380 71238 4394 71290
rect 4394 71238 4406 71290
rect 4406 71238 4436 71290
rect 4460 71238 4470 71290
rect 4470 71238 4516 71290
rect 4220 71236 4276 71238
rect 4300 71236 4356 71238
rect 4380 71236 4436 71238
rect 4460 71236 4516 71238
rect 4880 70746 4936 70748
rect 4960 70746 5016 70748
rect 5040 70746 5096 70748
rect 5120 70746 5176 70748
rect 4880 70694 4926 70746
rect 4926 70694 4936 70746
rect 4960 70694 4990 70746
rect 4990 70694 5002 70746
rect 5002 70694 5016 70746
rect 5040 70694 5054 70746
rect 5054 70694 5066 70746
rect 5066 70694 5096 70746
rect 5120 70694 5130 70746
rect 5130 70694 5176 70746
rect 4880 70692 4936 70694
rect 4960 70692 5016 70694
rect 5040 70692 5096 70694
rect 5120 70692 5176 70694
rect 4220 70202 4276 70204
rect 4300 70202 4356 70204
rect 4380 70202 4436 70204
rect 4460 70202 4516 70204
rect 4220 70150 4266 70202
rect 4266 70150 4276 70202
rect 4300 70150 4330 70202
rect 4330 70150 4342 70202
rect 4342 70150 4356 70202
rect 4380 70150 4394 70202
rect 4394 70150 4406 70202
rect 4406 70150 4436 70202
rect 4460 70150 4470 70202
rect 4470 70150 4516 70202
rect 4220 70148 4276 70150
rect 4300 70148 4356 70150
rect 4380 70148 4436 70150
rect 4460 70148 4516 70150
rect 2226 70080 2282 70136
rect 4880 69658 4936 69660
rect 4960 69658 5016 69660
rect 5040 69658 5096 69660
rect 5120 69658 5176 69660
rect 4880 69606 4926 69658
rect 4926 69606 4936 69658
rect 4960 69606 4990 69658
rect 4990 69606 5002 69658
rect 5002 69606 5016 69658
rect 5040 69606 5054 69658
rect 5054 69606 5066 69658
rect 5066 69606 5096 69658
rect 5120 69606 5130 69658
rect 5130 69606 5176 69658
rect 4880 69604 4936 69606
rect 4960 69604 5016 69606
rect 5040 69604 5096 69606
rect 5120 69604 5176 69606
rect 1306 69400 1362 69456
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 1214 68740 1270 68776
rect 1214 68720 1216 68740
rect 1216 68720 1268 68740
rect 1268 68720 1270 68740
rect 4880 68570 4936 68572
rect 4960 68570 5016 68572
rect 5040 68570 5096 68572
rect 5120 68570 5176 68572
rect 4880 68518 4926 68570
rect 4926 68518 4936 68570
rect 4960 68518 4990 68570
rect 4990 68518 5002 68570
rect 5002 68518 5016 68570
rect 5040 68518 5054 68570
rect 5054 68518 5066 68570
rect 5066 68518 5096 68570
rect 5120 68518 5130 68570
rect 5130 68518 5176 68570
rect 4880 68516 4936 68518
rect 4960 68516 5016 68518
rect 5040 68516 5096 68518
rect 5120 68516 5176 68518
rect 1306 68040 1362 68096
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 1122 67360 1178 67416
rect 846 66816 902 66872
rect 846 65900 848 65920
rect 848 65900 900 65920
rect 900 65900 902 65920
rect 846 65864 902 65900
rect 846 65456 902 65512
rect 1398 64640 1454 64696
rect 846 64096 902 64152
rect 846 63452 848 63472
rect 848 63452 900 63472
rect 900 63452 902 63472
rect 846 63416 902 63452
rect 846 62756 902 62792
rect 846 62736 848 62756
rect 848 62736 900 62756
rect 900 62736 902 62756
rect 1490 61920 1546 61976
rect 4880 67482 4936 67484
rect 4960 67482 5016 67484
rect 5040 67482 5096 67484
rect 5120 67482 5176 67484
rect 4880 67430 4926 67482
rect 4926 67430 4936 67482
rect 4960 67430 4990 67482
rect 4990 67430 5002 67482
rect 5002 67430 5016 67482
rect 5040 67430 5054 67482
rect 5054 67430 5066 67482
rect 5066 67430 5096 67482
rect 5120 67430 5130 67482
rect 5130 67430 5176 67482
rect 4880 67428 4936 67430
rect 4960 67428 5016 67430
rect 5040 67428 5096 67430
rect 5120 67428 5176 67430
rect 8022 67224 8078 67280
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 8390 101224 8446 101280
rect 8390 99456 8446 99512
rect 8390 98368 8446 98424
rect 8390 96736 8446 96792
rect 8390 95648 8446 95704
rect 8390 93880 8446 93936
rect 8942 69672 8998 69728
rect 8850 69536 8906 69592
rect 8206 67360 8262 67416
rect 9218 69808 9274 69864
rect 36082 124208 36138 124264
rect 37738 124208 37794 124264
rect 41326 124208 41382 124264
rect 77298 126404 77354 126440
rect 77298 126384 77300 126404
rect 77300 126384 77352 126404
rect 77352 126384 77354 126404
rect 45190 125976 45246 126032
rect 56782 125976 56838 126032
rect 61842 125704 61898 125760
rect 49698 125568 49754 125624
rect 59358 125568 59414 125624
rect 63958 125568 64014 125624
rect 64418 125160 64474 125216
rect 66320 126234 66376 126236
rect 66400 126234 66456 126236
rect 66480 126234 66536 126236
rect 66560 126234 66616 126236
rect 66320 126182 66366 126234
rect 66366 126182 66376 126234
rect 66400 126182 66430 126234
rect 66430 126182 66442 126234
rect 66442 126182 66456 126234
rect 66480 126182 66494 126234
rect 66494 126182 66506 126234
rect 66506 126182 66536 126234
rect 66560 126182 66570 126234
rect 66570 126182 66616 126234
rect 66320 126180 66376 126182
rect 66400 126180 66456 126182
rect 66480 126180 66536 126182
rect 66560 126180 66616 126182
rect 48502 124208 48558 124264
rect 66074 124208 66130 124264
rect 68558 124208 68614 124264
rect 71410 124208 71466 124264
rect 42338 124072 42394 124128
rect 86314 123936 86370 123992
rect 97040 126234 97096 126236
rect 97120 126234 97176 126236
rect 97200 126234 97256 126236
rect 97280 126234 97336 126236
rect 97040 126182 97086 126234
rect 97086 126182 97096 126234
rect 97120 126182 97150 126234
rect 97150 126182 97162 126234
rect 97162 126182 97176 126234
rect 97200 126182 97214 126234
rect 97214 126182 97226 126234
rect 97226 126182 97256 126234
rect 97280 126182 97290 126234
rect 97290 126182 97336 126234
rect 97040 126180 97096 126182
rect 97120 126180 97176 126182
rect 97200 126180 97256 126182
rect 97280 126180 97336 126182
rect 87326 123800 87382 123856
rect 96066 123800 96122 123856
rect 37462 69808 37518 69864
rect 38658 69808 38714 69864
rect 39762 69828 39818 69864
rect 39762 69808 39764 69828
rect 39764 69808 39816 69828
rect 39816 69808 39818 69828
rect 23294 69536 23350 69592
rect 23478 69536 23534 69592
rect 24674 69536 24730 69592
rect 25778 69536 25834 69592
rect 26974 69536 27030 69592
rect 28078 69536 28134 69592
rect 30470 69536 30526 69592
rect 31758 69536 31814 69592
rect 32862 69556 32918 69592
rect 32862 69536 32864 69556
rect 32864 69536 32916 69556
rect 32916 69536 32918 69556
rect 9402 69400 9458 69456
rect 23294 69264 23350 69320
rect 29550 69264 29606 69320
rect 33966 69536 34022 69592
rect 35162 69536 35218 69592
rect 36358 69536 36414 69592
rect 9126 67088 9182 67144
rect 8114 66680 8170 66736
rect 4880 66394 4936 66396
rect 4960 66394 5016 66396
rect 5040 66394 5096 66396
rect 5120 66394 5176 66396
rect 4880 66342 4926 66394
rect 4926 66342 4936 66394
rect 4960 66342 4990 66394
rect 4990 66342 5002 66394
rect 5002 66342 5016 66394
rect 5040 66342 5054 66394
rect 5054 66342 5066 66394
rect 5066 66342 5096 66394
rect 5120 66342 5130 66394
rect 5130 66342 5176 66394
rect 4880 66340 4936 66342
rect 4960 66340 5016 66342
rect 5040 66340 5096 66342
rect 5120 66340 5176 66342
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 4880 65306 4936 65308
rect 4960 65306 5016 65308
rect 5040 65306 5096 65308
rect 5120 65306 5176 65308
rect 4880 65254 4926 65306
rect 4926 65254 4936 65306
rect 4960 65254 4990 65306
rect 4990 65254 5002 65306
rect 5002 65254 5016 65306
rect 5040 65254 5054 65306
rect 5054 65254 5066 65306
rect 5066 65254 5096 65306
rect 5120 65254 5130 65306
rect 5130 65254 5176 65306
rect 4880 65252 4936 65254
rect 4960 65252 5016 65254
rect 5040 65252 5096 65254
rect 5120 65252 5176 65254
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 4880 64218 4936 64220
rect 4960 64218 5016 64220
rect 5040 64218 5096 64220
rect 5120 64218 5176 64220
rect 4880 64166 4926 64218
rect 4926 64166 4936 64218
rect 4960 64166 4990 64218
rect 4990 64166 5002 64218
rect 5002 64166 5016 64218
rect 5040 64166 5054 64218
rect 5054 64166 5066 64218
rect 5066 64166 5096 64218
rect 5120 64166 5130 64218
rect 5130 64166 5176 64218
rect 4880 64164 4936 64166
rect 4960 64164 5016 64166
rect 5040 64164 5096 64166
rect 5120 64164 5176 64166
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 4880 63130 4936 63132
rect 4960 63130 5016 63132
rect 5040 63130 5096 63132
rect 5120 63130 5176 63132
rect 4880 63078 4926 63130
rect 4926 63078 4936 63130
rect 4960 63078 4990 63130
rect 4990 63078 5002 63130
rect 5002 63078 5016 63130
rect 5040 63078 5054 63130
rect 5054 63078 5066 63130
rect 5066 63078 5096 63130
rect 5120 63078 5130 63130
rect 5130 63078 5176 63130
rect 4880 63076 4936 63078
rect 4960 63076 5016 63078
rect 5040 63076 5096 63078
rect 5120 63076 5176 63078
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 4880 62042 4936 62044
rect 4960 62042 5016 62044
rect 5040 62042 5096 62044
rect 5120 62042 5176 62044
rect 4880 61990 4926 62042
rect 4926 61990 4936 62042
rect 4960 61990 4990 62042
rect 4990 61990 5002 62042
rect 5002 61990 5016 62042
rect 5040 61990 5054 62042
rect 5054 61990 5066 62042
rect 5066 61990 5096 62042
rect 5120 61990 5130 62042
rect 5130 61990 5176 62042
rect 4880 61988 4936 61990
rect 4960 61988 5016 61990
rect 5040 61988 5096 61990
rect 5120 61988 5176 61990
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 1306 61240 1362 61296
rect 4880 60954 4936 60956
rect 4960 60954 5016 60956
rect 5040 60954 5096 60956
rect 5120 60954 5176 60956
rect 4880 60902 4926 60954
rect 4926 60902 4936 60954
rect 4960 60902 4990 60954
rect 4990 60902 5002 60954
rect 5002 60902 5016 60954
rect 5040 60902 5054 60954
rect 5054 60902 5066 60954
rect 5066 60902 5096 60954
rect 5120 60902 5130 60954
rect 5130 60902 5176 60954
rect 4880 60900 4936 60902
rect 4960 60900 5016 60902
rect 5040 60900 5096 60902
rect 5120 60900 5176 60902
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 4880 59866 4936 59868
rect 4960 59866 5016 59868
rect 5040 59866 5096 59868
rect 5120 59866 5176 59868
rect 4880 59814 4926 59866
rect 4926 59814 4936 59866
rect 4960 59814 4990 59866
rect 4990 59814 5002 59866
rect 5002 59814 5016 59866
rect 5040 59814 5054 59866
rect 5054 59814 5066 59866
rect 5066 59814 5096 59866
rect 5120 59814 5130 59866
rect 5130 59814 5176 59866
rect 4880 59812 4936 59814
rect 4960 59812 5016 59814
rect 5040 59812 5096 59814
rect 5120 59812 5176 59814
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4880 58778 4936 58780
rect 4960 58778 5016 58780
rect 5040 58778 5096 58780
rect 5120 58778 5176 58780
rect 4880 58726 4926 58778
rect 4926 58726 4936 58778
rect 4960 58726 4990 58778
rect 4990 58726 5002 58778
rect 5002 58726 5016 58778
rect 5040 58726 5054 58778
rect 5054 58726 5066 58778
rect 5066 58726 5096 58778
rect 5120 58726 5130 58778
rect 5130 58726 5176 58778
rect 4880 58724 4936 58726
rect 4960 58724 5016 58726
rect 5040 58724 5096 58726
rect 5120 58724 5176 58726
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4880 57690 4936 57692
rect 4960 57690 5016 57692
rect 5040 57690 5096 57692
rect 5120 57690 5176 57692
rect 4880 57638 4926 57690
rect 4926 57638 4936 57690
rect 4960 57638 4990 57690
rect 4990 57638 5002 57690
rect 5002 57638 5016 57690
rect 5040 57638 5054 57690
rect 5054 57638 5066 57690
rect 5066 57638 5096 57690
rect 5120 57638 5130 57690
rect 5130 57638 5176 57690
rect 4880 57636 4936 57638
rect 4960 57636 5016 57638
rect 5040 57636 5096 57638
rect 5120 57636 5176 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4880 56602 4936 56604
rect 4960 56602 5016 56604
rect 5040 56602 5096 56604
rect 5120 56602 5176 56604
rect 4880 56550 4926 56602
rect 4926 56550 4936 56602
rect 4960 56550 4990 56602
rect 4990 56550 5002 56602
rect 5002 56550 5016 56602
rect 5040 56550 5054 56602
rect 5054 56550 5066 56602
rect 5066 56550 5096 56602
rect 5120 56550 5130 56602
rect 5130 56550 5176 56602
rect 4880 56548 4936 56550
rect 4960 56548 5016 56550
rect 5040 56548 5096 56550
rect 5120 56548 5176 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4880 55514 4936 55516
rect 4960 55514 5016 55516
rect 5040 55514 5096 55516
rect 5120 55514 5176 55516
rect 4880 55462 4926 55514
rect 4926 55462 4936 55514
rect 4960 55462 4990 55514
rect 4990 55462 5002 55514
rect 5002 55462 5016 55514
rect 5040 55462 5054 55514
rect 5054 55462 5066 55514
rect 5066 55462 5096 55514
rect 5120 55462 5130 55514
rect 5130 55462 5176 55514
rect 4880 55460 4936 55462
rect 4960 55460 5016 55462
rect 5040 55460 5096 55462
rect 5120 55460 5176 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4880 54426 4936 54428
rect 4960 54426 5016 54428
rect 5040 54426 5096 54428
rect 5120 54426 5176 54428
rect 4880 54374 4926 54426
rect 4926 54374 4936 54426
rect 4960 54374 4990 54426
rect 4990 54374 5002 54426
rect 5002 54374 5016 54426
rect 5040 54374 5054 54426
rect 5054 54374 5066 54426
rect 5066 54374 5096 54426
rect 5120 54374 5130 54426
rect 5130 54374 5176 54426
rect 4880 54372 4936 54374
rect 4960 54372 5016 54374
rect 5040 54372 5096 54374
rect 5120 54372 5176 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4880 53338 4936 53340
rect 4960 53338 5016 53340
rect 5040 53338 5096 53340
rect 5120 53338 5176 53340
rect 4880 53286 4926 53338
rect 4926 53286 4936 53338
rect 4960 53286 4990 53338
rect 4990 53286 5002 53338
rect 5002 53286 5016 53338
rect 5040 53286 5054 53338
rect 5054 53286 5066 53338
rect 5066 53286 5096 53338
rect 5120 53286 5130 53338
rect 5130 53286 5176 53338
rect 4880 53284 4936 53286
rect 4960 53284 5016 53286
rect 5040 53284 5096 53286
rect 5120 53284 5176 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4880 52250 4936 52252
rect 4960 52250 5016 52252
rect 5040 52250 5096 52252
rect 5120 52250 5176 52252
rect 4880 52198 4926 52250
rect 4926 52198 4936 52250
rect 4960 52198 4990 52250
rect 4990 52198 5002 52250
rect 5002 52198 5016 52250
rect 5040 52198 5054 52250
rect 5054 52198 5066 52250
rect 5066 52198 5096 52250
rect 5120 52198 5130 52250
rect 5130 52198 5176 52250
rect 4880 52196 4936 52198
rect 4960 52196 5016 52198
rect 5040 52196 5096 52198
rect 5120 52196 5176 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4880 51162 4936 51164
rect 4960 51162 5016 51164
rect 5040 51162 5096 51164
rect 5120 51162 5176 51164
rect 4880 51110 4926 51162
rect 4926 51110 4936 51162
rect 4960 51110 4990 51162
rect 4990 51110 5002 51162
rect 5002 51110 5016 51162
rect 5040 51110 5054 51162
rect 5054 51110 5066 51162
rect 5066 51110 5096 51162
rect 5120 51110 5130 51162
rect 5130 51110 5176 51162
rect 4880 51108 4936 51110
rect 4960 51108 5016 51110
rect 5040 51108 5096 51110
rect 5120 51108 5176 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4880 50074 4936 50076
rect 4960 50074 5016 50076
rect 5040 50074 5096 50076
rect 5120 50074 5176 50076
rect 4880 50022 4926 50074
rect 4926 50022 4936 50074
rect 4960 50022 4990 50074
rect 4990 50022 5002 50074
rect 5002 50022 5016 50074
rect 5040 50022 5054 50074
rect 5054 50022 5066 50074
rect 5066 50022 5096 50074
rect 5120 50022 5130 50074
rect 5130 50022 5176 50074
rect 4880 50020 4936 50022
rect 4960 50020 5016 50022
rect 5040 50020 5096 50022
rect 5120 50020 5176 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4880 48986 4936 48988
rect 4960 48986 5016 48988
rect 5040 48986 5096 48988
rect 5120 48986 5176 48988
rect 4880 48934 4926 48986
rect 4926 48934 4936 48986
rect 4960 48934 4990 48986
rect 4990 48934 5002 48986
rect 5002 48934 5016 48986
rect 5040 48934 5054 48986
rect 5054 48934 5066 48986
rect 5066 48934 5096 48986
rect 5120 48934 5130 48986
rect 5130 48934 5176 48986
rect 4880 48932 4936 48934
rect 4960 48932 5016 48934
rect 5040 48932 5096 48934
rect 5120 48932 5176 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4880 47898 4936 47900
rect 4960 47898 5016 47900
rect 5040 47898 5096 47900
rect 5120 47898 5176 47900
rect 4880 47846 4926 47898
rect 4926 47846 4936 47898
rect 4960 47846 4990 47898
rect 4990 47846 5002 47898
rect 5002 47846 5016 47898
rect 5040 47846 5054 47898
rect 5054 47846 5066 47898
rect 5066 47846 5096 47898
rect 5120 47846 5130 47898
rect 5130 47846 5176 47898
rect 4880 47844 4936 47846
rect 4960 47844 5016 47846
rect 5040 47844 5096 47846
rect 5120 47844 5176 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 1214 41556 1216 41576
rect 1216 41556 1268 41576
rect 1268 41556 1270 41576
rect 1214 41520 1270 41556
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 5538 41248 5594 41304
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 5538 39616 5594 39672
rect 1398 39480 1454 39536
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 8390 38428 8392 38448
rect 8392 38428 8444 38448
rect 8444 38428 8446 38448
rect 8390 38392 8446 38428
rect 1214 38120 1270 38176
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 1398 36760 1454 36816
rect 9494 36668 9550 36724
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 9494 35585 9550 35641
rect 1306 35400 1362 35456
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 1398 34040 1454 34096
rect 5538 33904 5594 33960
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1306 15680 1362 15736
rect 9494 15425 9550 15481
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 16394 67652 16450 67688
rect 16394 67632 16396 67652
rect 16396 67632 16448 67652
rect 16448 67632 16450 67652
rect 19338 66952 19394 67008
rect 20350 66816 20406 66872
rect 28998 66952 29054 67008
rect 27066 66816 27122 66872
rect 29734 66836 29790 66872
rect 29734 66816 29736 66836
rect 29736 66816 29788 66836
rect 29788 66816 29790 66836
rect 33046 66580 33048 66600
rect 33048 66580 33100 66600
rect 33100 66580 33102 66600
rect 33046 66544 33102 66580
rect 35600 67482 35656 67484
rect 35680 67482 35736 67484
rect 35760 67482 35816 67484
rect 35840 67482 35896 67484
rect 35600 67430 35646 67482
rect 35646 67430 35656 67482
rect 35680 67430 35710 67482
rect 35710 67430 35722 67482
rect 35722 67430 35736 67482
rect 35760 67430 35774 67482
rect 35774 67430 35786 67482
rect 35786 67430 35816 67482
rect 35840 67430 35850 67482
rect 35850 67430 35896 67482
rect 35600 67428 35656 67430
rect 35680 67428 35736 67430
rect 35760 67428 35816 67430
rect 35840 67428 35896 67430
rect 40958 69844 40960 69864
rect 40960 69844 41012 69864
rect 41012 69844 41014 69864
rect 40958 69808 41014 69844
rect 43258 69808 43314 69864
rect 42154 69536 42210 69592
rect 65660 68026 65716 68028
rect 65740 68026 65796 68028
rect 65820 68026 65876 68028
rect 65900 68026 65956 68028
rect 65660 67974 65706 68026
rect 65706 67974 65716 68026
rect 65740 67974 65770 68026
rect 65770 67974 65782 68026
rect 65782 67974 65796 68026
rect 65820 67974 65834 68026
rect 65834 67974 65846 68026
rect 65846 67974 65876 68026
rect 65900 67974 65910 68026
rect 65910 67974 65956 68026
rect 65660 67972 65716 67974
rect 65740 67972 65796 67974
rect 65820 67972 65876 67974
rect 65900 67972 65956 67974
rect 40406 67496 40462 67552
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 33874 66544 33930 66600
rect 35346 66544 35402 66600
rect 35600 66394 35656 66396
rect 35680 66394 35736 66396
rect 35760 66394 35816 66396
rect 35840 66394 35896 66396
rect 35600 66342 35646 66394
rect 35646 66342 35656 66394
rect 35680 66342 35710 66394
rect 35710 66342 35722 66394
rect 35722 66342 35736 66394
rect 35760 66342 35774 66394
rect 35774 66342 35786 66394
rect 35786 66342 35816 66394
rect 35840 66342 35850 66394
rect 35850 66342 35896 66394
rect 35600 66340 35656 66342
rect 35680 66340 35736 66342
rect 35760 66340 35816 66342
rect 35840 66340 35896 66342
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 33506 65456 33562 65512
rect 39118 66680 39174 66736
rect 39026 66272 39082 66328
rect 66320 67482 66376 67484
rect 66400 67482 66456 67484
rect 66480 67482 66536 67484
rect 66560 67482 66616 67484
rect 66320 67430 66366 67482
rect 66366 67430 66376 67482
rect 66400 67430 66430 67482
rect 66430 67430 66442 67482
rect 66442 67430 66456 67482
rect 66480 67430 66494 67482
rect 66494 67430 66506 67482
rect 66506 67430 66536 67482
rect 66560 67430 66570 67482
rect 66570 67430 66616 67482
rect 66320 67428 66376 67430
rect 66400 67428 66456 67430
rect 66480 67428 66536 67430
rect 66560 67428 66616 67430
rect 46662 67260 46664 67280
rect 46664 67260 46716 67280
rect 46716 67260 46718 67280
rect 44454 67124 44456 67144
rect 44456 67124 44508 67144
rect 44508 67124 44510 67144
rect 44454 67088 44510 67124
rect 46662 67224 46718 67260
rect 45742 66136 45798 66192
rect 62394 67244 62450 67280
rect 62394 67224 62396 67244
rect 62396 67224 62448 67244
rect 62448 67224 62450 67244
rect 69018 67496 69074 67552
rect 62210 67108 62266 67144
rect 62210 67088 62212 67108
rect 62212 67088 62264 67108
rect 62264 67088 62266 67108
rect 47858 66544 47914 66600
rect 53654 65900 53656 65920
rect 53656 65900 53708 65920
rect 53708 65900 53710 65920
rect 53654 65864 53710 65900
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 35990 64096 36046 64152
rect 47490 64096 47546 64152
rect 63406 64096 63462 64152
rect 67546 66680 67602 66736
rect 67638 66564 67694 66600
rect 67638 66544 67640 66564
rect 67640 66544 67692 66564
rect 67692 66544 67694 66564
rect 69754 68176 69810 68232
rect 70398 66952 70454 67008
rect 90362 69808 90418 69864
rect 79966 67496 80022 67552
rect 75366 67380 75422 67416
rect 75366 67360 75368 67380
rect 75368 67360 75420 67380
rect 75420 67360 75422 67380
rect 66320 66394 66376 66396
rect 66400 66394 66456 66396
rect 66480 66394 66536 66396
rect 66560 66394 66616 66396
rect 66320 66342 66366 66394
rect 66366 66342 66376 66394
rect 66400 66342 66430 66394
rect 66430 66342 66442 66394
rect 66442 66342 66456 66394
rect 66480 66342 66494 66394
rect 66494 66342 66506 66394
rect 66506 66342 66536 66394
rect 66560 66342 66570 66394
rect 66570 66342 66616 66394
rect 66320 66340 66376 66342
rect 66400 66340 66456 66342
rect 66480 66340 66536 66342
rect 66560 66340 66616 66342
rect 66166 63960 66222 64016
rect 73710 66272 73766 66328
rect 84842 66700 84898 66736
rect 84842 66680 84844 66700
rect 84844 66680 84896 66700
rect 84896 66680 84898 66700
rect 84658 66580 84660 66600
rect 84660 66580 84712 66600
rect 84712 66580 84714 66600
rect 84658 66544 84714 66580
rect 85578 66952 85634 67008
rect 96894 69536 96950 69592
rect 90822 68720 90878 68776
rect 85394 66700 85450 66736
rect 85394 66680 85396 66700
rect 85396 66680 85448 66700
rect 85448 66680 85450 66700
rect 84934 65456 84990 65512
rect 87970 66444 87972 66464
rect 87972 66444 88024 66464
rect 88024 66444 88026 66464
rect 87970 66408 88026 66444
rect 88522 66408 88578 66464
rect 90914 67632 90970 67688
rect 90822 67532 90824 67552
rect 90824 67532 90876 67552
rect 90876 67532 90878 67552
rect 90822 67496 90878 67532
rect 91006 66272 91062 66328
rect 94778 67496 94834 67552
rect 95606 67768 95662 67824
rect 95330 67668 95332 67688
rect 95332 67668 95384 67688
rect 95384 67668 95386 67688
rect 95330 67632 95386 67668
rect 95790 67532 95792 67552
rect 95792 67532 95844 67552
rect 95844 67532 95846 67552
rect 95790 67496 95846 67532
rect 96380 68026 96436 68028
rect 96460 68026 96516 68028
rect 96540 68026 96596 68028
rect 96620 68026 96676 68028
rect 96380 67974 96426 68026
rect 96426 67974 96436 68026
rect 96460 67974 96490 68026
rect 96490 67974 96502 68026
rect 96502 67974 96516 68026
rect 96540 67974 96554 68026
rect 96554 67974 96566 68026
rect 96566 67974 96596 68026
rect 96620 67974 96630 68026
rect 96630 67974 96676 68026
rect 96380 67972 96436 67974
rect 96460 67972 96516 67974
rect 96540 67972 96596 67974
rect 96620 67972 96676 67974
rect 96618 67668 96620 67688
rect 96620 67668 96672 67688
rect 96672 67668 96674 67688
rect 96618 67632 96674 67668
rect 96710 67496 96766 67552
rect 96380 66938 96436 66940
rect 96460 66938 96516 66940
rect 96540 66938 96596 66940
rect 96620 66938 96676 66940
rect 96380 66886 96426 66938
rect 96426 66886 96436 66938
rect 96460 66886 96490 66938
rect 96490 66886 96502 66938
rect 96502 66886 96516 66938
rect 96540 66886 96554 66938
rect 96554 66886 96566 66938
rect 96566 66886 96596 66938
rect 96620 66886 96630 66938
rect 96630 66886 96676 66938
rect 96380 66884 96436 66886
rect 96460 66884 96516 66886
rect 96540 66884 96596 66886
rect 96620 66884 96676 66886
rect 75458 64096 75514 64152
rect 96380 65850 96436 65852
rect 96460 65850 96516 65852
rect 96540 65850 96596 65852
rect 96620 65850 96676 65852
rect 96380 65798 96426 65850
rect 96426 65798 96436 65850
rect 96460 65798 96490 65850
rect 96490 65798 96502 65850
rect 96502 65798 96516 65850
rect 96540 65798 96554 65850
rect 96554 65798 96566 65850
rect 96566 65798 96596 65850
rect 96620 65798 96630 65850
rect 96630 65798 96676 65850
rect 96380 65796 96436 65798
rect 96460 65796 96516 65798
rect 96540 65796 96596 65798
rect 96620 65796 96676 65798
rect 96986 67788 97042 67824
rect 96986 67768 96988 67788
rect 96988 67768 97040 67788
rect 97040 67768 97042 67788
rect 97040 67482 97096 67484
rect 97120 67482 97176 67484
rect 97200 67482 97256 67484
rect 97280 67482 97336 67484
rect 97040 67430 97086 67482
rect 97086 67430 97096 67482
rect 97120 67430 97150 67482
rect 97150 67430 97162 67482
rect 97162 67430 97176 67482
rect 97200 67430 97214 67482
rect 97214 67430 97226 67482
rect 97226 67430 97256 67482
rect 97280 67430 97290 67482
rect 97290 67430 97336 67482
rect 97040 67428 97096 67430
rect 97120 67428 97176 67430
rect 97200 67428 97256 67430
rect 97280 67428 97336 67430
rect 102046 83332 102102 83388
rect 105928 126778 105984 126780
rect 106008 126778 106064 126780
rect 106088 126778 106144 126780
rect 106168 126778 106224 126780
rect 105928 126726 105974 126778
rect 105974 126726 105984 126778
rect 106008 126726 106038 126778
rect 106038 126726 106050 126778
rect 106050 126726 106064 126778
rect 106088 126726 106102 126778
rect 106102 126726 106114 126778
rect 106114 126726 106144 126778
rect 106168 126726 106178 126778
rect 106178 126726 106224 126778
rect 105928 126724 105984 126726
rect 106008 126724 106064 126726
rect 106088 126724 106144 126726
rect 106168 126724 106224 126726
rect 102230 67496 102286 67552
rect 97040 66394 97096 66396
rect 97120 66394 97176 66396
rect 97200 66394 97256 66396
rect 97280 66394 97336 66396
rect 97040 66342 97086 66394
rect 97086 66342 97096 66394
rect 97120 66342 97150 66394
rect 97150 66342 97162 66394
rect 97162 66342 97176 66394
rect 97200 66342 97214 66394
rect 97214 66342 97226 66394
rect 97226 66342 97256 66394
rect 97280 66342 97290 66394
rect 97290 66342 97336 66394
rect 97040 66340 97096 66342
rect 97120 66340 97176 66342
rect 97200 66340 97256 66342
rect 97280 66340 97336 66342
rect 102138 67224 102194 67280
rect 106664 126234 106720 126236
rect 106744 126234 106800 126236
rect 106824 126234 106880 126236
rect 106904 126234 106960 126236
rect 106664 126182 106710 126234
rect 106710 126182 106720 126234
rect 106744 126182 106774 126234
rect 106774 126182 106786 126234
rect 106786 126182 106800 126234
rect 106824 126182 106838 126234
rect 106838 126182 106850 126234
rect 106850 126182 106880 126234
rect 106904 126182 106914 126234
rect 106914 126182 106960 126234
rect 106664 126180 106720 126182
rect 106744 126180 106800 126182
rect 106824 126180 106880 126182
rect 106904 126180 106960 126182
rect 102782 123800 102838 123856
rect 103058 82184 103114 82240
rect 102414 68176 102470 68232
rect 105928 125690 105984 125692
rect 106008 125690 106064 125692
rect 106088 125690 106144 125692
rect 106168 125690 106224 125692
rect 105928 125638 105974 125690
rect 105974 125638 105984 125690
rect 106008 125638 106038 125690
rect 106038 125638 106050 125690
rect 106050 125638 106064 125690
rect 106088 125638 106102 125690
rect 106102 125638 106114 125690
rect 106114 125638 106144 125690
rect 106168 125638 106178 125690
rect 106178 125638 106224 125690
rect 105928 125636 105984 125638
rect 106008 125636 106064 125638
rect 106088 125636 106144 125638
rect 106168 125636 106224 125638
rect 106664 125146 106720 125148
rect 106744 125146 106800 125148
rect 106824 125146 106880 125148
rect 106904 125146 106960 125148
rect 106664 125094 106710 125146
rect 106710 125094 106720 125146
rect 106744 125094 106774 125146
rect 106774 125094 106786 125146
rect 106786 125094 106800 125146
rect 106824 125094 106838 125146
rect 106838 125094 106850 125146
rect 106850 125094 106880 125146
rect 106904 125094 106914 125146
rect 106914 125094 106960 125146
rect 106664 125092 106720 125094
rect 106744 125092 106800 125094
rect 106824 125092 106880 125094
rect 106904 125092 106960 125094
rect 105928 124602 105984 124604
rect 106008 124602 106064 124604
rect 106088 124602 106144 124604
rect 106168 124602 106224 124604
rect 105928 124550 105974 124602
rect 105974 124550 105984 124602
rect 106008 124550 106038 124602
rect 106038 124550 106050 124602
rect 106050 124550 106064 124602
rect 106088 124550 106102 124602
rect 106102 124550 106114 124602
rect 106114 124550 106144 124602
rect 106168 124550 106178 124602
rect 106178 124550 106224 124602
rect 105928 124548 105984 124550
rect 106008 124548 106064 124550
rect 106088 124548 106144 124550
rect 106168 124548 106224 124550
rect 106664 124058 106720 124060
rect 106744 124058 106800 124060
rect 106824 124058 106880 124060
rect 106904 124058 106960 124060
rect 106664 124006 106710 124058
rect 106710 124006 106720 124058
rect 106744 124006 106774 124058
rect 106774 124006 106786 124058
rect 106786 124006 106800 124058
rect 106824 124006 106838 124058
rect 106838 124006 106850 124058
rect 106850 124006 106880 124058
rect 106904 124006 106914 124058
rect 106914 124006 106960 124058
rect 106664 124004 106720 124006
rect 106744 124004 106800 124006
rect 106824 124004 106880 124006
rect 106904 124004 106960 124006
rect 104714 123936 104770 123992
rect 104346 119720 104402 119776
rect 105928 123514 105984 123516
rect 106008 123514 106064 123516
rect 106088 123514 106144 123516
rect 106168 123514 106224 123516
rect 105928 123462 105974 123514
rect 105974 123462 105984 123514
rect 106008 123462 106038 123514
rect 106038 123462 106050 123514
rect 106050 123462 106064 123514
rect 106088 123462 106102 123514
rect 106102 123462 106114 123514
rect 106114 123462 106144 123514
rect 106168 123462 106178 123514
rect 106178 123462 106224 123514
rect 105928 123460 105984 123462
rect 106008 123460 106064 123462
rect 106088 123460 106144 123462
rect 106168 123460 106224 123462
rect 106664 122970 106720 122972
rect 106744 122970 106800 122972
rect 106824 122970 106880 122972
rect 106904 122970 106960 122972
rect 106664 122918 106710 122970
rect 106710 122918 106720 122970
rect 106744 122918 106774 122970
rect 106774 122918 106786 122970
rect 106786 122918 106800 122970
rect 106824 122918 106838 122970
rect 106838 122918 106850 122970
rect 106850 122918 106880 122970
rect 106904 122918 106914 122970
rect 106914 122918 106960 122970
rect 106664 122916 106720 122918
rect 106744 122916 106800 122918
rect 106824 122916 106880 122918
rect 106904 122916 106960 122918
rect 105928 122426 105984 122428
rect 106008 122426 106064 122428
rect 106088 122426 106144 122428
rect 106168 122426 106224 122428
rect 105928 122374 105974 122426
rect 105974 122374 105984 122426
rect 106008 122374 106038 122426
rect 106038 122374 106050 122426
rect 106050 122374 106064 122426
rect 106088 122374 106102 122426
rect 106102 122374 106114 122426
rect 106114 122374 106144 122426
rect 106168 122374 106178 122426
rect 106178 122374 106224 122426
rect 105928 122372 105984 122374
rect 106008 122372 106064 122374
rect 106088 122372 106144 122374
rect 106168 122372 106224 122374
rect 106664 121882 106720 121884
rect 106744 121882 106800 121884
rect 106824 121882 106880 121884
rect 106904 121882 106960 121884
rect 106664 121830 106710 121882
rect 106710 121830 106720 121882
rect 106744 121830 106774 121882
rect 106774 121830 106786 121882
rect 106786 121830 106800 121882
rect 106824 121830 106838 121882
rect 106838 121830 106850 121882
rect 106850 121830 106880 121882
rect 106904 121830 106914 121882
rect 106914 121830 106960 121882
rect 106664 121828 106720 121830
rect 106744 121828 106800 121830
rect 106824 121828 106880 121830
rect 106904 121828 106960 121830
rect 105928 121338 105984 121340
rect 106008 121338 106064 121340
rect 106088 121338 106144 121340
rect 106168 121338 106224 121340
rect 105928 121286 105974 121338
rect 105974 121286 105984 121338
rect 106008 121286 106038 121338
rect 106038 121286 106050 121338
rect 106050 121286 106064 121338
rect 106088 121286 106102 121338
rect 106102 121286 106114 121338
rect 106114 121286 106144 121338
rect 106168 121286 106178 121338
rect 106178 121286 106224 121338
rect 105928 121284 105984 121286
rect 106008 121284 106064 121286
rect 106088 121284 106144 121286
rect 106168 121284 106224 121286
rect 106664 120794 106720 120796
rect 106744 120794 106800 120796
rect 106824 120794 106880 120796
rect 106904 120794 106960 120796
rect 106664 120742 106710 120794
rect 106710 120742 106720 120794
rect 106744 120742 106774 120794
rect 106774 120742 106786 120794
rect 106786 120742 106800 120794
rect 106824 120742 106838 120794
rect 106838 120742 106850 120794
rect 106850 120742 106880 120794
rect 106904 120742 106914 120794
rect 106914 120742 106960 120794
rect 106664 120740 106720 120742
rect 106744 120740 106800 120742
rect 106824 120740 106880 120742
rect 106904 120740 106960 120742
rect 105928 120250 105984 120252
rect 106008 120250 106064 120252
rect 106088 120250 106144 120252
rect 106168 120250 106224 120252
rect 105928 120198 105974 120250
rect 105974 120198 105984 120250
rect 106008 120198 106038 120250
rect 106038 120198 106050 120250
rect 106050 120198 106064 120250
rect 106088 120198 106102 120250
rect 106102 120198 106114 120250
rect 106114 120198 106144 120250
rect 106168 120198 106178 120250
rect 106178 120198 106224 120250
rect 105928 120196 105984 120198
rect 106008 120196 106064 120198
rect 106088 120196 106144 120198
rect 106168 120196 106224 120198
rect 106664 119706 106720 119708
rect 106744 119706 106800 119708
rect 106824 119706 106880 119708
rect 106904 119706 106960 119708
rect 106664 119654 106710 119706
rect 106710 119654 106720 119706
rect 106744 119654 106774 119706
rect 106774 119654 106786 119706
rect 106786 119654 106800 119706
rect 106824 119654 106838 119706
rect 106838 119654 106850 119706
rect 106850 119654 106880 119706
rect 106904 119654 106914 119706
rect 106914 119654 106960 119706
rect 106664 119652 106720 119654
rect 106744 119652 106800 119654
rect 106824 119652 106880 119654
rect 106904 119652 106960 119654
rect 105928 119162 105984 119164
rect 106008 119162 106064 119164
rect 106088 119162 106144 119164
rect 106168 119162 106224 119164
rect 105928 119110 105974 119162
rect 105974 119110 105984 119162
rect 106008 119110 106038 119162
rect 106038 119110 106050 119162
rect 106050 119110 106064 119162
rect 106088 119110 106102 119162
rect 106102 119110 106114 119162
rect 106114 119110 106144 119162
rect 106168 119110 106178 119162
rect 106178 119110 106224 119162
rect 105928 119108 105984 119110
rect 106008 119108 106064 119110
rect 106088 119108 106144 119110
rect 106168 119108 106224 119110
rect 106664 118618 106720 118620
rect 106744 118618 106800 118620
rect 106824 118618 106880 118620
rect 106904 118618 106960 118620
rect 106664 118566 106710 118618
rect 106710 118566 106720 118618
rect 106744 118566 106774 118618
rect 106774 118566 106786 118618
rect 106786 118566 106800 118618
rect 106824 118566 106838 118618
rect 106838 118566 106850 118618
rect 106850 118566 106880 118618
rect 106904 118566 106914 118618
rect 106914 118566 106960 118618
rect 106664 118564 106720 118566
rect 106744 118564 106800 118566
rect 106824 118564 106880 118566
rect 106904 118564 106960 118566
rect 105928 118074 105984 118076
rect 106008 118074 106064 118076
rect 106088 118074 106144 118076
rect 106168 118074 106224 118076
rect 105928 118022 105974 118074
rect 105974 118022 105984 118074
rect 106008 118022 106038 118074
rect 106038 118022 106050 118074
rect 106050 118022 106064 118074
rect 106088 118022 106102 118074
rect 106102 118022 106114 118074
rect 106114 118022 106144 118074
rect 106168 118022 106178 118074
rect 106178 118022 106224 118074
rect 105928 118020 105984 118022
rect 106008 118020 106064 118022
rect 106088 118020 106144 118022
rect 106168 118020 106224 118022
rect 106664 117530 106720 117532
rect 106744 117530 106800 117532
rect 106824 117530 106880 117532
rect 106904 117530 106960 117532
rect 106664 117478 106710 117530
rect 106710 117478 106720 117530
rect 106744 117478 106774 117530
rect 106774 117478 106786 117530
rect 106786 117478 106800 117530
rect 106824 117478 106838 117530
rect 106838 117478 106850 117530
rect 106850 117478 106880 117530
rect 106904 117478 106914 117530
rect 106914 117478 106960 117530
rect 106664 117476 106720 117478
rect 106744 117476 106800 117478
rect 106824 117476 106880 117478
rect 106904 117476 106960 117478
rect 105928 116986 105984 116988
rect 106008 116986 106064 116988
rect 106088 116986 106144 116988
rect 106168 116986 106224 116988
rect 105928 116934 105974 116986
rect 105974 116934 105984 116986
rect 106008 116934 106038 116986
rect 106038 116934 106050 116986
rect 106050 116934 106064 116986
rect 106088 116934 106102 116986
rect 106102 116934 106114 116986
rect 106114 116934 106144 116986
rect 106168 116934 106178 116986
rect 106178 116934 106224 116986
rect 105928 116932 105984 116934
rect 106008 116932 106064 116934
rect 106088 116932 106144 116934
rect 106168 116932 106224 116934
rect 106664 116442 106720 116444
rect 106744 116442 106800 116444
rect 106824 116442 106880 116444
rect 106904 116442 106960 116444
rect 106664 116390 106710 116442
rect 106710 116390 106720 116442
rect 106744 116390 106774 116442
rect 106774 116390 106786 116442
rect 106786 116390 106800 116442
rect 106824 116390 106838 116442
rect 106838 116390 106850 116442
rect 106850 116390 106880 116442
rect 106904 116390 106914 116442
rect 106914 116390 106960 116442
rect 106664 116388 106720 116390
rect 106744 116388 106800 116390
rect 106824 116388 106880 116390
rect 106904 116388 106960 116390
rect 105928 115898 105984 115900
rect 106008 115898 106064 115900
rect 106088 115898 106144 115900
rect 106168 115898 106224 115900
rect 105928 115846 105974 115898
rect 105974 115846 105984 115898
rect 106008 115846 106038 115898
rect 106038 115846 106050 115898
rect 106050 115846 106064 115898
rect 106088 115846 106102 115898
rect 106102 115846 106114 115898
rect 106114 115846 106144 115898
rect 106168 115846 106178 115898
rect 106178 115846 106224 115898
rect 105928 115844 105984 115846
rect 106008 115844 106064 115846
rect 106088 115844 106144 115846
rect 106168 115844 106224 115846
rect 106664 115354 106720 115356
rect 106744 115354 106800 115356
rect 106824 115354 106880 115356
rect 106904 115354 106960 115356
rect 106664 115302 106710 115354
rect 106710 115302 106720 115354
rect 106744 115302 106774 115354
rect 106774 115302 106786 115354
rect 106786 115302 106800 115354
rect 106824 115302 106838 115354
rect 106838 115302 106850 115354
rect 106850 115302 106880 115354
rect 106904 115302 106914 115354
rect 106914 115302 106960 115354
rect 106664 115300 106720 115302
rect 106744 115300 106800 115302
rect 106824 115300 106880 115302
rect 106904 115300 106960 115302
rect 105928 114810 105984 114812
rect 106008 114810 106064 114812
rect 106088 114810 106144 114812
rect 106168 114810 106224 114812
rect 105928 114758 105974 114810
rect 105974 114758 105984 114810
rect 106008 114758 106038 114810
rect 106038 114758 106050 114810
rect 106050 114758 106064 114810
rect 106088 114758 106102 114810
rect 106102 114758 106114 114810
rect 106114 114758 106144 114810
rect 106168 114758 106178 114810
rect 106178 114758 106224 114810
rect 105928 114756 105984 114758
rect 106008 114756 106064 114758
rect 106088 114756 106144 114758
rect 106168 114756 106224 114758
rect 106664 114266 106720 114268
rect 106744 114266 106800 114268
rect 106824 114266 106880 114268
rect 106904 114266 106960 114268
rect 106664 114214 106710 114266
rect 106710 114214 106720 114266
rect 106744 114214 106774 114266
rect 106774 114214 106786 114266
rect 106786 114214 106800 114266
rect 106824 114214 106838 114266
rect 106838 114214 106850 114266
rect 106850 114214 106880 114266
rect 106904 114214 106914 114266
rect 106914 114214 106960 114266
rect 106664 114212 106720 114214
rect 106744 114212 106800 114214
rect 106824 114212 106880 114214
rect 106904 114212 106960 114214
rect 105928 113722 105984 113724
rect 106008 113722 106064 113724
rect 106088 113722 106144 113724
rect 106168 113722 106224 113724
rect 105928 113670 105974 113722
rect 105974 113670 105984 113722
rect 106008 113670 106038 113722
rect 106038 113670 106050 113722
rect 106050 113670 106064 113722
rect 106088 113670 106102 113722
rect 106102 113670 106114 113722
rect 106114 113670 106144 113722
rect 106168 113670 106178 113722
rect 106178 113670 106224 113722
rect 105928 113668 105984 113670
rect 106008 113668 106064 113670
rect 106088 113668 106144 113670
rect 106168 113668 106224 113670
rect 106664 113178 106720 113180
rect 106744 113178 106800 113180
rect 106824 113178 106880 113180
rect 106904 113178 106960 113180
rect 106664 113126 106710 113178
rect 106710 113126 106720 113178
rect 106744 113126 106774 113178
rect 106774 113126 106786 113178
rect 106786 113126 106800 113178
rect 106824 113126 106838 113178
rect 106838 113126 106850 113178
rect 106850 113126 106880 113178
rect 106904 113126 106914 113178
rect 106914 113126 106960 113178
rect 106664 113124 106720 113126
rect 106744 113124 106800 113126
rect 106824 113124 106880 113126
rect 106904 113124 106960 113126
rect 105928 112634 105984 112636
rect 106008 112634 106064 112636
rect 106088 112634 106144 112636
rect 106168 112634 106224 112636
rect 105928 112582 105974 112634
rect 105974 112582 105984 112634
rect 106008 112582 106038 112634
rect 106038 112582 106050 112634
rect 106050 112582 106064 112634
rect 106088 112582 106102 112634
rect 106102 112582 106114 112634
rect 106114 112582 106144 112634
rect 106168 112582 106178 112634
rect 106178 112582 106224 112634
rect 105928 112580 105984 112582
rect 106008 112580 106064 112582
rect 106088 112580 106144 112582
rect 106168 112580 106224 112582
rect 106664 112090 106720 112092
rect 106744 112090 106800 112092
rect 106824 112090 106880 112092
rect 106904 112090 106960 112092
rect 106664 112038 106710 112090
rect 106710 112038 106720 112090
rect 106744 112038 106774 112090
rect 106774 112038 106786 112090
rect 106786 112038 106800 112090
rect 106824 112038 106838 112090
rect 106838 112038 106850 112090
rect 106850 112038 106880 112090
rect 106904 112038 106914 112090
rect 106914 112038 106960 112090
rect 106664 112036 106720 112038
rect 106744 112036 106800 112038
rect 106824 112036 106880 112038
rect 106904 112036 106960 112038
rect 105928 111546 105984 111548
rect 106008 111546 106064 111548
rect 106088 111546 106144 111548
rect 106168 111546 106224 111548
rect 105928 111494 105974 111546
rect 105974 111494 105984 111546
rect 106008 111494 106038 111546
rect 106038 111494 106050 111546
rect 106050 111494 106064 111546
rect 106088 111494 106102 111546
rect 106102 111494 106114 111546
rect 106114 111494 106144 111546
rect 106168 111494 106178 111546
rect 106178 111494 106224 111546
rect 105928 111492 105984 111494
rect 106008 111492 106064 111494
rect 106088 111492 106144 111494
rect 106168 111492 106224 111494
rect 106664 111002 106720 111004
rect 106744 111002 106800 111004
rect 106824 111002 106880 111004
rect 106904 111002 106960 111004
rect 106664 110950 106710 111002
rect 106710 110950 106720 111002
rect 106744 110950 106774 111002
rect 106774 110950 106786 111002
rect 106786 110950 106800 111002
rect 106824 110950 106838 111002
rect 106838 110950 106850 111002
rect 106850 110950 106880 111002
rect 106904 110950 106914 111002
rect 106914 110950 106960 111002
rect 106664 110948 106720 110950
rect 106744 110948 106800 110950
rect 106824 110948 106880 110950
rect 106904 110948 106960 110950
rect 105928 110458 105984 110460
rect 106008 110458 106064 110460
rect 106088 110458 106144 110460
rect 106168 110458 106224 110460
rect 105928 110406 105974 110458
rect 105974 110406 105984 110458
rect 106008 110406 106038 110458
rect 106038 110406 106050 110458
rect 106050 110406 106064 110458
rect 106088 110406 106102 110458
rect 106102 110406 106114 110458
rect 106114 110406 106144 110458
rect 106168 110406 106178 110458
rect 106178 110406 106224 110458
rect 105928 110404 105984 110406
rect 106008 110404 106064 110406
rect 106088 110404 106144 110406
rect 106168 110404 106224 110406
rect 106664 109914 106720 109916
rect 106744 109914 106800 109916
rect 106824 109914 106880 109916
rect 106904 109914 106960 109916
rect 106664 109862 106710 109914
rect 106710 109862 106720 109914
rect 106744 109862 106774 109914
rect 106774 109862 106786 109914
rect 106786 109862 106800 109914
rect 106824 109862 106838 109914
rect 106838 109862 106850 109914
rect 106850 109862 106880 109914
rect 106904 109862 106914 109914
rect 106914 109862 106960 109914
rect 106664 109860 106720 109862
rect 106744 109860 106800 109862
rect 106824 109860 106880 109862
rect 106904 109860 106960 109862
rect 105928 109370 105984 109372
rect 106008 109370 106064 109372
rect 106088 109370 106144 109372
rect 106168 109370 106224 109372
rect 105928 109318 105974 109370
rect 105974 109318 105984 109370
rect 106008 109318 106038 109370
rect 106038 109318 106050 109370
rect 106050 109318 106064 109370
rect 106088 109318 106102 109370
rect 106102 109318 106114 109370
rect 106114 109318 106144 109370
rect 106168 109318 106178 109370
rect 106178 109318 106224 109370
rect 105928 109316 105984 109318
rect 106008 109316 106064 109318
rect 106088 109316 106144 109318
rect 106168 109316 106224 109318
rect 106664 108826 106720 108828
rect 106744 108826 106800 108828
rect 106824 108826 106880 108828
rect 106904 108826 106960 108828
rect 106664 108774 106710 108826
rect 106710 108774 106720 108826
rect 106744 108774 106774 108826
rect 106774 108774 106786 108826
rect 106786 108774 106800 108826
rect 106824 108774 106838 108826
rect 106838 108774 106850 108826
rect 106850 108774 106880 108826
rect 106904 108774 106914 108826
rect 106914 108774 106960 108826
rect 106664 108772 106720 108774
rect 106744 108772 106800 108774
rect 106824 108772 106880 108774
rect 106904 108772 106960 108774
rect 105928 108282 105984 108284
rect 106008 108282 106064 108284
rect 106088 108282 106144 108284
rect 106168 108282 106224 108284
rect 105928 108230 105974 108282
rect 105974 108230 105984 108282
rect 106008 108230 106038 108282
rect 106038 108230 106050 108282
rect 106050 108230 106064 108282
rect 106088 108230 106102 108282
rect 106102 108230 106114 108282
rect 106114 108230 106144 108282
rect 106168 108230 106178 108282
rect 106178 108230 106224 108282
rect 105928 108228 105984 108230
rect 106008 108228 106064 108230
rect 106088 108228 106144 108230
rect 106168 108228 106224 108230
rect 106664 107738 106720 107740
rect 106744 107738 106800 107740
rect 106824 107738 106880 107740
rect 106904 107738 106960 107740
rect 106664 107686 106710 107738
rect 106710 107686 106720 107738
rect 106744 107686 106774 107738
rect 106774 107686 106786 107738
rect 106786 107686 106800 107738
rect 106824 107686 106838 107738
rect 106838 107686 106850 107738
rect 106850 107686 106880 107738
rect 106904 107686 106914 107738
rect 106914 107686 106960 107738
rect 106664 107684 106720 107686
rect 106744 107684 106800 107686
rect 106824 107684 106880 107686
rect 106904 107684 106960 107686
rect 105928 107194 105984 107196
rect 106008 107194 106064 107196
rect 106088 107194 106144 107196
rect 106168 107194 106224 107196
rect 105928 107142 105974 107194
rect 105974 107142 105984 107194
rect 106008 107142 106038 107194
rect 106038 107142 106050 107194
rect 106050 107142 106064 107194
rect 106088 107142 106102 107194
rect 106102 107142 106114 107194
rect 106114 107142 106144 107194
rect 106168 107142 106178 107194
rect 106178 107142 106224 107194
rect 105928 107140 105984 107142
rect 106008 107140 106064 107142
rect 106088 107140 106144 107142
rect 106168 107140 106224 107142
rect 106664 106650 106720 106652
rect 106744 106650 106800 106652
rect 106824 106650 106880 106652
rect 106904 106650 106960 106652
rect 106664 106598 106710 106650
rect 106710 106598 106720 106650
rect 106744 106598 106774 106650
rect 106774 106598 106786 106650
rect 106786 106598 106800 106650
rect 106824 106598 106838 106650
rect 106838 106598 106850 106650
rect 106850 106598 106880 106650
rect 106904 106598 106914 106650
rect 106914 106598 106960 106650
rect 106664 106596 106720 106598
rect 106744 106596 106800 106598
rect 106824 106596 106880 106598
rect 106904 106596 106960 106598
rect 105928 106106 105984 106108
rect 106008 106106 106064 106108
rect 106088 106106 106144 106108
rect 106168 106106 106224 106108
rect 105928 106054 105974 106106
rect 105974 106054 105984 106106
rect 106008 106054 106038 106106
rect 106038 106054 106050 106106
rect 106050 106054 106064 106106
rect 106088 106054 106102 106106
rect 106102 106054 106114 106106
rect 106114 106054 106144 106106
rect 106168 106054 106178 106106
rect 106178 106054 106224 106106
rect 105928 106052 105984 106054
rect 106008 106052 106064 106054
rect 106088 106052 106144 106054
rect 106168 106052 106224 106054
rect 106664 105562 106720 105564
rect 106744 105562 106800 105564
rect 106824 105562 106880 105564
rect 106904 105562 106960 105564
rect 106664 105510 106710 105562
rect 106710 105510 106720 105562
rect 106744 105510 106774 105562
rect 106774 105510 106786 105562
rect 106786 105510 106800 105562
rect 106824 105510 106838 105562
rect 106838 105510 106850 105562
rect 106850 105510 106880 105562
rect 106904 105510 106914 105562
rect 106914 105510 106960 105562
rect 106664 105508 106720 105510
rect 106744 105508 106800 105510
rect 106824 105508 106880 105510
rect 106904 105508 106960 105510
rect 105928 105018 105984 105020
rect 106008 105018 106064 105020
rect 106088 105018 106144 105020
rect 106168 105018 106224 105020
rect 105928 104966 105974 105018
rect 105974 104966 105984 105018
rect 106008 104966 106038 105018
rect 106038 104966 106050 105018
rect 106050 104966 106064 105018
rect 106088 104966 106102 105018
rect 106102 104966 106114 105018
rect 106114 104966 106144 105018
rect 106168 104966 106178 105018
rect 106178 104966 106224 105018
rect 105928 104964 105984 104966
rect 106008 104964 106064 104966
rect 106088 104964 106144 104966
rect 106168 104964 106224 104966
rect 106664 104474 106720 104476
rect 106744 104474 106800 104476
rect 106824 104474 106880 104476
rect 106904 104474 106960 104476
rect 106664 104422 106710 104474
rect 106710 104422 106720 104474
rect 106744 104422 106774 104474
rect 106774 104422 106786 104474
rect 106786 104422 106800 104474
rect 106824 104422 106838 104474
rect 106838 104422 106850 104474
rect 106850 104422 106880 104474
rect 106904 104422 106914 104474
rect 106914 104422 106960 104474
rect 106664 104420 106720 104422
rect 106744 104420 106800 104422
rect 106824 104420 106880 104422
rect 106904 104420 106960 104422
rect 105928 103930 105984 103932
rect 106008 103930 106064 103932
rect 106088 103930 106144 103932
rect 106168 103930 106224 103932
rect 105928 103878 105974 103930
rect 105974 103878 105984 103930
rect 106008 103878 106038 103930
rect 106038 103878 106050 103930
rect 106050 103878 106064 103930
rect 106088 103878 106102 103930
rect 106102 103878 106114 103930
rect 106114 103878 106144 103930
rect 106168 103878 106178 103930
rect 106178 103878 106224 103930
rect 105928 103876 105984 103878
rect 106008 103876 106064 103878
rect 106088 103876 106144 103878
rect 106168 103876 106224 103878
rect 106664 103386 106720 103388
rect 106744 103386 106800 103388
rect 106824 103386 106880 103388
rect 106904 103386 106960 103388
rect 106664 103334 106710 103386
rect 106710 103334 106720 103386
rect 106744 103334 106774 103386
rect 106774 103334 106786 103386
rect 106786 103334 106800 103386
rect 106824 103334 106838 103386
rect 106838 103334 106850 103386
rect 106850 103334 106880 103386
rect 106904 103334 106914 103386
rect 106914 103334 106960 103386
rect 106664 103332 106720 103334
rect 106744 103332 106800 103334
rect 106824 103332 106880 103334
rect 106904 103332 106960 103334
rect 105928 102842 105984 102844
rect 106008 102842 106064 102844
rect 106088 102842 106144 102844
rect 106168 102842 106224 102844
rect 105928 102790 105974 102842
rect 105974 102790 105984 102842
rect 106008 102790 106038 102842
rect 106038 102790 106050 102842
rect 106050 102790 106064 102842
rect 106088 102790 106102 102842
rect 106102 102790 106114 102842
rect 106114 102790 106144 102842
rect 106168 102790 106178 102842
rect 106178 102790 106224 102842
rect 105928 102788 105984 102790
rect 106008 102788 106064 102790
rect 106088 102788 106144 102790
rect 106168 102788 106224 102790
rect 106664 102298 106720 102300
rect 106744 102298 106800 102300
rect 106824 102298 106880 102300
rect 106904 102298 106960 102300
rect 106664 102246 106710 102298
rect 106710 102246 106720 102298
rect 106744 102246 106774 102298
rect 106774 102246 106786 102298
rect 106786 102246 106800 102298
rect 106824 102246 106838 102298
rect 106838 102246 106850 102298
rect 106850 102246 106880 102298
rect 106904 102246 106914 102298
rect 106914 102246 106960 102298
rect 106664 102244 106720 102246
rect 106744 102244 106800 102246
rect 106824 102244 106880 102246
rect 106904 102244 106960 102246
rect 105928 101754 105984 101756
rect 106008 101754 106064 101756
rect 106088 101754 106144 101756
rect 106168 101754 106224 101756
rect 105928 101702 105974 101754
rect 105974 101702 105984 101754
rect 106008 101702 106038 101754
rect 106038 101702 106050 101754
rect 106050 101702 106064 101754
rect 106088 101702 106102 101754
rect 106102 101702 106114 101754
rect 106114 101702 106144 101754
rect 106168 101702 106178 101754
rect 106178 101702 106224 101754
rect 105928 101700 105984 101702
rect 106008 101700 106064 101702
rect 106088 101700 106144 101702
rect 106168 101700 106224 101702
rect 106664 101210 106720 101212
rect 106744 101210 106800 101212
rect 106824 101210 106880 101212
rect 106904 101210 106960 101212
rect 106664 101158 106710 101210
rect 106710 101158 106720 101210
rect 106744 101158 106774 101210
rect 106774 101158 106786 101210
rect 106786 101158 106800 101210
rect 106824 101158 106838 101210
rect 106838 101158 106850 101210
rect 106850 101158 106880 101210
rect 106904 101158 106914 101210
rect 106914 101158 106960 101210
rect 106664 101156 106720 101158
rect 106744 101156 106800 101158
rect 106824 101156 106880 101158
rect 106904 101156 106960 101158
rect 105928 100666 105984 100668
rect 106008 100666 106064 100668
rect 106088 100666 106144 100668
rect 106168 100666 106224 100668
rect 105928 100614 105974 100666
rect 105974 100614 105984 100666
rect 106008 100614 106038 100666
rect 106038 100614 106050 100666
rect 106050 100614 106064 100666
rect 106088 100614 106102 100666
rect 106102 100614 106114 100666
rect 106114 100614 106144 100666
rect 106168 100614 106178 100666
rect 106178 100614 106224 100666
rect 105928 100612 105984 100614
rect 106008 100612 106064 100614
rect 106088 100612 106144 100614
rect 106168 100612 106224 100614
rect 106664 100122 106720 100124
rect 106744 100122 106800 100124
rect 106824 100122 106880 100124
rect 106904 100122 106960 100124
rect 106664 100070 106710 100122
rect 106710 100070 106720 100122
rect 106744 100070 106774 100122
rect 106774 100070 106786 100122
rect 106786 100070 106800 100122
rect 106824 100070 106838 100122
rect 106838 100070 106850 100122
rect 106850 100070 106880 100122
rect 106904 100070 106914 100122
rect 106914 100070 106960 100122
rect 106664 100068 106720 100070
rect 106744 100068 106800 100070
rect 106824 100068 106880 100070
rect 106904 100068 106960 100070
rect 105928 99578 105984 99580
rect 106008 99578 106064 99580
rect 106088 99578 106144 99580
rect 106168 99578 106224 99580
rect 105928 99526 105974 99578
rect 105974 99526 105984 99578
rect 106008 99526 106038 99578
rect 106038 99526 106050 99578
rect 106050 99526 106064 99578
rect 106088 99526 106102 99578
rect 106102 99526 106114 99578
rect 106114 99526 106144 99578
rect 106168 99526 106178 99578
rect 106178 99526 106224 99578
rect 105928 99524 105984 99526
rect 106008 99524 106064 99526
rect 106088 99524 106144 99526
rect 106168 99524 106224 99526
rect 106664 99034 106720 99036
rect 106744 99034 106800 99036
rect 106824 99034 106880 99036
rect 106904 99034 106960 99036
rect 106664 98982 106710 99034
rect 106710 98982 106720 99034
rect 106744 98982 106774 99034
rect 106774 98982 106786 99034
rect 106786 98982 106800 99034
rect 106824 98982 106838 99034
rect 106838 98982 106850 99034
rect 106850 98982 106880 99034
rect 106904 98982 106914 99034
rect 106914 98982 106960 99034
rect 106664 98980 106720 98982
rect 106744 98980 106800 98982
rect 106824 98980 106880 98982
rect 106904 98980 106960 98982
rect 105928 98490 105984 98492
rect 106008 98490 106064 98492
rect 106088 98490 106144 98492
rect 106168 98490 106224 98492
rect 105928 98438 105974 98490
rect 105974 98438 105984 98490
rect 106008 98438 106038 98490
rect 106038 98438 106050 98490
rect 106050 98438 106064 98490
rect 106088 98438 106102 98490
rect 106102 98438 106114 98490
rect 106114 98438 106144 98490
rect 106168 98438 106178 98490
rect 106178 98438 106224 98490
rect 105928 98436 105984 98438
rect 106008 98436 106064 98438
rect 106088 98436 106144 98438
rect 106168 98436 106224 98438
rect 106664 97946 106720 97948
rect 106744 97946 106800 97948
rect 106824 97946 106880 97948
rect 106904 97946 106960 97948
rect 106664 97894 106710 97946
rect 106710 97894 106720 97946
rect 106744 97894 106774 97946
rect 106774 97894 106786 97946
rect 106786 97894 106800 97946
rect 106824 97894 106838 97946
rect 106838 97894 106850 97946
rect 106850 97894 106880 97946
rect 106904 97894 106914 97946
rect 106914 97894 106960 97946
rect 106664 97892 106720 97894
rect 106744 97892 106800 97894
rect 106824 97892 106880 97894
rect 106904 97892 106960 97894
rect 105928 97402 105984 97404
rect 106008 97402 106064 97404
rect 106088 97402 106144 97404
rect 106168 97402 106224 97404
rect 105928 97350 105974 97402
rect 105974 97350 105984 97402
rect 106008 97350 106038 97402
rect 106038 97350 106050 97402
rect 106050 97350 106064 97402
rect 106088 97350 106102 97402
rect 106102 97350 106114 97402
rect 106114 97350 106144 97402
rect 106168 97350 106178 97402
rect 106178 97350 106224 97402
rect 105928 97348 105984 97350
rect 106008 97348 106064 97350
rect 106088 97348 106144 97350
rect 106168 97348 106224 97350
rect 106664 96858 106720 96860
rect 106744 96858 106800 96860
rect 106824 96858 106880 96860
rect 106904 96858 106960 96860
rect 106664 96806 106710 96858
rect 106710 96806 106720 96858
rect 106744 96806 106774 96858
rect 106774 96806 106786 96858
rect 106786 96806 106800 96858
rect 106824 96806 106838 96858
rect 106838 96806 106850 96858
rect 106850 96806 106880 96858
rect 106904 96806 106914 96858
rect 106914 96806 106960 96858
rect 106664 96804 106720 96806
rect 106744 96804 106800 96806
rect 106824 96804 106880 96806
rect 106904 96804 106960 96806
rect 105928 96314 105984 96316
rect 106008 96314 106064 96316
rect 106088 96314 106144 96316
rect 106168 96314 106224 96316
rect 105928 96262 105974 96314
rect 105974 96262 105984 96314
rect 106008 96262 106038 96314
rect 106038 96262 106050 96314
rect 106050 96262 106064 96314
rect 106088 96262 106102 96314
rect 106102 96262 106114 96314
rect 106114 96262 106144 96314
rect 106168 96262 106178 96314
rect 106178 96262 106224 96314
rect 105928 96260 105984 96262
rect 106008 96260 106064 96262
rect 106088 96260 106144 96262
rect 106168 96260 106224 96262
rect 106664 95770 106720 95772
rect 106744 95770 106800 95772
rect 106824 95770 106880 95772
rect 106904 95770 106960 95772
rect 106664 95718 106710 95770
rect 106710 95718 106720 95770
rect 106744 95718 106774 95770
rect 106774 95718 106786 95770
rect 106786 95718 106800 95770
rect 106824 95718 106838 95770
rect 106838 95718 106850 95770
rect 106850 95718 106880 95770
rect 106904 95718 106914 95770
rect 106914 95718 106960 95770
rect 106664 95716 106720 95718
rect 106744 95716 106800 95718
rect 106824 95716 106880 95718
rect 106904 95716 106960 95718
rect 105928 95226 105984 95228
rect 106008 95226 106064 95228
rect 106088 95226 106144 95228
rect 106168 95226 106224 95228
rect 105928 95174 105974 95226
rect 105974 95174 105984 95226
rect 106008 95174 106038 95226
rect 106038 95174 106050 95226
rect 106050 95174 106064 95226
rect 106088 95174 106102 95226
rect 106102 95174 106114 95226
rect 106114 95174 106144 95226
rect 106168 95174 106178 95226
rect 106178 95174 106224 95226
rect 105928 95172 105984 95174
rect 106008 95172 106064 95174
rect 106088 95172 106144 95174
rect 106168 95172 106224 95174
rect 106664 94682 106720 94684
rect 106744 94682 106800 94684
rect 106824 94682 106880 94684
rect 106904 94682 106960 94684
rect 106664 94630 106710 94682
rect 106710 94630 106720 94682
rect 106744 94630 106774 94682
rect 106774 94630 106786 94682
rect 106786 94630 106800 94682
rect 106824 94630 106838 94682
rect 106838 94630 106850 94682
rect 106850 94630 106880 94682
rect 106904 94630 106914 94682
rect 106914 94630 106960 94682
rect 106664 94628 106720 94630
rect 106744 94628 106800 94630
rect 106824 94628 106880 94630
rect 106904 94628 106960 94630
rect 105928 94138 105984 94140
rect 106008 94138 106064 94140
rect 106088 94138 106144 94140
rect 106168 94138 106224 94140
rect 105928 94086 105974 94138
rect 105974 94086 105984 94138
rect 106008 94086 106038 94138
rect 106038 94086 106050 94138
rect 106050 94086 106064 94138
rect 106088 94086 106102 94138
rect 106102 94086 106114 94138
rect 106114 94086 106144 94138
rect 106168 94086 106178 94138
rect 106178 94086 106224 94138
rect 105928 94084 105984 94086
rect 106008 94084 106064 94086
rect 106088 94084 106144 94086
rect 106168 94084 106224 94086
rect 106664 93594 106720 93596
rect 106744 93594 106800 93596
rect 106824 93594 106880 93596
rect 106904 93594 106960 93596
rect 106664 93542 106710 93594
rect 106710 93542 106720 93594
rect 106744 93542 106774 93594
rect 106774 93542 106786 93594
rect 106786 93542 106800 93594
rect 106824 93542 106838 93594
rect 106838 93542 106850 93594
rect 106850 93542 106880 93594
rect 106904 93542 106914 93594
rect 106914 93542 106960 93594
rect 106664 93540 106720 93542
rect 106744 93540 106800 93542
rect 106824 93540 106880 93542
rect 106904 93540 106960 93542
rect 105928 93050 105984 93052
rect 106008 93050 106064 93052
rect 106088 93050 106144 93052
rect 106168 93050 106224 93052
rect 105928 92998 105974 93050
rect 105974 92998 105984 93050
rect 106008 92998 106038 93050
rect 106038 92998 106050 93050
rect 106050 92998 106064 93050
rect 106088 92998 106102 93050
rect 106102 92998 106114 93050
rect 106114 92998 106144 93050
rect 106168 92998 106178 93050
rect 106178 92998 106224 93050
rect 105928 92996 105984 92998
rect 106008 92996 106064 92998
rect 106088 92996 106144 92998
rect 106168 92996 106224 92998
rect 106664 92506 106720 92508
rect 106744 92506 106800 92508
rect 106824 92506 106880 92508
rect 106904 92506 106960 92508
rect 106664 92454 106710 92506
rect 106710 92454 106720 92506
rect 106744 92454 106774 92506
rect 106774 92454 106786 92506
rect 106786 92454 106800 92506
rect 106824 92454 106838 92506
rect 106838 92454 106850 92506
rect 106850 92454 106880 92506
rect 106904 92454 106914 92506
rect 106914 92454 106960 92506
rect 106664 92452 106720 92454
rect 106744 92452 106800 92454
rect 106824 92452 106880 92454
rect 106904 92452 106960 92454
rect 105928 91962 105984 91964
rect 106008 91962 106064 91964
rect 106088 91962 106144 91964
rect 106168 91962 106224 91964
rect 105928 91910 105974 91962
rect 105974 91910 105984 91962
rect 106008 91910 106038 91962
rect 106038 91910 106050 91962
rect 106050 91910 106064 91962
rect 106088 91910 106102 91962
rect 106102 91910 106114 91962
rect 106114 91910 106144 91962
rect 106168 91910 106178 91962
rect 106178 91910 106224 91962
rect 105928 91908 105984 91910
rect 106008 91908 106064 91910
rect 106088 91908 106144 91910
rect 106168 91908 106224 91910
rect 106664 91418 106720 91420
rect 106744 91418 106800 91420
rect 106824 91418 106880 91420
rect 106904 91418 106960 91420
rect 106664 91366 106710 91418
rect 106710 91366 106720 91418
rect 106744 91366 106774 91418
rect 106774 91366 106786 91418
rect 106786 91366 106800 91418
rect 106824 91366 106838 91418
rect 106838 91366 106850 91418
rect 106850 91366 106880 91418
rect 106904 91366 106914 91418
rect 106914 91366 106960 91418
rect 106664 91364 106720 91366
rect 106744 91364 106800 91366
rect 106824 91364 106880 91366
rect 106904 91364 106960 91366
rect 105928 90874 105984 90876
rect 106008 90874 106064 90876
rect 106088 90874 106144 90876
rect 106168 90874 106224 90876
rect 105928 90822 105974 90874
rect 105974 90822 105984 90874
rect 106008 90822 106038 90874
rect 106038 90822 106050 90874
rect 106050 90822 106064 90874
rect 106088 90822 106102 90874
rect 106102 90822 106114 90874
rect 106114 90822 106144 90874
rect 106168 90822 106178 90874
rect 106178 90822 106224 90874
rect 105928 90820 105984 90822
rect 106008 90820 106064 90822
rect 106088 90820 106144 90822
rect 106168 90820 106224 90822
rect 106664 90330 106720 90332
rect 106744 90330 106800 90332
rect 106824 90330 106880 90332
rect 106904 90330 106960 90332
rect 106664 90278 106710 90330
rect 106710 90278 106720 90330
rect 106744 90278 106774 90330
rect 106774 90278 106786 90330
rect 106786 90278 106800 90330
rect 106824 90278 106838 90330
rect 106838 90278 106850 90330
rect 106850 90278 106880 90330
rect 106904 90278 106914 90330
rect 106914 90278 106960 90330
rect 106664 90276 106720 90278
rect 106744 90276 106800 90278
rect 106824 90276 106880 90278
rect 106904 90276 106960 90278
rect 105928 89786 105984 89788
rect 106008 89786 106064 89788
rect 106088 89786 106144 89788
rect 106168 89786 106224 89788
rect 105928 89734 105974 89786
rect 105974 89734 105984 89786
rect 106008 89734 106038 89786
rect 106038 89734 106050 89786
rect 106050 89734 106064 89786
rect 106088 89734 106102 89786
rect 106102 89734 106114 89786
rect 106114 89734 106144 89786
rect 106168 89734 106178 89786
rect 106178 89734 106224 89786
rect 105928 89732 105984 89734
rect 106008 89732 106064 89734
rect 106088 89732 106144 89734
rect 106168 89732 106224 89734
rect 106664 89242 106720 89244
rect 106744 89242 106800 89244
rect 106824 89242 106880 89244
rect 106904 89242 106960 89244
rect 106664 89190 106710 89242
rect 106710 89190 106720 89242
rect 106744 89190 106774 89242
rect 106774 89190 106786 89242
rect 106786 89190 106800 89242
rect 106824 89190 106838 89242
rect 106838 89190 106850 89242
rect 106850 89190 106880 89242
rect 106904 89190 106914 89242
rect 106914 89190 106960 89242
rect 106664 89188 106720 89190
rect 106744 89188 106800 89190
rect 106824 89188 106880 89190
rect 106904 89188 106960 89190
rect 105928 88698 105984 88700
rect 106008 88698 106064 88700
rect 106088 88698 106144 88700
rect 106168 88698 106224 88700
rect 105928 88646 105974 88698
rect 105974 88646 105984 88698
rect 106008 88646 106038 88698
rect 106038 88646 106050 88698
rect 106050 88646 106064 88698
rect 106088 88646 106102 88698
rect 106102 88646 106114 88698
rect 106114 88646 106144 88698
rect 106168 88646 106178 88698
rect 106178 88646 106224 88698
rect 105928 88644 105984 88646
rect 106008 88644 106064 88646
rect 106088 88644 106144 88646
rect 106168 88644 106224 88646
rect 106664 88154 106720 88156
rect 106744 88154 106800 88156
rect 106824 88154 106880 88156
rect 106904 88154 106960 88156
rect 106664 88102 106710 88154
rect 106710 88102 106720 88154
rect 106744 88102 106774 88154
rect 106774 88102 106786 88154
rect 106786 88102 106800 88154
rect 106824 88102 106838 88154
rect 106838 88102 106850 88154
rect 106850 88102 106880 88154
rect 106904 88102 106914 88154
rect 106914 88102 106960 88154
rect 106664 88100 106720 88102
rect 106744 88100 106800 88102
rect 106824 88100 106880 88102
rect 106904 88100 106960 88102
rect 105928 87610 105984 87612
rect 106008 87610 106064 87612
rect 106088 87610 106144 87612
rect 106168 87610 106224 87612
rect 105928 87558 105974 87610
rect 105974 87558 105984 87610
rect 106008 87558 106038 87610
rect 106038 87558 106050 87610
rect 106050 87558 106064 87610
rect 106088 87558 106102 87610
rect 106102 87558 106114 87610
rect 106114 87558 106144 87610
rect 106168 87558 106178 87610
rect 106178 87558 106224 87610
rect 105928 87556 105984 87558
rect 106008 87556 106064 87558
rect 106088 87556 106144 87558
rect 106168 87556 106224 87558
rect 106664 87066 106720 87068
rect 106744 87066 106800 87068
rect 106824 87066 106880 87068
rect 106904 87066 106960 87068
rect 106664 87014 106710 87066
rect 106710 87014 106720 87066
rect 106744 87014 106774 87066
rect 106774 87014 106786 87066
rect 106786 87014 106800 87066
rect 106824 87014 106838 87066
rect 106838 87014 106850 87066
rect 106850 87014 106880 87066
rect 106904 87014 106914 87066
rect 106914 87014 106960 87066
rect 106664 87012 106720 87014
rect 106744 87012 106800 87014
rect 106824 87012 106880 87014
rect 106904 87012 106960 87014
rect 105928 86522 105984 86524
rect 106008 86522 106064 86524
rect 106088 86522 106144 86524
rect 106168 86522 106224 86524
rect 105928 86470 105974 86522
rect 105974 86470 105984 86522
rect 106008 86470 106038 86522
rect 106038 86470 106050 86522
rect 106050 86470 106064 86522
rect 106088 86470 106102 86522
rect 106102 86470 106114 86522
rect 106114 86470 106144 86522
rect 106168 86470 106178 86522
rect 106178 86470 106224 86522
rect 105928 86468 105984 86470
rect 106008 86468 106064 86470
rect 106088 86468 106144 86470
rect 106168 86468 106224 86470
rect 106664 85978 106720 85980
rect 106744 85978 106800 85980
rect 106824 85978 106880 85980
rect 106904 85978 106960 85980
rect 106664 85926 106710 85978
rect 106710 85926 106720 85978
rect 106744 85926 106774 85978
rect 106774 85926 106786 85978
rect 106786 85926 106800 85978
rect 106824 85926 106838 85978
rect 106838 85926 106850 85978
rect 106850 85926 106880 85978
rect 106904 85926 106914 85978
rect 106914 85926 106960 85978
rect 106664 85924 106720 85926
rect 106744 85924 106800 85926
rect 106824 85924 106880 85926
rect 106904 85924 106960 85926
rect 104622 85040 104678 85096
rect 102322 66680 102378 66736
rect 71870 63824 71926 63880
rect 96158 63824 96214 63880
rect 104530 69808 104586 69864
rect 104346 67088 104402 67144
rect 102598 25100 102600 25120
rect 102600 25100 102652 25120
rect 102652 25100 102654 25120
rect 102322 25032 102378 25088
rect 102598 25064 102654 25100
rect 102046 23332 102102 23388
rect 9586 9832 9642 9888
rect 16118 9832 16174 9888
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 103978 59744 104034 59800
rect 105928 85434 105984 85436
rect 106008 85434 106064 85436
rect 106088 85434 106144 85436
rect 106168 85434 106224 85436
rect 105928 85382 105974 85434
rect 105974 85382 105984 85434
rect 106008 85382 106038 85434
rect 106038 85382 106050 85434
rect 106050 85382 106064 85434
rect 106088 85382 106102 85434
rect 106102 85382 106114 85434
rect 106114 85382 106144 85434
rect 106168 85382 106178 85434
rect 106178 85382 106224 85434
rect 105928 85380 105984 85382
rect 106008 85380 106064 85382
rect 106088 85380 106144 85382
rect 106168 85380 106224 85382
rect 106664 84890 106720 84892
rect 106744 84890 106800 84892
rect 106824 84890 106880 84892
rect 106904 84890 106960 84892
rect 106664 84838 106710 84890
rect 106710 84838 106720 84890
rect 106744 84838 106774 84890
rect 106774 84838 106786 84890
rect 106786 84838 106800 84890
rect 106824 84838 106838 84890
rect 106838 84838 106850 84890
rect 106850 84838 106880 84890
rect 106904 84838 106914 84890
rect 106914 84838 106960 84890
rect 106664 84836 106720 84838
rect 106744 84836 106800 84838
rect 106824 84836 106880 84838
rect 106904 84836 106960 84838
rect 105928 84346 105984 84348
rect 106008 84346 106064 84348
rect 106088 84346 106144 84348
rect 106168 84346 106224 84348
rect 105928 84294 105974 84346
rect 105974 84294 105984 84346
rect 106008 84294 106038 84346
rect 106038 84294 106050 84346
rect 106050 84294 106064 84346
rect 106088 84294 106102 84346
rect 106102 84294 106114 84346
rect 106114 84294 106144 84346
rect 106168 84294 106178 84346
rect 106178 84294 106224 84346
rect 105928 84292 105984 84294
rect 106008 84292 106064 84294
rect 106088 84292 106144 84294
rect 106168 84292 106224 84294
rect 106664 83802 106720 83804
rect 106744 83802 106800 83804
rect 106824 83802 106880 83804
rect 106904 83802 106960 83804
rect 106664 83750 106710 83802
rect 106710 83750 106720 83802
rect 106744 83750 106774 83802
rect 106774 83750 106786 83802
rect 106786 83750 106800 83802
rect 106824 83750 106838 83802
rect 106838 83750 106850 83802
rect 106850 83750 106880 83802
rect 106904 83750 106914 83802
rect 106914 83750 106960 83802
rect 106664 83748 106720 83750
rect 106744 83748 106800 83750
rect 106824 83748 106880 83750
rect 106904 83748 106960 83750
rect 105928 83258 105984 83260
rect 106008 83258 106064 83260
rect 106088 83258 106144 83260
rect 106168 83258 106224 83260
rect 105928 83206 105974 83258
rect 105974 83206 105984 83258
rect 106008 83206 106038 83258
rect 106038 83206 106050 83258
rect 106050 83206 106064 83258
rect 106088 83206 106102 83258
rect 106102 83206 106114 83258
rect 106114 83206 106144 83258
rect 106168 83206 106178 83258
rect 106178 83206 106224 83258
rect 105928 83204 105984 83206
rect 106008 83204 106064 83206
rect 106088 83204 106144 83206
rect 106168 83204 106224 83206
rect 106664 82714 106720 82716
rect 106744 82714 106800 82716
rect 106824 82714 106880 82716
rect 106904 82714 106960 82716
rect 106664 82662 106710 82714
rect 106710 82662 106720 82714
rect 106744 82662 106774 82714
rect 106774 82662 106786 82714
rect 106786 82662 106800 82714
rect 106824 82662 106838 82714
rect 106838 82662 106850 82714
rect 106850 82662 106880 82714
rect 106904 82662 106914 82714
rect 106914 82662 106960 82714
rect 106664 82660 106720 82662
rect 106744 82660 106800 82662
rect 106824 82660 106880 82662
rect 106904 82660 106960 82662
rect 105928 82170 105984 82172
rect 106008 82170 106064 82172
rect 106088 82170 106144 82172
rect 106168 82170 106224 82172
rect 105928 82118 105974 82170
rect 105974 82118 105984 82170
rect 106008 82118 106038 82170
rect 106038 82118 106050 82170
rect 106050 82118 106064 82170
rect 106088 82118 106102 82170
rect 106102 82118 106114 82170
rect 106114 82118 106144 82170
rect 106168 82118 106178 82170
rect 106178 82118 106224 82170
rect 105928 82116 105984 82118
rect 106008 82116 106064 82118
rect 106088 82116 106144 82118
rect 106168 82116 106224 82118
rect 106664 81626 106720 81628
rect 106744 81626 106800 81628
rect 106824 81626 106880 81628
rect 106904 81626 106960 81628
rect 106664 81574 106710 81626
rect 106710 81574 106720 81626
rect 106744 81574 106774 81626
rect 106774 81574 106786 81626
rect 106786 81574 106800 81626
rect 106824 81574 106838 81626
rect 106838 81574 106850 81626
rect 106850 81574 106880 81626
rect 106904 81574 106914 81626
rect 106914 81574 106960 81626
rect 106664 81572 106720 81574
rect 106744 81572 106800 81574
rect 106824 81572 106880 81574
rect 106904 81572 106960 81574
rect 105928 81082 105984 81084
rect 106008 81082 106064 81084
rect 106088 81082 106144 81084
rect 106168 81082 106224 81084
rect 105928 81030 105974 81082
rect 105974 81030 105984 81082
rect 106008 81030 106038 81082
rect 106038 81030 106050 81082
rect 106050 81030 106064 81082
rect 106088 81030 106102 81082
rect 106102 81030 106114 81082
rect 106114 81030 106144 81082
rect 106168 81030 106178 81082
rect 106178 81030 106224 81082
rect 105928 81028 105984 81030
rect 106008 81028 106064 81030
rect 106088 81028 106144 81030
rect 106168 81028 106224 81030
rect 106664 80538 106720 80540
rect 106744 80538 106800 80540
rect 106824 80538 106880 80540
rect 106904 80538 106960 80540
rect 106664 80486 106710 80538
rect 106710 80486 106720 80538
rect 106744 80486 106774 80538
rect 106774 80486 106786 80538
rect 106786 80486 106800 80538
rect 106824 80486 106838 80538
rect 106838 80486 106850 80538
rect 106850 80486 106880 80538
rect 106904 80486 106914 80538
rect 106914 80486 106960 80538
rect 106664 80484 106720 80486
rect 106744 80484 106800 80486
rect 106824 80484 106880 80486
rect 106904 80484 106960 80486
rect 105928 79994 105984 79996
rect 106008 79994 106064 79996
rect 106088 79994 106144 79996
rect 106168 79994 106224 79996
rect 105928 79942 105974 79994
rect 105974 79942 105984 79994
rect 106008 79942 106038 79994
rect 106038 79942 106050 79994
rect 106050 79942 106064 79994
rect 106088 79942 106102 79994
rect 106102 79942 106114 79994
rect 106114 79942 106144 79994
rect 106168 79942 106178 79994
rect 106178 79942 106224 79994
rect 105928 79940 105984 79942
rect 106008 79940 106064 79942
rect 106088 79940 106144 79942
rect 106168 79940 106224 79942
rect 106664 79450 106720 79452
rect 106744 79450 106800 79452
rect 106824 79450 106880 79452
rect 106904 79450 106960 79452
rect 106664 79398 106710 79450
rect 106710 79398 106720 79450
rect 106744 79398 106774 79450
rect 106774 79398 106786 79450
rect 106786 79398 106800 79450
rect 106824 79398 106838 79450
rect 106838 79398 106850 79450
rect 106850 79398 106880 79450
rect 106904 79398 106914 79450
rect 106914 79398 106960 79450
rect 106664 79396 106720 79398
rect 106744 79396 106800 79398
rect 106824 79396 106880 79398
rect 106904 79396 106960 79398
rect 105928 78906 105984 78908
rect 106008 78906 106064 78908
rect 106088 78906 106144 78908
rect 106168 78906 106224 78908
rect 105928 78854 105974 78906
rect 105974 78854 105984 78906
rect 106008 78854 106038 78906
rect 106038 78854 106050 78906
rect 106050 78854 106064 78906
rect 106088 78854 106102 78906
rect 106102 78854 106114 78906
rect 106114 78854 106144 78906
rect 106168 78854 106178 78906
rect 106178 78854 106224 78906
rect 105928 78852 105984 78854
rect 106008 78852 106064 78854
rect 106088 78852 106144 78854
rect 106168 78852 106224 78854
rect 106664 78362 106720 78364
rect 106744 78362 106800 78364
rect 106824 78362 106880 78364
rect 106904 78362 106960 78364
rect 106664 78310 106710 78362
rect 106710 78310 106720 78362
rect 106744 78310 106774 78362
rect 106774 78310 106786 78362
rect 106786 78310 106800 78362
rect 106824 78310 106838 78362
rect 106838 78310 106850 78362
rect 106850 78310 106880 78362
rect 106904 78310 106914 78362
rect 106914 78310 106960 78362
rect 106664 78308 106720 78310
rect 106744 78308 106800 78310
rect 106824 78308 106880 78310
rect 106904 78308 106960 78310
rect 105928 77818 105984 77820
rect 106008 77818 106064 77820
rect 106088 77818 106144 77820
rect 106168 77818 106224 77820
rect 105928 77766 105974 77818
rect 105974 77766 105984 77818
rect 106008 77766 106038 77818
rect 106038 77766 106050 77818
rect 106050 77766 106064 77818
rect 106088 77766 106102 77818
rect 106102 77766 106114 77818
rect 106114 77766 106144 77818
rect 106168 77766 106178 77818
rect 106178 77766 106224 77818
rect 105928 77764 105984 77766
rect 106008 77764 106064 77766
rect 106088 77764 106144 77766
rect 106168 77764 106224 77766
rect 105928 76730 105984 76732
rect 106008 76730 106064 76732
rect 106088 76730 106144 76732
rect 106168 76730 106224 76732
rect 105928 76678 105974 76730
rect 105974 76678 105984 76730
rect 106008 76678 106038 76730
rect 106038 76678 106050 76730
rect 106050 76678 106064 76730
rect 106088 76678 106102 76730
rect 106102 76678 106114 76730
rect 106114 76678 106144 76730
rect 106168 76678 106178 76730
rect 106178 76678 106224 76730
rect 105928 76676 105984 76678
rect 106008 76676 106064 76678
rect 106088 76676 106144 76678
rect 106168 76676 106224 76678
rect 106664 77274 106720 77276
rect 106744 77274 106800 77276
rect 106824 77274 106880 77276
rect 106904 77274 106960 77276
rect 106664 77222 106710 77274
rect 106710 77222 106720 77274
rect 106744 77222 106774 77274
rect 106774 77222 106786 77274
rect 106786 77222 106800 77274
rect 106824 77222 106838 77274
rect 106838 77222 106850 77274
rect 106850 77222 106880 77274
rect 106904 77222 106914 77274
rect 106914 77222 106960 77274
rect 106664 77220 106720 77222
rect 106744 77220 106800 77222
rect 106824 77220 106880 77222
rect 106904 77220 106960 77222
rect 106664 76186 106720 76188
rect 106744 76186 106800 76188
rect 106824 76186 106880 76188
rect 106904 76186 106960 76188
rect 106664 76134 106710 76186
rect 106710 76134 106720 76186
rect 106744 76134 106774 76186
rect 106774 76134 106786 76186
rect 106786 76134 106800 76186
rect 106824 76134 106838 76186
rect 106838 76134 106850 76186
rect 106850 76134 106880 76186
rect 106904 76134 106914 76186
rect 106914 76134 106960 76186
rect 106664 76132 106720 76134
rect 106744 76132 106800 76134
rect 106824 76132 106880 76134
rect 106904 76132 106960 76134
rect 105928 75642 105984 75644
rect 106008 75642 106064 75644
rect 106088 75642 106144 75644
rect 106168 75642 106224 75644
rect 105928 75590 105974 75642
rect 105974 75590 105984 75642
rect 106008 75590 106038 75642
rect 106038 75590 106050 75642
rect 106050 75590 106064 75642
rect 106088 75590 106102 75642
rect 106102 75590 106114 75642
rect 106114 75590 106144 75642
rect 106168 75590 106178 75642
rect 106178 75590 106224 75642
rect 105928 75588 105984 75590
rect 106008 75588 106064 75590
rect 106088 75588 106144 75590
rect 106168 75588 106224 75590
rect 106664 75098 106720 75100
rect 106744 75098 106800 75100
rect 106824 75098 106880 75100
rect 106904 75098 106960 75100
rect 106664 75046 106710 75098
rect 106710 75046 106720 75098
rect 106744 75046 106774 75098
rect 106774 75046 106786 75098
rect 106786 75046 106800 75098
rect 106824 75046 106838 75098
rect 106838 75046 106850 75098
rect 106850 75046 106880 75098
rect 106904 75046 106914 75098
rect 106914 75046 106960 75098
rect 106664 75044 106720 75046
rect 106744 75044 106800 75046
rect 106824 75044 106880 75046
rect 106904 75044 106960 75046
rect 105928 74554 105984 74556
rect 106008 74554 106064 74556
rect 106088 74554 106144 74556
rect 106168 74554 106224 74556
rect 105928 74502 105974 74554
rect 105974 74502 105984 74554
rect 106008 74502 106038 74554
rect 106038 74502 106050 74554
rect 106050 74502 106064 74554
rect 106088 74502 106102 74554
rect 106102 74502 106114 74554
rect 106114 74502 106144 74554
rect 106168 74502 106178 74554
rect 106178 74502 106224 74554
rect 105928 74500 105984 74502
rect 106008 74500 106064 74502
rect 106088 74500 106144 74502
rect 106168 74500 106224 74502
rect 106664 74010 106720 74012
rect 106744 74010 106800 74012
rect 106824 74010 106880 74012
rect 106904 74010 106960 74012
rect 106664 73958 106710 74010
rect 106710 73958 106720 74010
rect 106744 73958 106774 74010
rect 106774 73958 106786 74010
rect 106786 73958 106800 74010
rect 106824 73958 106838 74010
rect 106838 73958 106850 74010
rect 106850 73958 106880 74010
rect 106904 73958 106914 74010
rect 106914 73958 106960 74010
rect 106664 73956 106720 73958
rect 106744 73956 106800 73958
rect 106824 73956 106880 73958
rect 106904 73956 106960 73958
rect 105928 73466 105984 73468
rect 106008 73466 106064 73468
rect 106088 73466 106144 73468
rect 106168 73466 106224 73468
rect 105928 73414 105974 73466
rect 105974 73414 105984 73466
rect 106008 73414 106038 73466
rect 106038 73414 106050 73466
rect 106050 73414 106064 73466
rect 106088 73414 106102 73466
rect 106102 73414 106114 73466
rect 106114 73414 106144 73466
rect 106168 73414 106178 73466
rect 106178 73414 106224 73466
rect 105928 73412 105984 73414
rect 106008 73412 106064 73414
rect 106088 73412 106144 73414
rect 106168 73412 106224 73414
rect 106664 72922 106720 72924
rect 106744 72922 106800 72924
rect 106824 72922 106880 72924
rect 106904 72922 106960 72924
rect 106664 72870 106710 72922
rect 106710 72870 106720 72922
rect 106744 72870 106774 72922
rect 106774 72870 106786 72922
rect 106786 72870 106800 72922
rect 106824 72870 106838 72922
rect 106838 72870 106850 72922
rect 106850 72870 106880 72922
rect 106904 72870 106914 72922
rect 106914 72870 106960 72922
rect 106664 72868 106720 72870
rect 106744 72868 106800 72870
rect 106824 72868 106880 72870
rect 106904 72868 106960 72870
rect 105928 72378 105984 72380
rect 106008 72378 106064 72380
rect 106088 72378 106144 72380
rect 106168 72378 106224 72380
rect 105928 72326 105974 72378
rect 105974 72326 105984 72378
rect 106008 72326 106038 72378
rect 106038 72326 106050 72378
rect 106050 72326 106064 72378
rect 106088 72326 106102 72378
rect 106102 72326 106114 72378
rect 106114 72326 106144 72378
rect 106168 72326 106178 72378
rect 106178 72326 106224 72378
rect 105928 72324 105984 72326
rect 106008 72324 106064 72326
rect 106088 72324 106144 72326
rect 106168 72324 106224 72326
rect 106664 71834 106720 71836
rect 106744 71834 106800 71836
rect 106824 71834 106880 71836
rect 106904 71834 106960 71836
rect 106664 71782 106710 71834
rect 106710 71782 106720 71834
rect 106744 71782 106774 71834
rect 106774 71782 106786 71834
rect 106786 71782 106800 71834
rect 106824 71782 106838 71834
rect 106838 71782 106850 71834
rect 106850 71782 106880 71834
rect 106904 71782 106914 71834
rect 106914 71782 106960 71834
rect 106664 71780 106720 71782
rect 106744 71780 106800 71782
rect 106824 71780 106880 71782
rect 106904 71780 106960 71782
rect 105928 71290 105984 71292
rect 106008 71290 106064 71292
rect 106088 71290 106144 71292
rect 106168 71290 106224 71292
rect 105928 71238 105974 71290
rect 105974 71238 105984 71290
rect 106008 71238 106038 71290
rect 106038 71238 106050 71290
rect 106050 71238 106064 71290
rect 106088 71238 106102 71290
rect 106102 71238 106114 71290
rect 106114 71238 106144 71290
rect 106168 71238 106178 71290
rect 106178 71238 106224 71290
rect 105928 71236 105984 71238
rect 106008 71236 106064 71238
rect 106088 71236 106144 71238
rect 106168 71236 106224 71238
rect 106664 70746 106720 70748
rect 106744 70746 106800 70748
rect 106824 70746 106880 70748
rect 106904 70746 106960 70748
rect 106664 70694 106710 70746
rect 106710 70694 106720 70746
rect 106744 70694 106774 70746
rect 106774 70694 106786 70746
rect 106786 70694 106800 70746
rect 106824 70694 106838 70746
rect 106838 70694 106850 70746
rect 106850 70694 106880 70746
rect 106904 70694 106914 70746
rect 106914 70694 106960 70746
rect 106664 70692 106720 70694
rect 106744 70692 106800 70694
rect 106824 70692 106880 70694
rect 106904 70692 106960 70694
rect 105928 70202 105984 70204
rect 106008 70202 106064 70204
rect 106088 70202 106144 70204
rect 106168 70202 106224 70204
rect 105928 70150 105974 70202
rect 105974 70150 105984 70202
rect 106008 70150 106038 70202
rect 106038 70150 106050 70202
rect 106050 70150 106064 70202
rect 106088 70150 106102 70202
rect 106102 70150 106114 70202
rect 106114 70150 106144 70202
rect 106168 70150 106178 70202
rect 106178 70150 106224 70202
rect 105928 70148 105984 70150
rect 106008 70148 106064 70150
rect 106088 70148 106144 70150
rect 106168 70148 106224 70150
rect 106664 69658 106720 69660
rect 106744 69658 106800 69660
rect 106824 69658 106880 69660
rect 106904 69658 106960 69660
rect 106664 69606 106710 69658
rect 106710 69606 106720 69658
rect 106744 69606 106774 69658
rect 106774 69606 106786 69658
rect 106786 69606 106800 69658
rect 106824 69606 106838 69658
rect 106838 69606 106850 69658
rect 106850 69606 106880 69658
rect 106904 69606 106914 69658
rect 106914 69606 106960 69658
rect 106664 69604 106720 69606
rect 106744 69604 106800 69606
rect 106824 69604 106880 69606
rect 106904 69604 106960 69606
rect 105928 69114 105984 69116
rect 106008 69114 106064 69116
rect 106088 69114 106144 69116
rect 106168 69114 106224 69116
rect 105928 69062 105974 69114
rect 105974 69062 105984 69114
rect 106008 69062 106038 69114
rect 106038 69062 106050 69114
rect 106050 69062 106064 69114
rect 106088 69062 106102 69114
rect 106102 69062 106114 69114
rect 106114 69062 106144 69114
rect 106168 69062 106178 69114
rect 106178 69062 106224 69114
rect 105928 69060 105984 69062
rect 106008 69060 106064 69062
rect 106088 69060 106144 69062
rect 106168 69060 106224 69062
rect 106664 68570 106720 68572
rect 106744 68570 106800 68572
rect 106824 68570 106880 68572
rect 106904 68570 106960 68572
rect 106664 68518 106710 68570
rect 106710 68518 106720 68570
rect 106744 68518 106774 68570
rect 106774 68518 106786 68570
rect 106786 68518 106800 68570
rect 106824 68518 106838 68570
rect 106838 68518 106850 68570
rect 106850 68518 106880 68570
rect 106904 68518 106914 68570
rect 106914 68518 106960 68570
rect 106664 68516 106720 68518
rect 106744 68516 106800 68518
rect 106824 68516 106880 68518
rect 106904 68516 106960 68518
rect 105928 68026 105984 68028
rect 106008 68026 106064 68028
rect 106088 68026 106144 68028
rect 106168 68026 106224 68028
rect 105928 67974 105974 68026
rect 105974 67974 105984 68026
rect 106008 67974 106038 68026
rect 106038 67974 106050 68026
rect 106050 67974 106064 68026
rect 106088 67974 106102 68026
rect 106102 67974 106114 68026
rect 106114 67974 106144 68026
rect 106168 67974 106178 68026
rect 106178 67974 106224 68026
rect 105928 67972 105984 67974
rect 106008 67972 106064 67974
rect 106088 67972 106144 67974
rect 106168 67972 106224 67974
rect 106664 67482 106720 67484
rect 106744 67482 106800 67484
rect 106824 67482 106880 67484
rect 106904 67482 106960 67484
rect 106664 67430 106710 67482
rect 106710 67430 106720 67482
rect 106744 67430 106774 67482
rect 106774 67430 106786 67482
rect 106786 67430 106800 67482
rect 106824 67430 106838 67482
rect 106838 67430 106850 67482
rect 106850 67430 106880 67482
rect 106904 67430 106914 67482
rect 106914 67430 106960 67482
rect 106664 67428 106720 67430
rect 106744 67428 106800 67430
rect 106824 67428 106880 67430
rect 106904 67428 106960 67430
rect 106186 66544 106242 66600
rect 106664 66394 106720 66396
rect 106744 66394 106800 66396
rect 106824 66394 106880 66396
rect 106904 66394 106960 66396
rect 106664 66342 106710 66394
rect 106710 66342 106720 66394
rect 106744 66342 106774 66394
rect 106774 66342 106786 66394
rect 106786 66342 106800 66394
rect 106824 66342 106838 66394
rect 106838 66342 106850 66394
rect 106850 66342 106880 66394
rect 106904 66342 106914 66394
rect 106914 66342 106960 66394
rect 106664 66340 106720 66342
rect 106744 66340 106800 66342
rect 106824 66340 106880 66342
rect 106904 66340 106960 66342
rect 105928 65850 105984 65852
rect 106008 65850 106064 65852
rect 106088 65850 106144 65852
rect 106168 65850 106224 65852
rect 105928 65798 105974 65850
rect 105974 65798 105984 65850
rect 106008 65798 106038 65850
rect 106038 65798 106050 65850
rect 106050 65798 106064 65850
rect 106088 65798 106102 65850
rect 106102 65798 106114 65850
rect 106114 65798 106144 65850
rect 106168 65798 106178 65850
rect 106178 65798 106224 65850
rect 105928 65796 105984 65798
rect 106008 65796 106064 65798
rect 106088 65796 106144 65798
rect 106168 65796 106224 65798
rect 108486 69400 108542 69456
rect 108486 68720 108542 68776
rect 108486 68076 108488 68096
rect 108488 68076 108540 68096
rect 108540 68076 108542 68096
rect 108486 68040 108542 68076
rect 108486 67360 108542 67416
rect 108486 66680 108542 66736
rect 108486 66020 108542 66056
rect 108486 66000 108488 66020
rect 108488 66000 108540 66020
rect 108540 66000 108542 66020
rect 108486 65356 108488 65376
rect 108488 65356 108540 65376
rect 108540 65356 108542 65376
rect 108486 65320 108542 65356
rect 106664 65306 106720 65308
rect 106744 65306 106800 65308
rect 106824 65306 106880 65308
rect 106904 65306 106960 65308
rect 106664 65254 106710 65306
rect 106710 65254 106720 65306
rect 106744 65254 106774 65306
rect 106774 65254 106786 65306
rect 106786 65254 106800 65306
rect 106824 65254 106838 65306
rect 106838 65254 106850 65306
rect 106850 65254 106880 65306
rect 106904 65254 106914 65306
rect 106914 65254 106960 65306
rect 106664 65252 106720 65254
rect 106744 65252 106800 65254
rect 106824 65252 106880 65254
rect 106904 65252 106960 65254
rect 105928 64762 105984 64764
rect 106008 64762 106064 64764
rect 106088 64762 106144 64764
rect 106168 64762 106224 64764
rect 105928 64710 105974 64762
rect 105974 64710 105984 64762
rect 106008 64710 106038 64762
rect 106038 64710 106050 64762
rect 106050 64710 106064 64762
rect 106088 64710 106102 64762
rect 106102 64710 106114 64762
rect 106114 64710 106144 64762
rect 106168 64710 106178 64762
rect 106178 64710 106224 64762
rect 105928 64708 105984 64710
rect 106008 64708 106064 64710
rect 106088 64708 106144 64710
rect 106168 64708 106224 64710
rect 108486 64640 108542 64696
rect 106664 64218 106720 64220
rect 106744 64218 106800 64220
rect 106824 64218 106880 64220
rect 106904 64218 106960 64220
rect 106664 64166 106710 64218
rect 106710 64166 106720 64218
rect 106744 64166 106774 64218
rect 106774 64166 106786 64218
rect 106786 64166 106800 64218
rect 106824 64166 106838 64218
rect 106838 64166 106850 64218
rect 106850 64166 106880 64218
rect 106904 64166 106914 64218
rect 106914 64166 106960 64218
rect 106664 64164 106720 64166
rect 106744 64164 106800 64166
rect 106824 64164 106880 64166
rect 106904 64164 106960 64166
rect 108486 63960 108542 64016
rect 105634 63824 105690 63880
rect 105928 63674 105984 63676
rect 106008 63674 106064 63676
rect 106088 63674 106144 63676
rect 106168 63674 106224 63676
rect 105928 63622 105974 63674
rect 105974 63622 105984 63674
rect 106008 63622 106038 63674
rect 106038 63622 106050 63674
rect 106050 63622 106064 63674
rect 106088 63622 106102 63674
rect 106102 63622 106114 63674
rect 106114 63622 106144 63674
rect 106168 63622 106178 63674
rect 106178 63622 106224 63674
rect 105928 63620 105984 63622
rect 106008 63620 106064 63622
rect 106088 63620 106144 63622
rect 106168 63620 106224 63622
rect 106664 63130 106720 63132
rect 106744 63130 106800 63132
rect 106824 63130 106880 63132
rect 106904 63130 106960 63132
rect 106664 63078 106710 63130
rect 106710 63078 106720 63130
rect 106744 63078 106774 63130
rect 106774 63078 106786 63130
rect 106786 63078 106800 63130
rect 106824 63078 106838 63130
rect 106838 63078 106850 63130
rect 106850 63078 106880 63130
rect 106904 63078 106914 63130
rect 106914 63078 106960 63130
rect 106664 63076 106720 63078
rect 106744 63076 106800 63078
rect 106824 63076 106880 63078
rect 106904 63076 106960 63078
rect 105928 62586 105984 62588
rect 106008 62586 106064 62588
rect 106088 62586 106144 62588
rect 106168 62586 106224 62588
rect 105928 62534 105974 62586
rect 105974 62534 105984 62586
rect 106008 62534 106038 62586
rect 106038 62534 106050 62586
rect 106050 62534 106064 62586
rect 106088 62534 106102 62586
rect 106102 62534 106114 62586
rect 106114 62534 106144 62586
rect 106168 62534 106178 62586
rect 106178 62534 106224 62586
rect 105928 62532 105984 62534
rect 106008 62532 106064 62534
rect 106088 62532 106144 62534
rect 106168 62532 106224 62534
rect 106664 62042 106720 62044
rect 106744 62042 106800 62044
rect 106824 62042 106880 62044
rect 106904 62042 106960 62044
rect 106664 61990 106710 62042
rect 106710 61990 106720 62042
rect 106744 61990 106774 62042
rect 106774 61990 106786 62042
rect 106786 61990 106800 62042
rect 106824 61990 106838 62042
rect 106838 61990 106850 62042
rect 106850 61990 106880 62042
rect 106904 61990 106914 62042
rect 106914 61990 106960 62042
rect 106664 61988 106720 61990
rect 106744 61988 106800 61990
rect 106824 61988 106880 61990
rect 106904 61988 106960 61990
rect 105928 61498 105984 61500
rect 106008 61498 106064 61500
rect 106088 61498 106144 61500
rect 106168 61498 106224 61500
rect 105928 61446 105974 61498
rect 105974 61446 105984 61498
rect 106008 61446 106038 61498
rect 106038 61446 106050 61498
rect 106050 61446 106064 61498
rect 106088 61446 106102 61498
rect 106102 61446 106114 61498
rect 106114 61446 106144 61498
rect 106168 61446 106178 61498
rect 106178 61446 106224 61498
rect 105928 61444 105984 61446
rect 106008 61444 106064 61446
rect 106088 61444 106144 61446
rect 106168 61444 106224 61446
rect 106664 60954 106720 60956
rect 106744 60954 106800 60956
rect 106824 60954 106880 60956
rect 106904 60954 106960 60956
rect 106664 60902 106710 60954
rect 106710 60902 106720 60954
rect 106744 60902 106774 60954
rect 106774 60902 106786 60954
rect 106786 60902 106800 60954
rect 106824 60902 106838 60954
rect 106838 60902 106850 60954
rect 106850 60902 106880 60954
rect 106904 60902 106914 60954
rect 106914 60902 106960 60954
rect 106664 60900 106720 60902
rect 106744 60900 106800 60902
rect 106824 60900 106880 60902
rect 106904 60900 106960 60902
rect 105928 60410 105984 60412
rect 106008 60410 106064 60412
rect 106088 60410 106144 60412
rect 106168 60410 106224 60412
rect 105928 60358 105974 60410
rect 105974 60358 105984 60410
rect 106008 60358 106038 60410
rect 106038 60358 106050 60410
rect 106050 60358 106064 60410
rect 106088 60358 106102 60410
rect 106102 60358 106114 60410
rect 106114 60358 106144 60410
rect 106168 60358 106178 60410
rect 106178 60358 106224 60410
rect 105928 60356 105984 60358
rect 106008 60356 106064 60358
rect 106088 60356 106144 60358
rect 106168 60356 106224 60358
rect 106664 59866 106720 59868
rect 106744 59866 106800 59868
rect 106824 59866 106880 59868
rect 106904 59866 106960 59868
rect 106664 59814 106710 59866
rect 106710 59814 106720 59866
rect 106744 59814 106774 59866
rect 106774 59814 106786 59866
rect 106786 59814 106800 59866
rect 106824 59814 106838 59866
rect 106838 59814 106850 59866
rect 106850 59814 106880 59866
rect 106904 59814 106914 59866
rect 106914 59814 106960 59866
rect 106664 59812 106720 59814
rect 106744 59812 106800 59814
rect 106824 59812 106880 59814
rect 106904 59812 106960 59814
rect 105928 59322 105984 59324
rect 106008 59322 106064 59324
rect 106088 59322 106144 59324
rect 106168 59322 106224 59324
rect 105928 59270 105974 59322
rect 105974 59270 105984 59322
rect 106008 59270 106038 59322
rect 106038 59270 106050 59322
rect 106050 59270 106064 59322
rect 106088 59270 106102 59322
rect 106102 59270 106114 59322
rect 106114 59270 106144 59322
rect 106168 59270 106178 59322
rect 106178 59270 106224 59322
rect 105928 59268 105984 59270
rect 106008 59268 106064 59270
rect 106088 59268 106144 59270
rect 106168 59268 106224 59270
rect 106664 58778 106720 58780
rect 106744 58778 106800 58780
rect 106824 58778 106880 58780
rect 106904 58778 106960 58780
rect 106664 58726 106710 58778
rect 106710 58726 106720 58778
rect 106744 58726 106774 58778
rect 106774 58726 106786 58778
rect 106786 58726 106800 58778
rect 106824 58726 106838 58778
rect 106838 58726 106850 58778
rect 106850 58726 106880 58778
rect 106904 58726 106914 58778
rect 106914 58726 106960 58778
rect 106664 58724 106720 58726
rect 106744 58724 106800 58726
rect 106824 58724 106880 58726
rect 106904 58724 106960 58726
rect 104346 22208 104402 22264
rect 105928 58234 105984 58236
rect 106008 58234 106064 58236
rect 106088 58234 106144 58236
rect 106168 58234 106224 58236
rect 105928 58182 105974 58234
rect 105974 58182 105984 58234
rect 106008 58182 106038 58234
rect 106038 58182 106050 58234
rect 106050 58182 106064 58234
rect 106088 58182 106102 58234
rect 106102 58182 106114 58234
rect 106114 58182 106144 58234
rect 106168 58182 106178 58234
rect 106178 58182 106224 58234
rect 105928 58180 105984 58182
rect 106008 58180 106064 58182
rect 106088 58180 106144 58182
rect 106168 58180 106224 58182
rect 106664 57690 106720 57692
rect 106744 57690 106800 57692
rect 106824 57690 106880 57692
rect 106904 57690 106960 57692
rect 106664 57638 106710 57690
rect 106710 57638 106720 57690
rect 106744 57638 106774 57690
rect 106774 57638 106786 57690
rect 106786 57638 106800 57690
rect 106824 57638 106838 57690
rect 106838 57638 106850 57690
rect 106850 57638 106880 57690
rect 106904 57638 106914 57690
rect 106914 57638 106960 57690
rect 106664 57636 106720 57638
rect 106744 57636 106800 57638
rect 106824 57636 106880 57638
rect 106904 57636 106960 57638
rect 105928 57146 105984 57148
rect 106008 57146 106064 57148
rect 106088 57146 106144 57148
rect 106168 57146 106224 57148
rect 105928 57094 105974 57146
rect 105974 57094 105984 57146
rect 106008 57094 106038 57146
rect 106038 57094 106050 57146
rect 106050 57094 106064 57146
rect 106088 57094 106102 57146
rect 106102 57094 106114 57146
rect 106114 57094 106144 57146
rect 106168 57094 106178 57146
rect 106178 57094 106224 57146
rect 105928 57092 105984 57094
rect 106008 57092 106064 57094
rect 106088 57092 106144 57094
rect 106168 57092 106224 57094
rect 106664 56602 106720 56604
rect 106744 56602 106800 56604
rect 106824 56602 106880 56604
rect 106904 56602 106960 56604
rect 106664 56550 106710 56602
rect 106710 56550 106720 56602
rect 106744 56550 106774 56602
rect 106774 56550 106786 56602
rect 106786 56550 106800 56602
rect 106824 56550 106838 56602
rect 106838 56550 106850 56602
rect 106850 56550 106880 56602
rect 106904 56550 106914 56602
rect 106914 56550 106960 56602
rect 106664 56548 106720 56550
rect 106744 56548 106800 56550
rect 106824 56548 106880 56550
rect 106904 56548 106960 56550
rect 105928 56058 105984 56060
rect 106008 56058 106064 56060
rect 106088 56058 106144 56060
rect 106168 56058 106224 56060
rect 105928 56006 105974 56058
rect 105974 56006 105984 56058
rect 106008 56006 106038 56058
rect 106038 56006 106050 56058
rect 106050 56006 106064 56058
rect 106088 56006 106102 56058
rect 106102 56006 106114 56058
rect 106114 56006 106144 56058
rect 106168 56006 106178 56058
rect 106178 56006 106224 56058
rect 105928 56004 105984 56006
rect 106008 56004 106064 56006
rect 106088 56004 106144 56006
rect 106168 56004 106224 56006
rect 106664 55514 106720 55516
rect 106744 55514 106800 55516
rect 106824 55514 106880 55516
rect 106904 55514 106960 55516
rect 106664 55462 106710 55514
rect 106710 55462 106720 55514
rect 106744 55462 106774 55514
rect 106774 55462 106786 55514
rect 106786 55462 106800 55514
rect 106824 55462 106838 55514
rect 106838 55462 106850 55514
rect 106850 55462 106880 55514
rect 106904 55462 106914 55514
rect 106914 55462 106960 55514
rect 106664 55460 106720 55462
rect 106744 55460 106800 55462
rect 106824 55460 106880 55462
rect 106904 55460 106960 55462
rect 105928 54970 105984 54972
rect 106008 54970 106064 54972
rect 106088 54970 106144 54972
rect 106168 54970 106224 54972
rect 105928 54918 105974 54970
rect 105974 54918 105984 54970
rect 106008 54918 106038 54970
rect 106038 54918 106050 54970
rect 106050 54918 106064 54970
rect 106088 54918 106102 54970
rect 106102 54918 106114 54970
rect 106114 54918 106144 54970
rect 106168 54918 106178 54970
rect 106178 54918 106224 54970
rect 105928 54916 105984 54918
rect 106008 54916 106064 54918
rect 106088 54916 106144 54918
rect 106168 54916 106224 54918
rect 106664 54426 106720 54428
rect 106744 54426 106800 54428
rect 106824 54426 106880 54428
rect 106904 54426 106960 54428
rect 106664 54374 106710 54426
rect 106710 54374 106720 54426
rect 106744 54374 106774 54426
rect 106774 54374 106786 54426
rect 106786 54374 106800 54426
rect 106824 54374 106838 54426
rect 106838 54374 106850 54426
rect 106850 54374 106880 54426
rect 106904 54374 106914 54426
rect 106914 54374 106960 54426
rect 106664 54372 106720 54374
rect 106744 54372 106800 54374
rect 106824 54372 106880 54374
rect 106904 54372 106960 54374
rect 105928 53882 105984 53884
rect 106008 53882 106064 53884
rect 106088 53882 106144 53884
rect 106168 53882 106224 53884
rect 105928 53830 105974 53882
rect 105974 53830 105984 53882
rect 106008 53830 106038 53882
rect 106038 53830 106050 53882
rect 106050 53830 106064 53882
rect 106088 53830 106102 53882
rect 106102 53830 106114 53882
rect 106114 53830 106144 53882
rect 106168 53830 106178 53882
rect 106178 53830 106224 53882
rect 105928 53828 105984 53830
rect 106008 53828 106064 53830
rect 106088 53828 106144 53830
rect 106168 53828 106224 53830
rect 106664 53338 106720 53340
rect 106744 53338 106800 53340
rect 106824 53338 106880 53340
rect 106904 53338 106960 53340
rect 106664 53286 106710 53338
rect 106710 53286 106720 53338
rect 106744 53286 106774 53338
rect 106774 53286 106786 53338
rect 106786 53286 106800 53338
rect 106824 53286 106838 53338
rect 106838 53286 106850 53338
rect 106850 53286 106880 53338
rect 106904 53286 106914 53338
rect 106914 53286 106960 53338
rect 106664 53284 106720 53286
rect 106744 53284 106800 53286
rect 106824 53284 106880 53286
rect 106904 53284 106960 53286
rect 105928 52794 105984 52796
rect 106008 52794 106064 52796
rect 106088 52794 106144 52796
rect 106168 52794 106224 52796
rect 105928 52742 105974 52794
rect 105974 52742 105984 52794
rect 106008 52742 106038 52794
rect 106038 52742 106050 52794
rect 106050 52742 106064 52794
rect 106088 52742 106102 52794
rect 106102 52742 106114 52794
rect 106114 52742 106144 52794
rect 106168 52742 106178 52794
rect 106178 52742 106224 52794
rect 105928 52740 105984 52742
rect 106008 52740 106064 52742
rect 106088 52740 106144 52742
rect 106168 52740 106224 52742
rect 106664 52250 106720 52252
rect 106744 52250 106800 52252
rect 106824 52250 106880 52252
rect 106904 52250 106960 52252
rect 106664 52198 106710 52250
rect 106710 52198 106720 52250
rect 106744 52198 106774 52250
rect 106774 52198 106786 52250
rect 106786 52198 106800 52250
rect 106824 52198 106838 52250
rect 106838 52198 106850 52250
rect 106850 52198 106880 52250
rect 106904 52198 106914 52250
rect 106914 52198 106960 52250
rect 106664 52196 106720 52198
rect 106744 52196 106800 52198
rect 106824 52196 106880 52198
rect 106904 52196 106960 52198
rect 105928 51706 105984 51708
rect 106008 51706 106064 51708
rect 106088 51706 106144 51708
rect 106168 51706 106224 51708
rect 105928 51654 105974 51706
rect 105974 51654 105984 51706
rect 106008 51654 106038 51706
rect 106038 51654 106050 51706
rect 106050 51654 106064 51706
rect 106088 51654 106102 51706
rect 106102 51654 106114 51706
rect 106114 51654 106144 51706
rect 106168 51654 106178 51706
rect 106178 51654 106224 51706
rect 105928 51652 105984 51654
rect 106008 51652 106064 51654
rect 106088 51652 106144 51654
rect 106168 51652 106224 51654
rect 106664 51162 106720 51164
rect 106744 51162 106800 51164
rect 106824 51162 106880 51164
rect 106904 51162 106960 51164
rect 106664 51110 106710 51162
rect 106710 51110 106720 51162
rect 106744 51110 106774 51162
rect 106774 51110 106786 51162
rect 106786 51110 106800 51162
rect 106824 51110 106838 51162
rect 106838 51110 106850 51162
rect 106850 51110 106880 51162
rect 106904 51110 106914 51162
rect 106914 51110 106960 51162
rect 106664 51108 106720 51110
rect 106744 51108 106800 51110
rect 106824 51108 106880 51110
rect 106904 51108 106960 51110
rect 105928 50618 105984 50620
rect 106008 50618 106064 50620
rect 106088 50618 106144 50620
rect 106168 50618 106224 50620
rect 105928 50566 105974 50618
rect 105974 50566 105984 50618
rect 106008 50566 106038 50618
rect 106038 50566 106050 50618
rect 106050 50566 106064 50618
rect 106088 50566 106102 50618
rect 106102 50566 106114 50618
rect 106114 50566 106144 50618
rect 106168 50566 106178 50618
rect 106178 50566 106224 50618
rect 105928 50564 105984 50566
rect 106008 50564 106064 50566
rect 106088 50564 106144 50566
rect 106168 50564 106224 50566
rect 106664 50074 106720 50076
rect 106744 50074 106800 50076
rect 106824 50074 106880 50076
rect 106904 50074 106960 50076
rect 106664 50022 106710 50074
rect 106710 50022 106720 50074
rect 106744 50022 106774 50074
rect 106774 50022 106786 50074
rect 106786 50022 106800 50074
rect 106824 50022 106838 50074
rect 106838 50022 106850 50074
rect 106850 50022 106880 50074
rect 106904 50022 106914 50074
rect 106914 50022 106960 50074
rect 106664 50020 106720 50022
rect 106744 50020 106800 50022
rect 106824 50020 106880 50022
rect 106904 50020 106960 50022
rect 105928 49530 105984 49532
rect 106008 49530 106064 49532
rect 106088 49530 106144 49532
rect 106168 49530 106224 49532
rect 105928 49478 105974 49530
rect 105974 49478 105984 49530
rect 106008 49478 106038 49530
rect 106038 49478 106050 49530
rect 106050 49478 106064 49530
rect 106088 49478 106102 49530
rect 106102 49478 106114 49530
rect 106114 49478 106144 49530
rect 106168 49478 106178 49530
rect 106178 49478 106224 49530
rect 105928 49476 105984 49478
rect 106008 49476 106064 49478
rect 106088 49476 106144 49478
rect 106168 49476 106224 49478
rect 106664 48986 106720 48988
rect 106744 48986 106800 48988
rect 106824 48986 106880 48988
rect 106904 48986 106960 48988
rect 106664 48934 106710 48986
rect 106710 48934 106720 48986
rect 106744 48934 106774 48986
rect 106774 48934 106786 48986
rect 106786 48934 106800 48986
rect 106824 48934 106838 48986
rect 106838 48934 106850 48986
rect 106850 48934 106880 48986
rect 106904 48934 106914 48986
rect 106914 48934 106960 48986
rect 106664 48932 106720 48934
rect 106744 48932 106800 48934
rect 106824 48932 106880 48934
rect 106904 48932 106960 48934
rect 105928 48442 105984 48444
rect 106008 48442 106064 48444
rect 106088 48442 106144 48444
rect 106168 48442 106224 48444
rect 105928 48390 105974 48442
rect 105974 48390 105984 48442
rect 106008 48390 106038 48442
rect 106038 48390 106050 48442
rect 106050 48390 106064 48442
rect 106088 48390 106102 48442
rect 106102 48390 106114 48442
rect 106114 48390 106144 48442
rect 106168 48390 106178 48442
rect 106178 48390 106224 48442
rect 105928 48388 105984 48390
rect 106008 48388 106064 48390
rect 106088 48388 106144 48390
rect 106168 48388 106224 48390
rect 106664 47898 106720 47900
rect 106744 47898 106800 47900
rect 106824 47898 106880 47900
rect 106904 47898 106960 47900
rect 106664 47846 106710 47898
rect 106710 47846 106720 47898
rect 106744 47846 106774 47898
rect 106774 47846 106786 47898
rect 106786 47846 106800 47898
rect 106824 47846 106838 47898
rect 106838 47846 106850 47898
rect 106850 47846 106880 47898
rect 106904 47846 106914 47898
rect 106914 47846 106960 47898
rect 106664 47844 106720 47846
rect 106744 47844 106800 47846
rect 106824 47844 106880 47846
rect 106904 47844 106960 47846
rect 105928 47354 105984 47356
rect 106008 47354 106064 47356
rect 106088 47354 106144 47356
rect 106168 47354 106224 47356
rect 105928 47302 105974 47354
rect 105974 47302 105984 47354
rect 106008 47302 106038 47354
rect 106038 47302 106050 47354
rect 106050 47302 106064 47354
rect 106088 47302 106102 47354
rect 106102 47302 106114 47354
rect 106114 47302 106144 47354
rect 106168 47302 106178 47354
rect 106178 47302 106224 47354
rect 105928 47300 105984 47302
rect 106008 47300 106064 47302
rect 106088 47300 106144 47302
rect 106168 47300 106224 47302
rect 106664 46810 106720 46812
rect 106744 46810 106800 46812
rect 106824 46810 106880 46812
rect 106904 46810 106960 46812
rect 106664 46758 106710 46810
rect 106710 46758 106720 46810
rect 106744 46758 106774 46810
rect 106774 46758 106786 46810
rect 106786 46758 106800 46810
rect 106824 46758 106838 46810
rect 106838 46758 106850 46810
rect 106850 46758 106880 46810
rect 106904 46758 106914 46810
rect 106914 46758 106960 46810
rect 106664 46756 106720 46758
rect 106744 46756 106800 46758
rect 106824 46756 106880 46758
rect 106904 46756 106960 46758
rect 105928 46266 105984 46268
rect 106008 46266 106064 46268
rect 106088 46266 106144 46268
rect 106168 46266 106224 46268
rect 105928 46214 105974 46266
rect 105974 46214 105984 46266
rect 106008 46214 106038 46266
rect 106038 46214 106050 46266
rect 106050 46214 106064 46266
rect 106088 46214 106102 46266
rect 106102 46214 106114 46266
rect 106114 46214 106144 46266
rect 106168 46214 106178 46266
rect 106178 46214 106224 46266
rect 105928 46212 105984 46214
rect 106008 46212 106064 46214
rect 106088 46212 106144 46214
rect 106168 46212 106224 46214
rect 106664 45722 106720 45724
rect 106744 45722 106800 45724
rect 106824 45722 106880 45724
rect 106904 45722 106960 45724
rect 106664 45670 106710 45722
rect 106710 45670 106720 45722
rect 106744 45670 106774 45722
rect 106774 45670 106786 45722
rect 106786 45670 106800 45722
rect 106824 45670 106838 45722
rect 106838 45670 106850 45722
rect 106850 45670 106880 45722
rect 106904 45670 106914 45722
rect 106914 45670 106960 45722
rect 106664 45668 106720 45670
rect 106744 45668 106800 45670
rect 106824 45668 106880 45670
rect 106904 45668 106960 45670
rect 105928 45178 105984 45180
rect 106008 45178 106064 45180
rect 106088 45178 106144 45180
rect 106168 45178 106224 45180
rect 105928 45126 105974 45178
rect 105974 45126 105984 45178
rect 106008 45126 106038 45178
rect 106038 45126 106050 45178
rect 106050 45126 106064 45178
rect 106088 45126 106102 45178
rect 106102 45126 106114 45178
rect 106114 45126 106144 45178
rect 106168 45126 106178 45178
rect 106178 45126 106224 45178
rect 105928 45124 105984 45126
rect 106008 45124 106064 45126
rect 106088 45124 106144 45126
rect 106168 45124 106224 45126
rect 108486 51040 108542 51096
rect 106664 44634 106720 44636
rect 106744 44634 106800 44636
rect 106824 44634 106880 44636
rect 106904 44634 106960 44636
rect 106664 44582 106710 44634
rect 106710 44582 106720 44634
rect 106744 44582 106774 44634
rect 106774 44582 106786 44634
rect 106786 44582 106800 44634
rect 106824 44582 106838 44634
rect 106838 44582 106850 44634
rect 106850 44582 106880 44634
rect 106904 44582 106914 44634
rect 106914 44582 106960 44634
rect 106664 44580 106720 44582
rect 106744 44580 106800 44582
rect 106824 44580 106880 44582
rect 106904 44580 106960 44582
rect 105928 44090 105984 44092
rect 106008 44090 106064 44092
rect 106088 44090 106144 44092
rect 106168 44090 106224 44092
rect 105928 44038 105974 44090
rect 105974 44038 105984 44090
rect 106008 44038 106038 44090
rect 106038 44038 106050 44090
rect 106050 44038 106064 44090
rect 106088 44038 106102 44090
rect 106102 44038 106114 44090
rect 106114 44038 106144 44090
rect 106168 44038 106178 44090
rect 106178 44038 106224 44090
rect 105928 44036 105984 44038
rect 106008 44036 106064 44038
rect 106088 44036 106144 44038
rect 106168 44036 106224 44038
rect 106664 43546 106720 43548
rect 106744 43546 106800 43548
rect 106824 43546 106880 43548
rect 106904 43546 106960 43548
rect 106664 43494 106710 43546
rect 106710 43494 106720 43546
rect 106744 43494 106774 43546
rect 106774 43494 106786 43546
rect 106786 43494 106800 43546
rect 106824 43494 106838 43546
rect 106838 43494 106850 43546
rect 106850 43494 106880 43546
rect 106904 43494 106914 43546
rect 106914 43494 106960 43546
rect 106664 43492 106720 43494
rect 106744 43492 106800 43494
rect 106824 43492 106880 43494
rect 106904 43492 106960 43494
rect 105928 43002 105984 43004
rect 106008 43002 106064 43004
rect 106088 43002 106144 43004
rect 106168 43002 106224 43004
rect 105928 42950 105974 43002
rect 105974 42950 105984 43002
rect 106008 42950 106038 43002
rect 106038 42950 106050 43002
rect 106050 42950 106064 43002
rect 106088 42950 106102 43002
rect 106102 42950 106114 43002
rect 106114 42950 106144 43002
rect 106168 42950 106178 43002
rect 106178 42950 106224 43002
rect 105928 42948 105984 42950
rect 106008 42948 106064 42950
rect 106088 42948 106144 42950
rect 106168 42948 106224 42950
rect 106664 42458 106720 42460
rect 106744 42458 106800 42460
rect 106824 42458 106880 42460
rect 106904 42458 106960 42460
rect 106664 42406 106710 42458
rect 106710 42406 106720 42458
rect 106744 42406 106774 42458
rect 106774 42406 106786 42458
rect 106786 42406 106800 42458
rect 106824 42406 106838 42458
rect 106838 42406 106850 42458
rect 106850 42406 106880 42458
rect 106904 42406 106914 42458
rect 106914 42406 106960 42458
rect 106664 42404 106720 42406
rect 106744 42404 106800 42406
rect 106824 42404 106880 42406
rect 106904 42404 106960 42406
rect 105928 41914 105984 41916
rect 106008 41914 106064 41916
rect 106088 41914 106144 41916
rect 106168 41914 106224 41916
rect 105928 41862 105974 41914
rect 105974 41862 105984 41914
rect 106008 41862 106038 41914
rect 106038 41862 106050 41914
rect 106050 41862 106064 41914
rect 106088 41862 106102 41914
rect 106102 41862 106114 41914
rect 106114 41862 106144 41914
rect 106168 41862 106178 41914
rect 106178 41862 106224 41914
rect 105928 41860 105984 41862
rect 106008 41860 106064 41862
rect 106088 41860 106144 41862
rect 106168 41860 106224 41862
rect 106664 41370 106720 41372
rect 106744 41370 106800 41372
rect 106824 41370 106880 41372
rect 106904 41370 106960 41372
rect 106664 41318 106710 41370
rect 106710 41318 106720 41370
rect 106744 41318 106774 41370
rect 106774 41318 106786 41370
rect 106786 41318 106800 41370
rect 106824 41318 106838 41370
rect 106838 41318 106850 41370
rect 106850 41318 106880 41370
rect 106904 41318 106914 41370
rect 106914 41318 106960 41370
rect 106664 41316 106720 41318
rect 106744 41316 106800 41318
rect 106824 41316 106880 41318
rect 106904 41316 106960 41318
rect 105928 40826 105984 40828
rect 106008 40826 106064 40828
rect 106088 40826 106144 40828
rect 106168 40826 106224 40828
rect 105928 40774 105974 40826
rect 105974 40774 105984 40826
rect 106008 40774 106038 40826
rect 106038 40774 106050 40826
rect 106050 40774 106064 40826
rect 106088 40774 106102 40826
rect 106102 40774 106114 40826
rect 106114 40774 106144 40826
rect 106168 40774 106178 40826
rect 106178 40774 106224 40826
rect 105928 40772 105984 40774
rect 106008 40772 106064 40774
rect 106088 40772 106144 40774
rect 106168 40772 106224 40774
rect 106664 40282 106720 40284
rect 106744 40282 106800 40284
rect 106824 40282 106880 40284
rect 106904 40282 106960 40284
rect 106664 40230 106710 40282
rect 106710 40230 106720 40282
rect 106744 40230 106774 40282
rect 106774 40230 106786 40282
rect 106786 40230 106800 40282
rect 106824 40230 106838 40282
rect 106838 40230 106850 40282
rect 106850 40230 106880 40282
rect 106904 40230 106914 40282
rect 106914 40230 106960 40282
rect 106664 40228 106720 40230
rect 106744 40228 106800 40230
rect 106824 40228 106880 40230
rect 106904 40228 106960 40230
rect 105928 39738 105984 39740
rect 106008 39738 106064 39740
rect 106088 39738 106144 39740
rect 106168 39738 106224 39740
rect 105928 39686 105974 39738
rect 105974 39686 105984 39738
rect 106008 39686 106038 39738
rect 106038 39686 106050 39738
rect 106050 39686 106064 39738
rect 106088 39686 106102 39738
rect 106102 39686 106114 39738
rect 106114 39686 106144 39738
rect 106168 39686 106178 39738
rect 106178 39686 106224 39738
rect 105928 39684 105984 39686
rect 106008 39684 106064 39686
rect 106088 39684 106144 39686
rect 106168 39684 106224 39686
rect 106664 39194 106720 39196
rect 106744 39194 106800 39196
rect 106824 39194 106880 39196
rect 106904 39194 106960 39196
rect 106664 39142 106710 39194
rect 106710 39142 106720 39194
rect 106744 39142 106774 39194
rect 106774 39142 106786 39194
rect 106786 39142 106800 39194
rect 106824 39142 106838 39194
rect 106838 39142 106850 39194
rect 106850 39142 106880 39194
rect 106904 39142 106914 39194
rect 106914 39142 106960 39194
rect 106664 39140 106720 39142
rect 106744 39140 106800 39142
rect 106824 39140 106880 39142
rect 106904 39140 106960 39142
rect 105928 38650 105984 38652
rect 106008 38650 106064 38652
rect 106088 38650 106144 38652
rect 106168 38650 106224 38652
rect 105928 38598 105974 38650
rect 105974 38598 105984 38650
rect 106008 38598 106038 38650
rect 106038 38598 106050 38650
rect 106050 38598 106064 38650
rect 106088 38598 106102 38650
rect 106102 38598 106114 38650
rect 106114 38598 106144 38650
rect 106168 38598 106178 38650
rect 106178 38598 106224 38650
rect 105928 38596 105984 38598
rect 106008 38596 106064 38598
rect 106088 38596 106144 38598
rect 106168 38596 106224 38598
rect 106664 38106 106720 38108
rect 106744 38106 106800 38108
rect 106824 38106 106880 38108
rect 106904 38106 106960 38108
rect 106664 38054 106710 38106
rect 106710 38054 106720 38106
rect 106744 38054 106774 38106
rect 106774 38054 106786 38106
rect 106786 38054 106800 38106
rect 106824 38054 106838 38106
rect 106838 38054 106850 38106
rect 106850 38054 106880 38106
rect 106904 38054 106914 38106
rect 106914 38054 106960 38106
rect 106664 38052 106720 38054
rect 106744 38052 106800 38054
rect 106824 38052 106880 38054
rect 106904 38052 106960 38054
rect 105928 37562 105984 37564
rect 106008 37562 106064 37564
rect 106088 37562 106144 37564
rect 106168 37562 106224 37564
rect 105928 37510 105974 37562
rect 105974 37510 105984 37562
rect 106008 37510 106038 37562
rect 106038 37510 106050 37562
rect 106050 37510 106064 37562
rect 106088 37510 106102 37562
rect 106102 37510 106114 37562
rect 106114 37510 106144 37562
rect 106168 37510 106178 37562
rect 106178 37510 106224 37562
rect 105928 37508 105984 37510
rect 106008 37508 106064 37510
rect 106088 37508 106144 37510
rect 106168 37508 106224 37510
rect 106664 37018 106720 37020
rect 106744 37018 106800 37020
rect 106824 37018 106880 37020
rect 106904 37018 106960 37020
rect 106664 36966 106710 37018
rect 106710 36966 106720 37018
rect 106744 36966 106774 37018
rect 106774 36966 106786 37018
rect 106786 36966 106800 37018
rect 106824 36966 106838 37018
rect 106838 36966 106850 37018
rect 106850 36966 106880 37018
rect 106904 36966 106914 37018
rect 106914 36966 106960 37018
rect 106664 36964 106720 36966
rect 106744 36964 106800 36966
rect 106824 36964 106880 36966
rect 106904 36964 106960 36966
rect 105928 36474 105984 36476
rect 106008 36474 106064 36476
rect 106088 36474 106144 36476
rect 106168 36474 106224 36476
rect 105928 36422 105974 36474
rect 105974 36422 105984 36474
rect 106008 36422 106038 36474
rect 106038 36422 106050 36474
rect 106050 36422 106064 36474
rect 106088 36422 106102 36474
rect 106102 36422 106114 36474
rect 106114 36422 106144 36474
rect 106168 36422 106178 36474
rect 106178 36422 106224 36474
rect 105928 36420 105984 36422
rect 106008 36420 106064 36422
rect 106088 36420 106144 36422
rect 106168 36420 106224 36422
rect 106664 35930 106720 35932
rect 106744 35930 106800 35932
rect 106824 35930 106880 35932
rect 106904 35930 106960 35932
rect 106664 35878 106710 35930
rect 106710 35878 106720 35930
rect 106744 35878 106774 35930
rect 106774 35878 106786 35930
rect 106786 35878 106800 35930
rect 106824 35878 106838 35930
rect 106838 35878 106850 35930
rect 106850 35878 106880 35930
rect 106904 35878 106914 35930
rect 106914 35878 106960 35930
rect 106664 35876 106720 35878
rect 106744 35876 106800 35878
rect 106824 35876 106880 35878
rect 106904 35876 106960 35878
rect 105928 35386 105984 35388
rect 106008 35386 106064 35388
rect 106088 35386 106144 35388
rect 106168 35386 106224 35388
rect 105928 35334 105974 35386
rect 105974 35334 105984 35386
rect 106008 35334 106038 35386
rect 106038 35334 106050 35386
rect 106050 35334 106064 35386
rect 106088 35334 106102 35386
rect 106102 35334 106114 35386
rect 106114 35334 106144 35386
rect 106168 35334 106178 35386
rect 106178 35334 106224 35386
rect 105928 35332 105984 35334
rect 106008 35332 106064 35334
rect 106088 35332 106144 35334
rect 106168 35332 106224 35334
rect 106664 34842 106720 34844
rect 106744 34842 106800 34844
rect 106824 34842 106880 34844
rect 106904 34842 106960 34844
rect 106664 34790 106710 34842
rect 106710 34790 106720 34842
rect 106744 34790 106774 34842
rect 106774 34790 106786 34842
rect 106786 34790 106800 34842
rect 106824 34790 106838 34842
rect 106838 34790 106850 34842
rect 106850 34790 106880 34842
rect 106904 34790 106914 34842
rect 106914 34790 106960 34842
rect 106664 34788 106720 34790
rect 106744 34788 106800 34790
rect 106824 34788 106880 34790
rect 106904 34788 106960 34790
rect 105928 34298 105984 34300
rect 106008 34298 106064 34300
rect 106088 34298 106144 34300
rect 106168 34298 106224 34300
rect 105928 34246 105974 34298
rect 105974 34246 105984 34298
rect 106008 34246 106038 34298
rect 106038 34246 106050 34298
rect 106050 34246 106064 34298
rect 106088 34246 106102 34298
rect 106102 34246 106114 34298
rect 106114 34246 106144 34298
rect 106168 34246 106178 34298
rect 106178 34246 106224 34298
rect 105928 34244 105984 34246
rect 106008 34244 106064 34246
rect 106088 34244 106144 34246
rect 106168 34244 106224 34246
rect 106664 33754 106720 33756
rect 106744 33754 106800 33756
rect 106824 33754 106880 33756
rect 106904 33754 106960 33756
rect 106664 33702 106710 33754
rect 106710 33702 106720 33754
rect 106744 33702 106774 33754
rect 106774 33702 106786 33754
rect 106786 33702 106800 33754
rect 106824 33702 106838 33754
rect 106838 33702 106850 33754
rect 106850 33702 106880 33754
rect 106904 33702 106914 33754
rect 106914 33702 106960 33754
rect 106664 33700 106720 33702
rect 106744 33700 106800 33702
rect 106824 33700 106880 33702
rect 106904 33700 106960 33702
rect 105928 33210 105984 33212
rect 106008 33210 106064 33212
rect 106088 33210 106144 33212
rect 106168 33210 106224 33212
rect 105928 33158 105974 33210
rect 105974 33158 105984 33210
rect 106008 33158 106038 33210
rect 106038 33158 106050 33210
rect 106050 33158 106064 33210
rect 106088 33158 106102 33210
rect 106102 33158 106114 33210
rect 106114 33158 106144 33210
rect 106168 33158 106178 33210
rect 106178 33158 106224 33210
rect 105928 33156 105984 33158
rect 106008 33156 106064 33158
rect 106088 33156 106144 33158
rect 106168 33156 106224 33158
rect 106664 32666 106720 32668
rect 106744 32666 106800 32668
rect 106824 32666 106880 32668
rect 106904 32666 106960 32668
rect 106664 32614 106710 32666
rect 106710 32614 106720 32666
rect 106744 32614 106774 32666
rect 106774 32614 106786 32666
rect 106786 32614 106800 32666
rect 106824 32614 106838 32666
rect 106838 32614 106850 32666
rect 106850 32614 106880 32666
rect 106904 32614 106914 32666
rect 106914 32614 106960 32666
rect 106664 32612 106720 32614
rect 106744 32612 106800 32614
rect 106824 32612 106880 32614
rect 106904 32612 106960 32614
rect 105928 32122 105984 32124
rect 106008 32122 106064 32124
rect 106088 32122 106144 32124
rect 106168 32122 106224 32124
rect 105928 32070 105974 32122
rect 105974 32070 105984 32122
rect 106008 32070 106038 32122
rect 106038 32070 106050 32122
rect 106050 32070 106064 32122
rect 106088 32070 106102 32122
rect 106102 32070 106114 32122
rect 106114 32070 106144 32122
rect 106168 32070 106178 32122
rect 106178 32070 106224 32122
rect 105928 32068 105984 32070
rect 106008 32068 106064 32070
rect 106088 32068 106144 32070
rect 106168 32068 106224 32070
rect 106664 31578 106720 31580
rect 106744 31578 106800 31580
rect 106824 31578 106880 31580
rect 106904 31578 106960 31580
rect 106664 31526 106710 31578
rect 106710 31526 106720 31578
rect 106744 31526 106774 31578
rect 106774 31526 106786 31578
rect 106786 31526 106800 31578
rect 106824 31526 106838 31578
rect 106838 31526 106850 31578
rect 106850 31526 106880 31578
rect 106904 31526 106914 31578
rect 106914 31526 106960 31578
rect 106664 31524 106720 31526
rect 106744 31524 106800 31526
rect 106824 31524 106880 31526
rect 106904 31524 106960 31526
rect 105928 31034 105984 31036
rect 106008 31034 106064 31036
rect 106088 31034 106144 31036
rect 106168 31034 106224 31036
rect 105928 30982 105974 31034
rect 105974 30982 105984 31034
rect 106008 30982 106038 31034
rect 106038 30982 106050 31034
rect 106050 30982 106064 31034
rect 106088 30982 106102 31034
rect 106102 30982 106114 31034
rect 106114 30982 106144 31034
rect 106168 30982 106178 31034
rect 106178 30982 106224 31034
rect 105928 30980 105984 30982
rect 106008 30980 106064 30982
rect 106088 30980 106144 30982
rect 106168 30980 106224 30982
rect 106664 30490 106720 30492
rect 106744 30490 106800 30492
rect 106824 30490 106880 30492
rect 106904 30490 106960 30492
rect 106664 30438 106710 30490
rect 106710 30438 106720 30490
rect 106744 30438 106774 30490
rect 106774 30438 106786 30490
rect 106786 30438 106800 30490
rect 106824 30438 106838 30490
rect 106838 30438 106850 30490
rect 106850 30438 106880 30490
rect 106904 30438 106914 30490
rect 106914 30438 106960 30490
rect 106664 30436 106720 30438
rect 106744 30436 106800 30438
rect 106824 30436 106880 30438
rect 106904 30436 106960 30438
rect 105928 29946 105984 29948
rect 106008 29946 106064 29948
rect 106088 29946 106144 29948
rect 106168 29946 106224 29948
rect 105928 29894 105974 29946
rect 105974 29894 105984 29946
rect 106008 29894 106038 29946
rect 106038 29894 106050 29946
rect 106050 29894 106064 29946
rect 106088 29894 106102 29946
rect 106102 29894 106114 29946
rect 106114 29894 106144 29946
rect 106168 29894 106178 29946
rect 106178 29894 106224 29946
rect 105928 29892 105984 29894
rect 106008 29892 106064 29894
rect 106088 29892 106144 29894
rect 106168 29892 106224 29894
rect 106664 29402 106720 29404
rect 106744 29402 106800 29404
rect 106824 29402 106880 29404
rect 106904 29402 106960 29404
rect 106664 29350 106710 29402
rect 106710 29350 106720 29402
rect 106744 29350 106774 29402
rect 106774 29350 106786 29402
rect 106786 29350 106800 29402
rect 106824 29350 106838 29402
rect 106838 29350 106850 29402
rect 106850 29350 106880 29402
rect 106904 29350 106914 29402
rect 106914 29350 106960 29402
rect 106664 29348 106720 29350
rect 106744 29348 106800 29350
rect 106824 29348 106880 29350
rect 106904 29348 106960 29350
rect 105928 28858 105984 28860
rect 106008 28858 106064 28860
rect 106088 28858 106144 28860
rect 106168 28858 106224 28860
rect 105928 28806 105974 28858
rect 105974 28806 105984 28858
rect 106008 28806 106038 28858
rect 106038 28806 106050 28858
rect 106050 28806 106064 28858
rect 106088 28806 106102 28858
rect 106102 28806 106114 28858
rect 106114 28806 106144 28858
rect 106168 28806 106178 28858
rect 106178 28806 106224 28858
rect 105928 28804 105984 28806
rect 106008 28804 106064 28806
rect 106088 28804 106144 28806
rect 106168 28804 106224 28806
rect 106664 28314 106720 28316
rect 106744 28314 106800 28316
rect 106824 28314 106880 28316
rect 106904 28314 106960 28316
rect 106664 28262 106710 28314
rect 106710 28262 106720 28314
rect 106744 28262 106774 28314
rect 106774 28262 106786 28314
rect 106786 28262 106800 28314
rect 106824 28262 106838 28314
rect 106838 28262 106850 28314
rect 106850 28262 106880 28314
rect 106904 28262 106914 28314
rect 106914 28262 106960 28314
rect 106664 28260 106720 28262
rect 106744 28260 106800 28262
rect 106824 28260 106880 28262
rect 106904 28260 106960 28262
rect 105928 27770 105984 27772
rect 106008 27770 106064 27772
rect 106088 27770 106144 27772
rect 106168 27770 106224 27772
rect 105928 27718 105974 27770
rect 105974 27718 105984 27770
rect 106008 27718 106038 27770
rect 106038 27718 106050 27770
rect 106050 27718 106064 27770
rect 106088 27718 106102 27770
rect 106102 27718 106114 27770
rect 106114 27718 106144 27770
rect 106168 27718 106178 27770
rect 106178 27718 106224 27770
rect 105928 27716 105984 27718
rect 106008 27716 106064 27718
rect 106088 27716 106144 27718
rect 106168 27716 106224 27718
rect 106664 27226 106720 27228
rect 106744 27226 106800 27228
rect 106824 27226 106880 27228
rect 106904 27226 106960 27228
rect 106664 27174 106710 27226
rect 106710 27174 106720 27226
rect 106744 27174 106774 27226
rect 106774 27174 106786 27226
rect 106786 27174 106800 27226
rect 106824 27174 106838 27226
rect 106838 27174 106850 27226
rect 106850 27174 106880 27226
rect 106904 27174 106914 27226
rect 106914 27174 106960 27226
rect 106664 27172 106720 27174
rect 106744 27172 106800 27174
rect 106824 27172 106880 27174
rect 106904 27172 106960 27174
rect 105928 26682 105984 26684
rect 106008 26682 106064 26684
rect 106088 26682 106144 26684
rect 106168 26682 106224 26684
rect 105928 26630 105974 26682
rect 105974 26630 105984 26682
rect 106008 26630 106038 26682
rect 106038 26630 106050 26682
rect 106050 26630 106064 26682
rect 106088 26630 106102 26682
rect 106102 26630 106114 26682
rect 106114 26630 106144 26682
rect 106168 26630 106178 26682
rect 106178 26630 106224 26682
rect 105928 26628 105984 26630
rect 106008 26628 106064 26630
rect 106088 26628 106144 26630
rect 106168 26628 106224 26630
rect 106664 26138 106720 26140
rect 106744 26138 106800 26140
rect 106824 26138 106880 26140
rect 106904 26138 106960 26140
rect 106664 26086 106710 26138
rect 106710 26086 106720 26138
rect 106744 26086 106774 26138
rect 106774 26086 106786 26138
rect 106786 26086 106800 26138
rect 106824 26086 106838 26138
rect 106838 26086 106850 26138
rect 106850 26086 106880 26138
rect 106904 26086 106914 26138
rect 106914 26086 106960 26138
rect 106664 26084 106720 26086
rect 106744 26084 106800 26086
rect 106824 26084 106880 26086
rect 106904 26084 106960 26086
rect 105928 25594 105984 25596
rect 106008 25594 106064 25596
rect 106088 25594 106144 25596
rect 106168 25594 106224 25596
rect 105928 25542 105974 25594
rect 105974 25542 105984 25594
rect 106008 25542 106038 25594
rect 106038 25542 106050 25594
rect 106050 25542 106064 25594
rect 106088 25542 106102 25594
rect 106102 25542 106114 25594
rect 106114 25542 106144 25594
rect 106168 25542 106178 25594
rect 106178 25542 106224 25594
rect 105928 25540 105984 25542
rect 106008 25540 106064 25542
rect 106088 25540 106144 25542
rect 106168 25540 106224 25542
rect 106664 25050 106720 25052
rect 106744 25050 106800 25052
rect 106824 25050 106880 25052
rect 106904 25050 106960 25052
rect 106664 24998 106710 25050
rect 106710 24998 106720 25050
rect 106744 24998 106774 25050
rect 106774 24998 106786 25050
rect 106786 24998 106800 25050
rect 106824 24998 106838 25050
rect 106838 24998 106850 25050
rect 106850 24998 106880 25050
rect 106904 24998 106914 25050
rect 106914 24998 106960 25050
rect 106664 24996 106720 24998
rect 106744 24996 106800 24998
rect 106824 24996 106880 24998
rect 106904 24996 106960 24998
rect 105928 24506 105984 24508
rect 106008 24506 106064 24508
rect 106088 24506 106144 24508
rect 106168 24506 106224 24508
rect 105928 24454 105974 24506
rect 105974 24454 105984 24506
rect 106008 24454 106038 24506
rect 106038 24454 106050 24506
rect 106050 24454 106064 24506
rect 106088 24454 106102 24506
rect 106102 24454 106114 24506
rect 106114 24454 106144 24506
rect 106168 24454 106178 24506
rect 106178 24454 106224 24506
rect 105928 24452 105984 24454
rect 106008 24452 106064 24454
rect 106088 24452 106144 24454
rect 106168 24452 106224 24454
rect 106664 23962 106720 23964
rect 106744 23962 106800 23964
rect 106824 23962 106880 23964
rect 106904 23962 106960 23964
rect 106664 23910 106710 23962
rect 106710 23910 106720 23962
rect 106744 23910 106774 23962
rect 106774 23910 106786 23962
rect 106786 23910 106800 23962
rect 106824 23910 106838 23962
rect 106838 23910 106850 23962
rect 106850 23910 106880 23962
rect 106904 23910 106914 23962
rect 106914 23910 106960 23962
rect 106664 23908 106720 23910
rect 106744 23908 106800 23910
rect 106824 23908 106880 23910
rect 106904 23908 106960 23910
rect 105928 23418 105984 23420
rect 106008 23418 106064 23420
rect 106088 23418 106144 23420
rect 106168 23418 106224 23420
rect 105928 23366 105974 23418
rect 105974 23366 105984 23418
rect 106008 23366 106038 23418
rect 106038 23366 106050 23418
rect 106050 23366 106064 23418
rect 106088 23366 106102 23418
rect 106102 23366 106114 23418
rect 106114 23366 106144 23418
rect 106168 23366 106178 23418
rect 106178 23366 106224 23418
rect 105928 23364 105984 23366
rect 106008 23364 106064 23366
rect 106088 23364 106144 23366
rect 106168 23364 106224 23366
rect 106664 22874 106720 22876
rect 106744 22874 106800 22876
rect 106824 22874 106880 22876
rect 106904 22874 106960 22876
rect 106664 22822 106710 22874
rect 106710 22822 106720 22874
rect 106744 22822 106774 22874
rect 106774 22822 106786 22874
rect 106786 22822 106800 22874
rect 106824 22822 106838 22874
rect 106838 22822 106850 22874
rect 106850 22822 106880 22874
rect 106904 22822 106914 22874
rect 106914 22822 106960 22874
rect 106664 22820 106720 22822
rect 106744 22820 106800 22822
rect 106824 22820 106880 22822
rect 106904 22820 106960 22822
rect 105928 22330 105984 22332
rect 106008 22330 106064 22332
rect 106088 22330 106144 22332
rect 106168 22330 106224 22332
rect 105928 22278 105974 22330
rect 105974 22278 105984 22330
rect 106008 22278 106038 22330
rect 106038 22278 106050 22330
rect 106050 22278 106064 22330
rect 106088 22278 106102 22330
rect 106102 22278 106114 22330
rect 106114 22278 106144 22330
rect 106168 22278 106178 22330
rect 106178 22278 106224 22330
rect 105928 22276 105984 22278
rect 106008 22276 106064 22278
rect 106088 22276 106144 22278
rect 106168 22276 106224 22278
rect 106664 21786 106720 21788
rect 106744 21786 106800 21788
rect 106824 21786 106880 21788
rect 106904 21786 106960 21788
rect 106664 21734 106710 21786
rect 106710 21734 106720 21786
rect 106744 21734 106774 21786
rect 106774 21734 106786 21786
rect 106786 21734 106800 21786
rect 106824 21734 106838 21786
rect 106838 21734 106850 21786
rect 106850 21734 106880 21786
rect 106904 21734 106914 21786
rect 106914 21734 106960 21786
rect 106664 21732 106720 21734
rect 106744 21732 106800 21734
rect 106824 21732 106880 21734
rect 106904 21732 106960 21734
rect 105928 21242 105984 21244
rect 106008 21242 106064 21244
rect 106088 21242 106144 21244
rect 106168 21242 106224 21244
rect 105928 21190 105974 21242
rect 105974 21190 105984 21242
rect 106008 21190 106038 21242
rect 106038 21190 106050 21242
rect 106050 21190 106064 21242
rect 106088 21190 106102 21242
rect 106102 21190 106114 21242
rect 106114 21190 106144 21242
rect 106168 21190 106178 21242
rect 106178 21190 106224 21242
rect 105928 21188 105984 21190
rect 106008 21188 106064 21190
rect 106088 21188 106144 21190
rect 106168 21188 106224 21190
rect 106664 20698 106720 20700
rect 106744 20698 106800 20700
rect 106824 20698 106880 20700
rect 106904 20698 106960 20700
rect 106664 20646 106710 20698
rect 106710 20646 106720 20698
rect 106744 20646 106774 20698
rect 106774 20646 106786 20698
rect 106786 20646 106800 20698
rect 106824 20646 106838 20698
rect 106838 20646 106850 20698
rect 106850 20646 106880 20698
rect 106904 20646 106914 20698
rect 106914 20646 106960 20698
rect 106664 20644 106720 20646
rect 106744 20644 106800 20646
rect 106824 20644 106880 20646
rect 106904 20644 106960 20646
rect 105928 20154 105984 20156
rect 106008 20154 106064 20156
rect 106088 20154 106144 20156
rect 106168 20154 106224 20156
rect 105928 20102 105974 20154
rect 105974 20102 105984 20154
rect 106008 20102 106038 20154
rect 106038 20102 106050 20154
rect 106050 20102 106064 20154
rect 106088 20102 106102 20154
rect 106102 20102 106114 20154
rect 106114 20102 106144 20154
rect 106168 20102 106178 20154
rect 106178 20102 106224 20154
rect 105928 20100 105984 20102
rect 106008 20100 106064 20102
rect 106088 20100 106144 20102
rect 106168 20100 106224 20102
rect 106664 19610 106720 19612
rect 106744 19610 106800 19612
rect 106824 19610 106880 19612
rect 106904 19610 106960 19612
rect 106664 19558 106710 19610
rect 106710 19558 106720 19610
rect 106744 19558 106774 19610
rect 106774 19558 106786 19610
rect 106786 19558 106800 19610
rect 106824 19558 106838 19610
rect 106838 19558 106850 19610
rect 106850 19558 106880 19610
rect 106904 19558 106914 19610
rect 106914 19558 106960 19610
rect 106664 19556 106720 19558
rect 106744 19556 106800 19558
rect 106824 19556 106880 19558
rect 106904 19556 106960 19558
rect 105928 19066 105984 19068
rect 106008 19066 106064 19068
rect 106088 19066 106144 19068
rect 106168 19066 106224 19068
rect 105928 19014 105974 19066
rect 105974 19014 105984 19066
rect 106008 19014 106038 19066
rect 106038 19014 106050 19066
rect 106050 19014 106064 19066
rect 106088 19014 106102 19066
rect 106102 19014 106114 19066
rect 106114 19014 106144 19066
rect 106168 19014 106178 19066
rect 106178 19014 106224 19066
rect 105928 19012 105984 19014
rect 106008 19012 106064 19014
rect 106088 19012 106144 19014
rect 106168 19012 106224 19014
rect 106664 18522 106720 18524
rect 106744 18522 106800 18524
rect 106824 18522 106880 18524
rect 106904 18522 106960 18524
rect 106664 18470 106710 18522
rect 106710 18470 106720 18522
rect 106744 18470 106774 18522
rect 106774 18470 106786 18522
rect 106786 18470 106800 18522
rect 106824 18470 106838 18522
rect 106838 18470 106850 18522
rect 106850 18470 106880 18522
rect 106904 18470 106914 18522
rect 106914 18470 106960 18522
rect 106664 18468 106720 18470
rect 106744 18468 106800 18470
rect 106824 18468 106880 18470
rect 106904 18468 106960 18470
rect 105928 17978 105984 17980
rect 106008 17978 106064 17980
rect 106088 17978 106144 17980
rect 106168 17978 106224 17980
rect 105928 17926 105974 17978
rect 105974 17926 105984 17978
rect 106008 17926 106038 17978
rect 106038 17926 106050 17978
rect 106050 17926 106064 17978
rect 106088 17926 106102 17978
rect 106102 17926 106114 17978
rect 106114 17926 106144 17978
rect 106168 17926 106178 17978
rect 106178 17926 106224 17978
rect 105928 17924 105984 17926
rect 106008 17924 106064 17926
rect 106088 17924 106144 17926
rect 106168 17924 106224 17926
rect 106664 17434 106720 17436
rect 106744 17434 106800 17436
rect 106824 17434 106880 17436
rect 106904 17434 106960 17436
rect 106664 17382 106710 17434
rect 106710 17382 106720 17434
rect 106744 17382 106774 17434
rect 106774 17382 106786 17434
rect 106786 17382 106800 17434
rect 106824 17382 106838 17434
rect 106838 17382 106850 17434
rect 106850 17382 106880 17434
rect 106904 17382 106914 17434
rect 106914 17382 106960 17434
rect 106664 17380 106720 17382
rect 106744 17380 106800 17382
rect 106824 17380 106880 17382
rect 106904 17380 106960 17382
rect 105928 16890 105984 16892
rect 106008 16890 106064 16892
rect 106088 16890 106144 16892
rect 106168 16890 106224 16892
rect 105928 16838 105974 16890
rect 105974 16838 105984 16890
rect 106008 16838 106038 16890
rect 106038 16838 106050 16890
rect 106050 16838 106064 16890
rect 106088 16838 106102 16890
rect 106102 16838 106114 16890
rect 106114 16838 106144 16890
rect 106168 16838 106178 16890
rect 106178 16838 106224 16890
rect 105928 16836 105984 16838
rect 106008 16836 106064 16838
rect 106088 16836 106144 16838
rect 106168 16836 106224 16838
rect 106664 16346 106720 16348
rect 106744 16346 106800 16348
rect 106824 16346 106880 16348
rect 106904 16346 106960 16348
rect 106664 16294 106710 16346
rect 106710 16294 106720 16346
rect 106744 16294 106774 16346
rect 106774 16294 106786 16346
rect 106786 16294 106800 16346
rect 106824 16294 106838 16346
rect 106838 16294 106850 16346
rect 106850 16294 106880 16346
rect 106904 16294 106914 16346
rect 106914 16294 106960 16346
rect 106664 16292 106720 16294
rect 106744 16292 106800 16294
rect 106824 16292 106880 16294
rect 106904 16292 106960 16294
rect 105928 15802 105984 15804
rect 106008 15802 106064 15804
rect 106088 15802 106144 15804
rect 106168 15802 106224 15804
rect 105928 15750 105974 15802
rect 105974 15750 105984 15802
rect 106008 15750 106038 15802
rect 106038 15750 106050 15802
rect 106050 15750 106064 15802
rect 106088 15750 106102 15802
rect 106102 15750 106114 15802
rect 106114 15750 106144 15802
rect 106168 15750 106178 15802
rect 106178 15750 106224 15802
rect 105928 15748 105984 15750
rect 106008 15748 106064 15750
rect 106088 15748 106144 15750
rect 106168 15748 106224 15750
rect 106664 15258 106720 15260
rect 106744 15258 106800 15260
rect 106824 15258 106880 15260
rect 106904 15258 106960 15260
rect 106664 15206 106710 15258
rect 106710 15206 106720 15258
rect 106744 15206 106774 15258
rect 106774 15206 106786 15258
rect 106786 15206 106800 15258
rect 106824 15206 106838 15258
rect 106838 15206 106850 15258
rect 106850 15206 106880 15258
rect 106904 15206 106914 15258
rect 106914 15206 106960 15258
rect 106664 15204 106720 15206
rect 106744 15204 106800 15206
rect 106824 15204 106880 15206
rect 106904 15204 106960 15206
rect 105928 14714 105984 14716
rect 106008 14714 106064 14716
rect 106088 14714 106144 14716
rect 106168 14714 106224 14716
rect 105928 14662 105974 14714
rect 105974 14662 105984 14714
rect 106008 14662 106038 14714
rect 106038 14662 106050 14714
rect 106050 14662 106064 14714
rect 106088 14662 106102 14714
rect 106102 14662 106114 14714
rect 106114 14662 106144 14714
rect 106168 14662 106178 14714
rect 106178 14662 106224 14714
rect 105928 14660 105984 14662
rect 106008 14660 106064 14662
rect 106088 14660 106144 14662
rect 106168 14660 106224 14662
rect 106664 14170 106720 14172
rect 106744 14170 106800 14172
rect 106824 14170 106880 14172
rect 106904 14170 106960 14172
rect 106664 14118 106710 14170
rect 106710 14118 106720 14170
rect 106744 14118 106774 14170
rect 106774 14118 106786 14170
rect 106786 14118 106800 14170
rect 106824 14118 106838 14170
rect 106838 14118 106850 14170
rect 106850 14118 106880 14170
rect 106904 14118 106914 14170
rect 106914 14118 106960 14170
rect 106664 14116 106720 14118
rect 106744 14116 106800 14118
rect 106824 14116 106880 14118
rect 106904 14116 106960 14118
rect 105928 13626 105984 13628
rect 106008 13626 106064 13628
rect 106088 13626 106144 13628
rect 106168 13626 106224 13628
rect 105928 13574 105974 13626
rect 105974 13574 105984 13626
rect 106008 13574 106038 13626
rect 106038 13574 106050 13626
rect 106050 13574 106064 13626
rect 106088 13574 106102 13626
rect 106102 13574 106114 13626
rect 106114 13574 106144 13626
rect 106168 13574 106178 13626
rect 106178 13574 106224 13626
rect 105928 13572 105984 13574
rect 106008 13572 106064 13574
rect 106088 13572 106144 13574
rect 106168 13572 106224 13574
rect 106664 13082 106720 13084
rect 106744 13082 106800 13084
rect 106824 13082 106880 13084
rect 106904 13082 106960 13084
rect 106664 13030 106710 13082
rect 106710 13030 106720 13082
rect 106744 13030 106774 13082
rect 106774 13030 106786 13082
rect 106786 13030 106800 13082
rect 106824 13030 106838 13082
rect 106838 13030 106850 13082
rect 106850 13030 106880 13082
rect 106904 13030 106914 13082
rect 106914 13030 106960 13082
rect 106664 13028 106720 13030
rect 106744 13028 106800 13030
rect 106824 13028 106880 13030
rect 106904 13028 106960 13030
rect 105928 12538 105984 12540
rect 106008 12538 106064 12540
rect 106088 12538 106144 12540
rect 106168 12538 106224 12540
rect 105928 12486 105974 12538
rect 105974 12486 105984 12538
rect 106008 12486 106038 12538
rect 106038 12486 106050 12538
rect 106050 12486 106064 12538
rect 106088 12486 106102 12538
rect 106102 12486 106114 12538
rect 106114 12486 106144 12538
rect 106168 12486 106178 12538
rect 106178 12486 106224 12538
rect 105928 12484 105984 12486
rect 106008 12484 106064 12486
rect 106088 12484 106144 12486
rect 106168 12484 106224 12486
rect 106664 11994 106720 11996
rect 106744 11994 106800 11996
rect 106824 11994 106880 11996
rect 106904 11994 106960 11996
rect 106664 11942 106710 11994
rect 106710 11942 106720 11994
rect 106744 11942 106774 11994
rect 106774 11942 106786 11994
rect 106786 11942 106800 11994
rect 106824 11942 106838 11994
rect 106838 11942 106850 11994
rect 106850 11942 106880 11994
rect 106904 11942 106914 11994
rect 106914 11942 106960 11994
rect 106664 11940 106720 11942
rect 106744 11940 106800 11942
rect 106824 11940 106880 11942
rect 106904 11940 106960 11942
rect 105928 11450 105984 11452
rect 106008 11450 106064 11452
rect 106088 11450 106144 11452
rect 106168 11450 106224 11452
rect 105928 11398 105974 11450
rect 105974 11398 105984 11450
rect 106008 11398 106038 11450
rect 106038 11398 106050 11450
rect 106050 11398 106064 11450
rect 106088 11398 106102 11450
rect 106102 11398 106114 11450
rect 106114 11398 106144 11450
rect 106168 11398 106178 11450
rect 106178 11398 106224 11450
rect 105928 11396 105984 11398
rect 106008 11396 106064 11398
rect 106088 11396 106144 11398
rect 106168 11396 106224 11398
rect 106664 10906 106720 10908
rect 106744 10906 106800 10908
rect 106824 10906 106880 10908
rect 106904 10906 106960 10908
rect 106664 10854 106710 10906
rect 106710 10854 106720 10906
rect 106744 10854 106774 10906
rect 106774 10854 106786 10906
rect 106786 10854 106800 10906
rect 106824 10854 106838 10906
rect 106838 10854 106850 10906
rect 106850 10854 106880 10906
rect 106904 10854 106914 10906
rect 106914 10854 106960 10906
rect 106664 10852 106720 10854
rect 106744 10852 106800 10854
rect 106824 10852 106880 10854
rect 106904 10852 106960 10854
rect 105928 10362 105984 10364
rect 106008 10362 106064 10364
rect 106088 10362 106144 10364
rect 106168 10362 106224 10364
rect 105928 10310 105974 10362
rect 105974 10310 105984 10362
rect 106008 10310 106038 10362
rect 106038 10310 106050 10362
rect 106050 10310 106064 10362
rect 106088 10310 106102 10362
rect 106102 10310 106114 10362
rect 106114 10310 106144 10362
rect 106168 10310 106178 10362
rect 106178 10310 106224 10362
rect 105928 10308 105984 10310
rect 106008 10308 106064 10310
rect 106088 10308 106144 10310
rect 106168 10308 106224 10310
rect 90822 9832 90878 9888
rect 104806 9832 104862 9888
rect 106664 9818 106720 9820
rect 106744 9818 106800 9820
rect 106824 9818 106880 9820
rect 106904 9818 106960 9820
rect 106664 9766 106710 9818
rect 106710 9766 106720 9818
rect 106744 9766 106774 9818
rect 106774 9766 106786 9818
rect 106786 9766 106800 9818
rect 106824 9766 106838 9818
rect 106838 9766 106850 9818
rect 106850 9766 106880 9818
rect 106904 9766 106914 9818
rect 106914 9766 106960 9818
rect 106664 9764 106720 9766
rect 106744 9764 106800 9766
rect 106824 9764 106880 9766
rect 106904 9764 106960 9766
rect 90730 9696 90786 9752
rect 23478 8200 23534 8256
rect 24766 8200 24822 8256
rect 25870 8200 25926 8256
rect 27158 8200 27214 8256
rect 28446 8200 28502 8256
rect 29274 8200 29330 8256
rect 30562 8200 30618 8256
rect 31666 8200 31722 8256
rect 32954 8200 33010 8256
rect 34242 8200 34298 8256
rect 35438 8200 35494 8256
rect 36358 8200 36414 8256
rect 37462 8200 37518 8256
rect 38750 8200 38806 8256
rect 41326 8200 41382 8256
rect 42154 8200 42210 8256
rect 43442 8200 43498 8256
rect 90638 8200 90694 8256
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 39946 4528 40002 4584
rect 66320 7642 66376 7644
rect 66400 7642 66456 7644
rect 66480 7642 66536 7644
rect 66560 7642 66616 7644
rect 66320 7590 66366 7642
rect 66366 7590 66376 7642
rect 66400 7590 66430 7642
rect 66430 7590 66442 7642
rect 66442 7590 66456 7642
rect 66480 7590 66494 7642
rect 66494 7590 66506 7642
rect 66506 7590 66536 7642
rect 66560 7590 66570 7642
rect 66570 7590 66616 7642
rect 66320 7588 66376 7590
rect 66400 7588 66456 7590
rect 66480 7588 66536 7590
rect 66560 7588 66616 7590
rect 105928 9274 105984 9276
rect 106008 9274 106064 9276
rect 106088 9274 106144 9276
rect 106168 9274 106224 9276
rect 105928 9222 105974 9274
rect 105974 9222 105984 9274
rect 106008 9222 106038 9274
rect 106038 9222 106050 9274
rect 106050 9222 106064 9274
rect 106088 9222 106102 9274
rect 106102 9222 106114 9274
rect 106114 9222 106144 9274
rect 106168 9222 106178 9274
rect 106178 9222 106224 9274
rect 105928 9220 105984 9222
rect 106008 9220 106064 9222
rect 106088 9220 106144 9222
rect 106168 9220 106224 9222
rect 106664 8730 106720 8732
rect 106744 8730 106800 8732
rect 106824 8730 106880 8732
rect 106904 8730 106960 8732
rect 106664 8678 106710 8730
rect 106710 8678 106720 8730
rect 106744 8678 106774 8730
rect 106774 8678 106786 8730
rect 106786 8678 106800 8730
rect 106824 8678 106838 8730
rect 106838 8678 106850 8730
rect 106850 8678 106880 8730
rect 106904 8678 106914 8730
rect 106914 8678 106960 8730
rect 106664 8676 106720 8678
rect 106744 8676 106800 8678
rect 106824 8676 106880 8678
rect 106904 8676 106960 8678
rect 91006 8200 91062 8256
rect 105928 8186 105984 8188
rect 106008 8186 106064 8188
rect 106088 8186 106144 8188
rect 106168 8186 106224 8188
rect 105928 8134 105974 8186
rect 105974 8134 105984 8186
rect 106008 8134 106038 8186
rect 106038 8134 106050 8186
rect 106050 8134 106064 8186
rect 106088 8134 106102 8186
rect 106102 8134 106114 8186
rect 106114 8134 106144 8186
rect 106168 8134 106178 8186
rect 106178 8134 106224 8186
rect 105928 8132 105984 8134
rect 106008 8132 106064 8134
rect 106088 8132 106144 8134
rect 106168 8132 106224 8134
rect 97040 7642 97096 7644
rect 97120 7642 97176 7644
rect 97200 7642 97256 7644
rect 97280 7642 97336 7644
rect 97040 7590 97086 7642
rect 97086 7590 97096 7642
rect 97120 7590 97150 7642
rect 97150 7590 97162 7642
rect 97162 7590 97176 7642
rect 97200 7590 97214 7642
rect 97214 7590 97226 7642
rect 97226 7590 97256 7642
rect 97280 7590 97290 7642
rect 97290 7590 97336 7642
rect 97040 7588 97096 7590
rect 97120 7588 97176 7590
rect 97200 7588 97256 7590
rect 97280 7588 97336 7590
rect 106664 7642 106720 7644
rect 106744 7642 106800 7644
rect 106824 7642 106880 7644
rect 106904 7642 106960 7644
rect 106664 7590 106710 7642
rect 106710 7590 106720 7642
rect 106744 7590 106774 7642
rect 106774 7590 106786 7642
rect 106786 7590 106800 7642
rect 106824 7590 106838 7642
rect 106838 7590 106850 7642
rect 106850 7590 106880 7642
rect 106904 7590 106914 7642
rect 106914 7590 106960 7642
rect 106664 7588 106720 7590
rect 106744 7588 106800 7590
rect 106824 7588 106880 7590
rect 106904 7588 106960 7590
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 96380 7098 96436 7100
rect 96460 7098 96516 7100
rect 96540 7098 96596 7100
rect 96620 7098 96676 7100
rect 96380 7046 96426 7098
rect 96426 7046 96436 7098
rect 96460 7046 96490 7098
rect 96490 7046 96502 7098
rect 96502 7046 96516 7098
rect 96540 7046 96554 7098
rect 96554 7046 96566 7098
rect 96566 7046 96596 7098
rect 96620 7046 96630 7098
rect 96630 7046 96676 7098
rect 96380 7044 96436 7046
rect 96460 7044 96516 7046
rect 96540 7044 96596 7046
rect 96620 7044 96676 7046
rect 105928 7098 105984 7100
rect 106008 7098 106064 7100
rect 106088 7098 106144 7100
rect 106168 7098 106224 7100
rect 105928 7046 105974 7098
rect 105974 7046 105984 7098
rect 106008 7046 106038 7098
rect 106038 7046 106050 7098
rect 106050 7046 106064 7098
rect 106088 7046 106102 7098
rect 106102 7046 106114 7098
rect 106114 7046 106144 7098
rect 106168 7046 106178 7098
rect 106178 7046 106224 7098
rect 105928 7044 105984 7046
rect 106008 7044 106064 7046
rect 106088 7044 106144 7046
rect 106168 7044 106224 7046
rect 66320 6554 66376 6556
rect 66400 6554 66456 6556
rect 66480 6554 66536 6556
rect 66560 6554 66616 6556
rect 66320 6502 66366 6554
rect 66366 6502 66376 6554
rect 66400 6502 66430 6554
rect 66430 6502 66442 6554
rect 66442 6502 66456 6554
rect 66480 6502 66494 6554
rect 66494 6502 66506 6554
rect 66506 6502 66536 6554
rect 66560 6502 66570 6554
rect 66570 6502 66616 6554
rect 66320 6500 66376 6502
rect 66400 6500 66456 6502
rect 66480 6500 66536 6502
rect 66560 6500 66616 6502
rect 97040 6554 97096 6556
rect 97120 6554 97176 6556
rect 97200 6554 97256 6556
rect 97280 6554 97336 6556
rect 97040 6502 97086 6554
rect 97086 6502 97096 6554
rect 97120 6502 97150 6554
rect 97150 6502 97162 6554
rect 97162 6502 97176 6554
rect 97200 6502 97214 6554
rect 97214 6502 97226 6554
rect 97226 6502 97256 6554
rect 97280 6502 97290 6554
rect 97290 6502 97336 6554
rect 97040 6500 97096 6502
rect 97120 6500 97176 6502
rect 97200 6500 97256 6502
rect 97280 6500 97336 6502
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 96380 6010 96436 6012
rect 96460 6010 96516 6012
rect 96540 6010 96596 6012
rect 96620 6010 96676 6012
rect 96380 5958 96426 6010
rect 96426 5958 96436 6010
rect 96460 5958 96490 6010
rect 96490 5958 96502 6010
rect 96502 5958 96516 6010
rect 96540 5958 96554 6010
rect 96554 5958 96566 6010
rect 96566 5958 96596 6010
rect 96620 5958 96630 6010
rect 96630 5958 96676 6010
rect 96380 5956 96436 5958
rect 96460 5956 96516 5958
rect 96540 5956 96596 5958
rect 96620 5956 96676 5958
rect 66320 5466 66376 5468
rect 66400 5466 66456 5468
rect 66480 5466 66536 5468
rect 66560 5466 66616 5468
rect 66320 5414 66366 5466
rect 66366 5414 66376 5466
rect 66400 5414 66430 5466
rect 66430 5414 66442 5466
rect 66442 5414 66456 5466
rect 66480 5414 66494 5466
rect 66494 5414 66506 5466
rect 66506 5414 66536 5466
rect 66560 5414 66570 5466
rect 66570 5414 66616 5466
rect 66320 5412 66376 5414
rect 66400 5412 66456 5414
rect 66480 5412 66536 5414
rect 66560 5412 66616 5414
rect 97040 5466 97096 5468
rect 97120 5466 97176 5468
rect 97200 5466 97256 5468
rect 97280 5466 97336 5468
rect 97040 5414 97086 5466
rect 97086 5414 97096 5466
rect 97120 5414 97150 5466
rect 97150 5414 97162 5466
rect 97162 5414 97176 5466
rect 97200 5414 97214 5466
rect 97214 5414 97226 5466
rect 97226 5414 97256 5466
rect 97280 5414 97290 5466
rect 97290 5414 97336 5466
rect 97040 5412 97096 5414
rect 97120 5412 97176 5414
rect 97200 5412 97256 5414
rect 97280 5412 97336 5414
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 96380 4922 96436 4924
rect 96460 4922 96516 4924
rect 96540 4922 96596 4924
rect 96620 4922 96676 4924
rect 96380 4870 96426 4922
rect 96426 4870 96436 4922
rect 96460 4870 96490 4922
rect 96490 4870 96502 4922
rect 96502 4870 96516 4922
rect 96540 4870 96554 4922
rect 96554 4870 96566 4922
rect 96566 4870 96596 4922
rect 96620 4870 96630 4922
rect 96630 4870 96676 4922
rect 96380 4868 96436 4870
rect 96460 4868 96516 4870
rect 96540 4868 96596 4870
rect 96620 4868 96676 4870
rect 66320 4378 66376 4380
rect 66400 4378 66456 4380
rect 66480 4378 66536 4380
rect 66560 4378 66616 4380
rect 66320 4326 66366 4378
rect 66366 4326 66376 4378
rect 66400 4326 66430 4378
rect 66430 4326 66442 4378
rect 66442 4326 66456 4378
rect 66480 4326 66494 4378
rect 66494 4326 66506 4378
rect 66506 4326 66536 4378
rect 66560 4326 66570 4378
rect 66570 4326 66616 4378
rect 66320 4324 66376 4326
rect 66400 4324 66456 4326
rect 66480 4324 66536 4326
rect 66560 4324 66616 4326
rect 97040 4378 97096 4380
rect 97120 4378 97176 4380
rect 97200 4378 97256 4380
rect 97280 4378 97336 4380
rect 97040 4326 97086 4378
rect 97086 4326 97096 4378
rect 97120 4326 97150 4378
rect 97150 4326 97162 4378
rect 97162 4326 97176 4378
rect 97200 4326 97214 4378
rect 97214 4326 97226 4378
rect 97226 4326 97256 4378
rect 97280 4326 97290 4378
rect 97290 4326 97336 4378
rect 97040 4324 97096 4326
rect 97120 4324 97176 4326
rect 97200 4324 97256 4326
rect 97280 4324 97336 4326
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 96380 3834 96436 3836
rect 96460 3834 96516 3836
rect 96540 3834 96596 3836
rect 96620 3834 96676 3836
rect 96380 3782 96426 3834
rect 96426 3782 96436 3834
rect 96460 3782 96490 3834
rect 96490 3782 96502 3834
rect 96502 3782 96516 3834
rect 96540 3782 96554 3834
rect 96554 3782 96566 3834
rect 96566 3782 96596 3834
rect 96620 3782 96630 3834
rect 96630 3782 96676 3834
rect 96380 3780 96436 3782
rect 96460 3780 96516 3782
rect 96540 3780 96596 3782
rect 96620 3780 96676 3782
rect 66320 3290 66376 3292
rect 66400 3290 66456 3292
rect 66480 3290 66536 3292
rect 66560 3290 66616 3292
rect 66320 3238 66366 3290
rect 66366 3238 66376 3290
rect 66400 3238 66430 3290
rect 66430 3238 66442 3290
rect 66442 3238 66456 3290
rect 66480 3238 66494 3290
rect 66494 3238 66506 3290
rect 66506 3238 66536 3290
rect 66560 3238 66570 3290
rect 66570 3238 66616 3290
rect 66320 3236 66376 3238
rect 66400 3236 66456 3238
rect 66480 3236 66536 3238
rect 66560 3236 66616 3238
rect 97040 3290 97096 3292
rect 97120 3290 97176 3292
rect 97200 3290 97256 3292
rect 97280 3290 97336 3292
rect 97040 3238 97086 3290
rect 97086 3238 97096 3290
rect 97120 3238 97150 3290
rect 97150 3238 97162 3290
rect 97162 3238 97176 3290
rect 97200 3238 97214 3290
rect 97214 3238 97226 3290
rect 97226 3238 97256 3290
rect 97280 3238 97290 3290
rect 97290 3238 97336 3290
rect 97040 3236 97096 3238
rect 97120 3236 97176 3238
rect 97200 3236 97256 3238
rect 97280 3236 97336 3238
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 96380 2746 96436 2748
rect 96460 2746 96516 2748
rect 96540 2746 96596 2748
rect 96620 2746 96676 2748
rect 96380 2694 96426 2746
rect 96426 2694 96436 2746
rect 96460 2694 96490 2746
rect 96490 2694 96502 2746
rect 96502 2694 96516 2746
rect 96540 2694 96554 2746
rect 96554 2694 96566 2746
rect 96566 2694 96596 2746
rect 96620 2694 96630 2746
rect 96630 2694 96676 2746
rect 96380 2692 96436 2694
rect 96460 2692 96516 2694
rect 96540 2692 96596 2694
rect 96620 2692 96676 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 66320 2202 66376 2204
rect 66400 2202 66456 2204
rect 66480 2202 66536 2204
rect 66560 2202 66616 2204
rect 66320 2150 66366 2202
rect 66366 2150 66376 2202
rect 66400 2150 66430 2202
rect 66430 2150 66442 2202
rect 66442 2150 66456 2202
rect 66480 2150 66494 2202
rect 66494 2150 66506 2202
rect 66506 2150 66536 2202
rect 66560 2150 66570 2202
rect 66570 2150 66616 2202
rect 66320 2148 66376 2150
rect 66400 2148 66456 2150
rect 66480 2148 66536 2150
rect 66560 2148 66616 2150
rect 97040 2202 97096 2204
rect 97120 2202 97176 2204
rect 97200 2202 97256 2204
rect 97280 2202 97336 2204
rect 97040 2150 97086 2202
rect 97086 2150 97096 2202
rect 97120 2150 97150 2202
rect 97150 2150 97162 2202
rect 97162 2150 97176 2202
rect 97200 2150 97214 2202
rect 97214 2150 97226 2202
rect 97226 2150 97256 2202
rect 97280 2150 97290 2202
rect 97290 2150 97336 2202
rect 97040 2148 97096 2150
rect 97120 2148 97176 2150
rect 97200 2148 97256 2150
rect 97280 2148 97336 2150
<< metal3 >>
rect 4870 127328 5186 127329
rect 4870 127264 4876 127328
rect 4940 127264 4956 127328
rect 5020 127264 5036 127328
rect 5100 127264 5116 127328
rect 5180 127264 5186 127328
rect 4870 127263 5186 127264
rect 35590 127328 35906 127329
rect 35590 127264 35596 127328
rect 35660 127264 35676 127328
rect 35740 127264 35756 127328
rect 35820 127264 35836 127328
rect 35900 127264 35906 127328
rect 35590 127263 35906 127264
rect 66310 127328 66626 127329
rect 66310 127264 66316 127328
rect 66380 127264 66396 127328
rect 66460 127264 66476 127328
rect 66540 127264 66556 127328
rect 66620 127264 66626 127328
rect 66310 127263 66626 127264
rect 97030 127328 97346 127329
rect 97030 127264 97036 127328
rect 97100 127264 97116 127328
rect 97180 127264 97196 127328
rect 97260 127264 97276 127328
rect 97340 127264 97346 127328
rect 97030 127263 97346 127264
rect 4210 126784 4526 126785
rect 4210 126720 4216 126784
rect 4280 126720 4296 126784
rect 4360 126720 4376 126784
rect 4440 126720 4456 126784
rect 4520 126720 4526 126784
rect 4210 126719 4526 126720
rect 34930 126784 35246 126785
rect 34930 126720 34936 126784
rect 35000 126720 35016 126784
rect 35080 126720 35096 126784
rect 35160 126720 35176 126784
rect 35240 126720 35246 126784
rect 34930 126719 35246 126720
rect 65650 126784 65966 126785
rect 65650 126720 65656 126784
rect 65720 126720 65736 126784
rect 65800 126720 65816 126784
rect 65880 126720 65896 126784
rect 65960 126720 65966 126784
rect 65650 126719 65966 126720
rect 96370 126784 96686 126785
rect 96370 126720 96376 126784
rect 96440 126720 96456 126784
rect 96520 126720 96536 126784
rect 96600 126720 96616 126784
rect 96680 126720 96686 126784
rect 96370 126719 96686 126720
rect 105918 126784 106234 126785
rect 105918 126720 105924 126784
rect 105988 126720 106004 126784
rect 106068 126720 106084 126784
rect 106148 126720 106164 126784
rect 106228 126720 106234 126784
rect 105918 126719 106234 126720
rect 73470 126380 73476 126444
rect 73540 126442 73546 126444
rect 77293 126442 77359 126445
rect 73540 126440 77359 126442
rect 73540 126384 77298 126440
rect 77354 126384 77359 126440
rect 73540 126382 77359 126384
rect 73540 126380 73546 126382
rect 77293 126379 77359 126382
rect 4870 126240 5186 126241
rect 4870 126176 4876 126240
rect 4940 126176 4956 126240
rect 5020 126176 5036 126240
rect 5100 126176 5116 126240
rect 5180 126176 5186 126240
rect 4870 126175 5186 126176
rect 35590 126240 35906 126241
rect 35590 126176 35596 126240
rect 35660 126176 35676 126240
rect 35740 126176 35756 126240
rect 35820 126176 35836 126240
rect 35900 126176 35906 126240
rect 35590 126175 35906 126176
rect 66310 126240 66626 126241
rect 66310 126176 66316 126240
rect 66380 126176 66396 126240
rect 66460 126176 66476 126240
rect 66540 126176 66556 126240
rect 66620 126176 66626 126240
rect 66310 126175 66626 126176
rect 97030 126240 97346 126241
rect 97030 126176 97036 126240
rect 97100 126176 97116 126240
rect 97180 126176 97196 126240
rect 97260 126176 97276 126240
rect 97340 126176 97346 126240
rect 97030 126175 97346 126176
rect 106654 126240 106970 126241
rect 106654 126176 106660 126240
rect 106724 126176 106740 126240
rect 106804 126176 106820 126240
rect 106884 126176 106900 126240
rect 106964 126176 106970 126240
rect 106654 126175 106970 126176
rect 45185 126034 45251 126037
rect 46054 126034 46060 126036
rect 45185 126032 46060 126034
rect 45185 125976 45190 126032
rect 45246 125976 46060 126032
rect 45185 125974 46060 125976
rect 45185 125971 45251 125974
rect 46054 125972 46060 125974
rect 46124 125972 46130 126036
rect 53598 125972 53604 126036
rect 53668 126034 53674 126036
rect 56777 126034 56843 126037
rect 53668 126032 56843 126034
rect 53668 125976 56782 126032
rect 56838 125976 56843 126032
rect 53668 125974 56843 125976
rect 53668 125972 53674 125974
rect 56777 125971 56843 125974
rect 58566 125700 58572 125764
rect 58636 125762 58642 125764
rect 61837 125762 61903 125765
rect 58636 125760 61903 125762
rect 58636 125704 61842 125760
rect 61898 125704 61903 125760
rect 58636 125702 61903 125704
rect 58636 125700 58642 125702
rect 61837 125699 61903 125702
rect 4210 125696 4526 125697
rect 4210 125632 4216 125696
rect 4280 125632 4296 125696
rect 4360 125632 4376 125696
rect 4440 125632 4456 125696
rect 4520 125632 4526 125696
rect 4210 125631 4526 125632
rect 105918 125696 106234 125697
rect 105918 125632 105924 125696
rect 105988 125632 106004 125696
rect 106068 125632 106084 125696
rect 106148 125632 106164 125696
rect 106228 125632 106234 125696
rect 105918 125631 106234 125632
rect 49693 125626 49759 125629
rect 51022 125626 51028 125628
rect 49693 125624 51028 125626
rect 49693 125568 49698 125624
rect 49754 125568 51028 125624
rect 49693 125566 51028 125568
rect 49693 125563 49759 125566
rect 51022 125564 51028 125566
rect 51092 125564 51098 125628
rect 55990 125564 55996 125628
rect 56060 125626 56066 125628
rect 59353 125626 59419 125629
rect 56060 125624 59419 125626
rect 56060 125568 59358 125624
rect 59414 125568 59419 125624
rect 56060 125566 59419 125568
rect 56060 125564 56066 125566
rect 59353 125563 59419 125566
rect 61142 125564 61148 125628
rect 61212 125626 61218 125628
rect 63953 125626 64019 125629
rect 61212 125624 64019 125626
rect 61212 125568 63958 125624
rect 64014 125568 64019 125624
rect 61212 125566 64019 125568
rect 61212 125564 61218 125566
rect 63953 125563 64019 125566
rect 63534 125156 63540 125220
rect 63604 125218 63610 125220
rect 64413 125218 64479 125221
rect 63604 125216 64479 125218
rect 63604 125160 64418 125216
rect 64474 125160 64479 125216
rect 63604 125158 64479 125160
rect 63604 125156 63610 125158
rect 64413 125155 64479 125158
rect 4870 125152 5186 125153
rect 4870 125088 4876 125152
rect 4940 125088 4956 125152
rect 5020 125088 5036 125152
rect 5100 125088 5116 125152
rect 5180 125088 5186 125152
rect 4870 125087 5186 125088
rect 106654 125152 106970 125153
rect 106654 125088 106660 125152
rect 106724 125088 106740 125152
rect 106804 125088 106820 125152
rect 106884 125088 106900 125152
rect 106964 125088 106970 125152
rect 106654 125087 106970 125088
rect 4210 124608 4526 124609
rect 4210 124544 4216 124608
rect 4280 124544 4296 124608
rect 4360 124544 4376 124608
rect 4440 124544 4456 124608
rect 4520 124544 4526 124608
rect 4210 124543 4526 124544
rect 105918 124608 106234 124609
rect 105918 124544 105924 124608
rect 105988 124544 106004 124608
rect 106068 124544 106084 124608
rect 106148 124544 106164 124608
rect 106228 124544 106234 124608
rect 105918 124543 106234 124544
rect 36077 124268 36143 124269
rect 36069 124266 36075 124268
rect 35986 124206 36075 124266
rect 36069 124204 36075 124206
rect 36139 124204 36145 124268
rect 37733 124266 37799 124269
rect 38565 124266 38571 124268
rect 37733 124264 38571 124266
rect 37733 124208 37738 124264
rect 37794 124208 38571 124264
rect 37733 124206 38571 124208
rect 36077 124203 36143 124204
rect 37733 124203 37799 124206
rect 38565 124204 38571 124206
rect 38635 124204 38641 124268
rect 41061 124204 41067 124268
rect 41131 124266 41137 124268
rect 41321 124266 41387 124269
rect 41131 124264 41387 124266
rect 41131 124208 41326 124264
rect 41382 124208 41387 124264
rect 41131 124206 41387 124208
rect 41131 124204 41137 124206
rect 41321 124203 41387 124206
rect 48497 124268 48563 124269
rect 66069 124268 66135 124269
rect 68553 124268 68619 124269
rect 48497 124264 48544 124268
rect 48608 124266 48614 124268
rect 66021 124266 66027 124268
rect 48497 124208 48502 124264
rect 48497 124204 48544 124208
rect 48608 124206 48654 124266
rect 65978 124206 66027 124266
rect 66091 124264 66135 124268
rect 68517 124266 68523 124268
rect 66130 124208 66135 124264
rect 48608 124204 48614 124206
rect 66021 124204 66027 124206
rect 66091 124204 66135 124208
rect 68462 124206 68523 124266
rect 68587 124264 68619 124268
rect 68614 124208 68619 124264
rect 68517 124204 68523 124206
rect 68587 124204 68619 124208
rect 71013 124204 71019 124268
rect 71083 124266 71089 124268
rect 71405 124266 71471 124269
rect 71083 124264 71471 124266
rect 71083 124208 71410 124264
rect 71466 124208 71471 124264
rect 71083 124206 71471 124208
rect 71083 124204 71089 124206
rect 48497 124203 48563 124204
rect 66069 124203 66135 124204
rect 68553 124203 68619 124204
rect 71405 124203 71471 124206
rect 42333 124130 42399 124133
rect 43557 124130 43563 124132
rect 42333 124128 43563 124130
rect 42333 124072 42338 124128
rect 42394 124072 43563 124128
rect 42333 124070 43563 124072
rect 42333 124067 42399 124070
rect 43557 124068 43563 124070
rect 43627 124068 43633 124132
rect 4870 124064 5186 124065
rect 4870 124000 4876 124064
rect 4940 124000 4956 124064
rect 5020 124000 5036 124064
rect 5100 124000 5116 124064
rect 5180 124000 5186 124064
rect 4870 123999 5186 124000
rect 106654 124064 106970 124065
rect 106654 124000 106660 124064
rect 106724 124000 106740 124064
rect 106804 124000 106820 124064
rect 106884 124000 106900 124064
rect 106964 124000 106970 124064
rect 106654 123999 106970 124000
rect 86136 123932 86142 123996
rect 86206 123994 86212 123996
rect 86309 123994 86375 123997
rect 104709 123994 104775 123997
rect 86206 123992 104775 123994
rect 86206 123936 86314 123992
rect 86370 123936 104714 123992
rect 104770 123936 104775 123992
rect 86206 123934 104775 123936
rect 86206 123932 86212 123934
rect 86309 123931 86375 123934
rect 104709 123931 104775 123934
rect 87321 123860 87387 123861
rect 87304 123858 87310 123860
rect 87230 123798 87310 123858
rect 87374 123856 87387 123860
rect 87382 123800 87387 123856
rect 87304 123796 87310 123798
rect 87374 123796 87387 123800
rect 87321 123795 87387 123796
rect 96061 123860 96127 123861
rect 96061 123856 96108 123860
rect 96172 123858 96178 123860
rect 102777 123858 102843 123861
rect 96172 123856 102843 123858
rect 96061 123800 96066 123856
rect 96172 123800 102782 123856
rect 102838 123800 102843 123856
rect 96061 123796 96108 123800
rect 96172 123798 102843 123800
rect 96172 123796 96178 123798
rect 96061 123795 96127 123796
rect 102777 123795 102843 123798
rect 4210 123520 4526 123521
rect 4210 123456 4216 123520
rect 4280 123456 4296 123520
rect 4360 123456 4376 123520
rect 4440 123456 4456 123520
rect 4520 123456 4526 123520
rect 4210 123455 4526 123456
rect 105918 123520 106234 123521
rect 105918 123456 105924 123520
rect 105988 123456 106004 123520
rect 106068 123456 106084 123520
rect 106148 123456 106164 123520
rect 106228 123456 106234 123520
rect 105918 123455 106234 123456
rect 4870 122976 5186 122977
rect 4870 122912 4876 122976
rect 4940 122912 4956 122976
rect 5020 122912 5036 122976
rect 5100 122912 5116 122976
rect 5180 122912 5186 122976
rect 4870 122911 5186 122912
rect 106654 122976 106970 122977
rect 106654 122912 106660 122976
rect 106724 122912 106740 122976
rect 106804 122912 106820 122976
rect 106884 122912 106900 122976
rect 106964 122912 106970 122976
rect 106654 122911 106970 122912
rect 4210 122432 4526 122433
rect 4210 122368 4216 122432
rect 4280 122368 4296 122432
rect 4360 122368 4376 122432
rect 4440 122368 4456 122432
rect 4520 122368 4526 122432
rect 4210 122367 4526 122368
rect 105918 122432 106234 122433
rect 105918 122368 105924 122432
rect 105988 122368 106004 122432
rect 106068 122368 106084 122432
rect 106148 122368 106164 122432
rect 106228 122368 106234 122432
rect 105918 122367 106234 122368
rect 4870 121888 5186 121889
rect 4870 121824 4876 121888
rect 4940 121824 4956 121888
rect 5020 121824 5036 121888
rect 5100 121824 5116 121888
rect 5180 121824 5186 121888
rect 4870 121823 5186 121824
rect 106654 121888 106970 121889
rect 106654 121824 106660 121888
rect 106724 121824 106740 121888
rect 106804 121824 106820 121888
rect 106884 121824 106900 121888
rect 106964 121824 106970 121888
rect 106654 121823 106970 121824
rect 4210 121344 4526 121345
rect 4210 121280 4216 121344
rect 4280 121280 4296 121344
rect 4360 121280 4376 121344
rect 4440 121280 4456 121344
rect 4520 121280 4526 121344
rect 4210 121279 4526 121280
rect 105918 121344 106234 121345
rect 105918 121280 105924 121344
rect 105988 121280 106004 121344
rect 106068 121280 106084 121344
rect 106148 121280 106164 121344
rect 106228 121280 106234 121344
rect 105918 121279 106234 121280
rect 4870 120800 5186 120801
rect 4870 120736 4876 120800
rect 4940 120736 4956 120800
rect 5020 120736 5036 120800
rect 5100 120736 5116 120800
rect 5180 120736 5186 120800
rect 4870 120735 5186 120736
rect 106654 120800 106970 120801
rect 106654 120736 106660 120800
rect 106724 120736 106740 120800
rect 106804 120736 106820 120800
rect 106884 120736 106900 120800
rect 106964 120736 106970 120800
rect 106654 120735 106970 120736
rect 4210 120256 4526 120257
rect 4210 120192 4216 120256
rect 4280 120192 4296 120256
rect 4360 120192 4376 120256
rect 4440 120192 4456 120256
rect 4520 120192 4526 120256
rect 4210 120191 4526 120192
rect 105918 120256 106234 120257
rect 105918 120192 105924 120256
rect 105988 120192 106004 120256
rect 106068 120192 106084 120256
rect 106148 120192 106164 120256
rect 106228 120192 106234 120256
rect 105918 120191 106234 120192
rect 104341 119778 104407 119781
rect 102550 119776 104407 119778
rect 102550 119768 104346 119776
rect 101948 119720 104346 119768
rect 104402 119720 104407 119776
rect 101948 119718 104407 119720
rect 4870 119712 5186 119713
rect 4870 119648 4876 119712
rect 4940 119648 4956 119712
rect 5020 119648 5036 119712
rect 5100 119648 5116 119712
rect 5180 119648 5186 119712
rect 101948 119708 102610 119718
rect 104341 119715 104407 119718
rect 106654 119712 106970 119713
rect 4870 119647 5186 119648
rect 106654 119648 106660 119712
rect 106724 119648 106740 119712
rect 106804 119648 106820 119712
rect 106884 119648 106900 119712
rect 106964 119648 106970 119712
rect 106654 119647 106970 119648
rect 4210 119168 4526 119169
rect 4210 119104 4216 119168
rect 4280 119104 4296 119168
rect 4360 119104 4376 119168
rect 4440 119104 4456 119168
rect 4520 119104 4526 119168
rect 4210 119103 4526 119104
rect 105918 119168 106234 119169
rect 105918 119104 105924 119168
rect 105988 119104 106004 119168
rect 106068 119104 106084 119168
rect 106148 119104 106164 119168
rect 106228 119104 106234 119168
rect 105918 119103 106234 119104
rect 4870 118624 5186 118625
rect 4870 118560 4876 118624
rect 4940 118560 4956 118624
rect 5020 118560 5036 118624
rect 5100 118560 5116 118624
rect 5180 118560 5186 118624
rect 4870 118559 5186 118560
rect 106654 118624 106970 118625
rect 106654 118560 106660 118624
rect 106724 118560 106740 118624
rect 106804 118560 106820 118624
rect 106884 118560 106900 118624
rect 106964 118560 106970 118624
rect 106654 118559 106970 118560
rect 4210 118080 4526 118081
rect 4210 118016 4216 118080
rect 4280 118016 4296 118080
rect 4360 118016 4376 118080
rect 4440 118016 4456 118080
rect 4520 118016 4526 118080
rect 4210 118015 4526 118016
rect 105918 118080 106234 118081
rect 105918 118016 105924 118080
rect 105988 118016 106004 118080
rect 106068 118016 106084 118080
rect 106148 118016 106164 118080
rect 106228 118016 106234 118080
rect 105918 118015 106234 118016
rect 4870 117536 5186 117537
rect 4870 117472 4876 117536
rect 4940 117472 4956 117536
rect 5020 117472 5036 117536
rect 5100 117472 5116 117536
rect 5180 117472 5186 117536
rect 4870 117471 5186 117472
rect 106654 117536 106970 117537
rect 106654 117472 106660 117536
rect 106724 117472 106740 117536
rect 106804 117472 106820 117536
rect 106884 117472 106900 117536
rect 106964 117472 106970 117536
rect 106654 117471 106970 117472
rect 4210 116992 4526 116993
rect 4210 116928 4216 116992
rect 4280 116928 4296 116992
rect 4360 116928 4376 116992
rect 4440 116928 4456 116992
rect 4520 116928 4526 116992
rect 4210 116927 4526 116928
rect 105918 116992 106234 116993
rect 105918 116928 105924 116992
rect 105988 116928 106004 116992
rect 106068 116928 106084 116992
rect 106148 116928 106164 116992
rect 106228 116928 106234 116992
rect 105918 116927 106234 116928
rect 4870 116448 5186 116449
rect 4870 116384 4876 116448
rect 4940 116384 4956 116448
rect 5020 116384 5036 116448
rect 5100 116384 5116 116448
rect 5180 116384 5186 116448
rect 4870 116383 5186 116384
rect 106654 116448 106970 116449
rect 106654 116384 106660 116448
rect 106724 116384 106740 116448
rect 106804 116384 106820 116448
rect 106884 116384 106900 116448
rect 106964 116384 106970 116448
rect 106654 116383 106970 116384
rect 4210 115904 4526 115905
rect 4210 115840 4216 115904
rect 4280 115840 4296 115904
rect 4360 115840 4376 115904
rect 4440 115840 4456 115904
rect 4520 115840 4526 115904
rect 4210 115839 4526 115840
rect 105918 115904 106234 115905
rect 105918 115840 105924 115904
rect 105988 115840 106004 115904
rect 106068 115840 106084 115904
rect 106148 115840 106164 115904
rect 106228 115840 106234 115904
rect 105918 115839 106234 115840
rect 4870 115360 5186 115361
rect 4870 115296 4876 115360
rect 4940 115296 4956 115360
rect 5020 115296 5036 115360
rect 5100 115296 5116 115360
rect 5180 115296 5186 115360
rect 4870 115295 5186 115296
rect 106654 115360 106970 115361
rect 106654 115296 106660 115360
rect 106724 115296 106740 115360
rect 106804 115296 106820 115360
rect 106884 115296 106900 115360
rect 106964 115296 106970 115360
rect 106654 115295 106970 115296
rect 4210 114816 4526 114817
rect 4210 114752 4216 114816
rect 4280 114752 4296 114816
rect 4360 114752 4376 114816
rect 4440 114752 4456 114816
rect 4520 114752 4526 114816
rect 4210 114751 4526 114752
rect 105918 114816 106234 114817
rect 105918 114752 105924 114816
rect 105988 114752 106004 114816
rect 106068 114752 106084 114816
rect 106148 114752 106164 114816
rect 106228 114752 106234 114816
rect 105918 114751 106234 114752
rect 4870 114272 5186 114273
rect 4870 114208 4876 114272
rect 4940 114208 4956 114272
rect 5020 114208 5036 114272
rect 5100 114208 5116 114272
rect 5180 114208 5186 114272
rect 4870 114207 5186 114208
rect 106654 114272 106970 114273
rect 106654 114208 106660 114272
rect 106724 114208 106740 114272
rect 106804 114208 106820 114272
rect 106884 114208 106900 114272
rect 106964 114208 106970 114272
rect 106654 114207 106970 114208
rect 4210 113728 4526 113729
rect 4210 113664 4216 113728
rect 4280 113664 4296 113728
rect 4360 113664 4376 113728
rect 4440 113664 4456 113728
rect 4520 113664 4526 113728
rect 4210 113663 4526 113664
rect 105918 113728 106234 113729
rect 105918 113664 105924 113728
rect 105988 113664 106004 113728
rect 106068 113664 106084 113728
rect 106148 113664 106164 113728
rect 106228 113664 106234 113728
rect 105918 113663 106234 113664
rect 4870 113184 5186 113185
rect 4870 113120 4876 113184
rect 4940 113120 4956 113184
rect 5020 113120 5036 113184
rect 5100 113120 5116 113184
rect 5180 113120 5186 113184
rect 4870 113119 5186 113120
rect 106654 113184 106970 113185
rect 106654 113120 106660 113184
rect 106724 113120 106740 113184
rect 106804 113120 106820 113184
rect 106884 113120 106900 113184
rect 106964 113120 106970 113184
rect 106654 113119 106970 113120
rect 4210 112640 4526 112641
rect 4210 112576 4216 112640
rect 4280 112576 4296 112640
rect 4360 112576 4376 112640
rect 4440 112576 4456 112640
rect 4520 112576 4526 112640
rect 4210 112575 4526 112576
rect 105918 112640 106234 112641
rect 105918 112576 105924 112640
rect 105988 112576 106004 112640
rect 106068 112576 106084 112640
rect 106148 112576 106164 112640
rect 106228 112576 106234 112640
rect 105918 112575 106234 112576
rect 4870 112096 5186 112097
rect 4870 112032 4876 112096
rect 4940 112032 4956 112096
rect 5020 112032 5036 112096
rect 5100 112032 5116 112096
rect 5180 112032 5186 112096
rect 4870 112031 5186 112032
rect 106654 112096 106970 112097
rect 106654 112032 106660 112096
rect 106724 112032 106740 112096
rect 106804 112032 106820 112096
rect 106884 112032 106900 112096
rect 106964 112032 106970 112096
rect 106654 112031 106970 112032
rect 4210 111552 4526 111553
rect 4210 111488 4216 111552
rect 4280 111488 4296 111552
rect 4360 111488 4376 111552
rect 4440 111488 4456 111552
rect 4520 111488 4526 111552
rect 4210 111487 4526 111488
rect 105918 111552 106234 111553
rect 105918 111488 105924 111552
rect 105988 111488 106004 111552
rect 106068 111488 106084 111552
rect 106148 111488 106164 111552
rect 106228 111488 106234 111552
rect 105918 111487 106234 111488
rect 4870 111008 5186 111009
rect 4870 110944 4876 111008
rect 4940 110944 4956 111008
rect 5020 110944 5036 111008
rect 5100 110944 5116 111008
rect 5180 110944 5186 111008
rect 4870 110943 5186 110944
rect 106654 111008 106970 111009
rect 106654 110944 106660 111008
rect 106724 110944 106740 111008
rect 106804 110944 106820 111008
rect 106884 110944 106900 111008
rect 106964 110944 106970 111008
rect 106654 110943 106970 110944
rect 4210 110464 4526 110465
rect 4210 110400 4216 110464
rect 4280 110400 4296 110464
rect 4360 110400 4376 110464
rect 4440 110400 4456 110464
rect 4520 110400 4526 110464
rect 4210 110399 4526 110400
rect 105918 110464 106234 110465
rect 105918 110400 105924 110464
rect 105988 110400 106004 110464
rect 106068 110400 106084 110464
rect 106148 110400 106164 110464
rect 106228 110400 106234 110464
rect 105918 110399 106234 110400
rect 4870 109920 5186 109921
rect 4870 109856 4876 109920
rect 4940 109856 4956 109920
rect 5020 109856 5036 109920
rect 5100 109856 5116 109920
rect 5180 109856 5186 109920
rect 4870 109855 5186 109856
rect 106654 109920 106970 109921
rect 106654 109856 106660 109920
rect 106724 109856 106740 109920
rect 106804 109856 106820 109920
rect 106884 109856 106900 109920
rect 106964 109856 106970 109920
rect 106654 109855 106970 109856
rect 4210 109376 4526 109377
rect 4210 109312 4216 109376
rect 4280 109312 4296 109376
rect 4360 109312 4376 109376
rect 4440 109312 4456 109376
rect 4520 109312 4526 109376
rect 4210 109311 4526 109312
rect 105918 109376 106234 109377
rect 105918 109312 105924 109376
rect 105988 109312 106004 109376
rect 106068 109312 106084 109376
rect 106148 109312 106164 109376
rect 106228 109312 106234 109376
rect 105918 109311 106234 109312
rect 4870 108832 5186 108833
rect 4870 108768 4876 108832
rect 4940 108768 4956 108832
rect 5020 108768 5036 108832
rect 5100 108768 5116 108832
rect 5180 108768 5186 108832
rect 4870 108767 5186 108768
rect 106654 108832 106970 108833
rect 106654 108768 106660 108832
rect 106724 108768 106740 108832
rect 106804 108768 106820 108832
rect 106884 108768 106900 108832
rect 106964 108768 106970 108832
rect 106654 108767 106970 108768
rect 4210 108288 4526 108289
rect 4210 108224 4216 108288
rect 4280 108224 4296 108288
rect 4360 108224 4376 108288
rect 4440 108224 4456 108288
rect 4520 108224 4526 108288
rect 4210 108223 4526 108224
rect 105918 108288 106234 108289
rect 105918 108224 105924 108288
rect 105988 108224 106004 108288
rect 106068 108224 106084 108288
rect 106148 108224 106164 108288
rect 106228 108224 106234 108288
rect 105918 108223 106234 108224
rect 4870 107744 5186 107745
rect 4870 107680 4876 107744
rect 4940 107680 4956 107744
rect 5020 107680 5036 107744
rect 5100 107680 5116 107744
rect 5180 107680 5186 107744
rect 4870 107679 5186 107680
rect 106654 107744 106970 107745
rect 106654 107680 106660 107744
rect 106724 107680 106740 107744
rect 106804 107680 106820 107744
rect 106884 107680 106900 107744
rect 106964 107680 106970 107744
rect 106654 107679 106970 107680
rect 4210 107200 4526 107201
rect 4210 107136 4216 107200
rect 4280 107136 4296 107200
rect 4360 107136 4376 107200
rect 4440 107136 4456 107200
rect 4520 107136 4526 107200
rect 4210 107135 4526 107136
rect 105918 107200 106234 107201
rect 105918 107136 105924 107200
rect 105988 107136 106004 107200
rect 106068 107136 106084 107200
rect 106148 107136 106164 107200
rect 106228 107136 106234 107200
rect 105918 107135 106234 107136
rect 4870 106656 5186 106657
rect 4870 106592 4876 106656
rect 4940 106592 4956 106656
rect 5020 106592 5036 106656
rect 5100 106592 5116 106656
rect 5180 106592 5186 106656
rect 4870 106591 5186 106592
rect 106654 106656 106970 106657
rect 106654 106592 106660 106656
rect 106724 106592 106740 106656
rect 106804 106592 106820 106656
rect 106884 106592 106900 106656
rect 106964 106592 106970 106656
rect 106654 106591 106970 106592
rect 4210 106112 4526 106113
rect 4210 106048 4216 106112
rect 4280 106048 4296 106112
rect 4360 106048 4376 106112
rect 4440 106048 4456 106112
rect 4520 106048 4526 106112
rect 4210 106047 4526 106048
rect 105918 106112 106234 106113
rect 105918 106048 105924 106112
rect 105988 106048 106004 106112
rect 106068 106048 106084 106112
rect 106148 106048 106164 106112
rect 106228 106048 106234 106112
rect 105918 106047 106234 106048
rect 4870 105568 5186 105569
rect 4870 105504 4876 105568
rect 4940 105504 4956 105568
rect 5020 105504 5036 105568
rect 5100 105504 5116 105568
rect 5180 105504 5186 105568
rect 4870 105503 5186 105504
rect 106654 105568 106970 105569
rect 106654 105504 106660 105568
rect 106724 105504 106740 105568
rect 106804 105504 106820 105568
rect 106884 105504 106900 105568
rect 106964 105504 106970 105568
rect 106654 105503 106970 105504
rect 4210 105024 4526 105025
rect 4210 104960 4216 105024
rect 4280 104960 4296 105024
rect 4360 104960 4376 105024
rect 4440 104960 4456 105024
rect 4520 104960 4526 105024
rect 4210 104959 4526 104960
rect 105918 105024 106234 105025
rect 105918 104960 105924 105024
rect 105988 104960 106004 105024
rect 106068 104960 106084 105024
rect 106148 104960 106164 105024
rect 106228 104960 106234 105024
rect 105918 104959 106234 104960
rect 4870 104480 5186 104481
rect 4870 104416 4876 104480
rect 4940 104416 4956 104480
rect 5020 104416 5036 104480
rect 5100 104416 5116 104480
rect 5180 104416 5186 104480
rect 4870 104415 5186 104416
rect 106654 104480 106970 104481
rect 106654 104416 106660 104480
rect 106724 104416 106740 104480
rect 106804 104416 106820 104480
rect 106884 104416 106900 104480
rect 106964 104416 106970 104480
rect 106654 104415 106970 104416
rect 4210 103936 4526 103937
rect 4210 103872 4216 103936
rect 4280 103872 4296 103936
rect 4360 103872 4376 103936
rect 4440 103872 4456 103936
rect 4520 103872 4526 103936
rect 4210 103871 4526 103872
rect 105918 103936 106234 103937
rect 105918 103872 105924 103936
rect 105988 103872 106004 103936
rect 106068 103872 106084 103936
rect 106148 103872 106164 103936
rect 106228 103872 106234 103936
rect 105918 103871 106234 103872
rect 4870 103392 5186 103393
rect 4870 103328 4876 103392
rect 4940 103328 4956 103392
rect 5020 103328 5036 103392
rect 5100 103328 5116 103392
rect 5180 103328 5186 103392
rect 4870 103327 5186 103328
rect 106654 103392 106970 103393
rect 106654 103328 106660 103392
rect 106724 103328 106740 103392
rect 106804 103328 106820 103392
rect 106884 103328 106900 103392
rect 106964 103328 106970 103392
rect 106654 103327 106970 103328
rect 4210 102848 4526 102849
rect 4210 102784 4216 102848
rect 4280 102784 4296 102848
rect 4360 102784 4376 102848
rect 4440 102784 4456 102848
rect 4520 102784 4526 102848
rect 4210 102783 4526 102784
rect 105918 102848 106234 102849
rect 105918 102784 105924 102848
rect 105988 102784 106004 102848
rect 106068 102784 106084 102848
rect 106148 102784 106164 102848
rect 106228 102784 106234 102848
rect 105918 102783 106234 102784
rect 4870 102304 5186 102305
rect 4870 102240 4876 102304
rect 4940 102240 4956 102304
rect 5020 102240 5036 102304
rect 5100 102240 5116 102304
rect 5180 102240 5186 102304
rect 4870 102239 5186 102240
rect 106654 102304 106970 102305
rect 106654 102240 106660 102304
rect 106724 102240 106740 102304
rect 106804 102240 106820 102304
rect 106884 102240 106900 102304
rect 106964 102240 106970 102304
rect 106654 102239 106970 102240
rect 4210 101760 4526 101761
rect 4210 101696 4216 101760
rect 4280 101696 4296 101760
rect 4360 101696 4376 101760
rect 4440 101696 4456 101760
rect 4520 101696 4526 101760
rect 4210 101695 4526 101696
rect 105918 101760 106234 101761
rect 105918 101696 105924 101760
rect 105988 101696 106004 101760
rect 106068 101696 106084 101760
rect 106148 101696 106164 101760
rect 106228 101696 106234 101760
rect 105918 101695 106234 101696
rect 0 101418 800 101448
rect 1209 101418 1275 101421
rect 0 101416 1275 101418
rect 0 101360 1214 101416
rect 1270 101360 1275 101416
rect 0 101358 1275 101360
rect 0 101328 800 101358
rect 1209 101355 1275 101358
rect 8385 101282 8451 101285
rect 8385 101280 9506 101282
rect 8385 101224 8390 101280
rect 8446 101254 9506 101280
rect 8446 101224 10028 101254
rect 8385 101222 10028 101224
rect 8385 101219 8451 101222
rect 4870 101216 5186 101217
rect 4870 101152 4876 101216
rect 4940 101152 4956 101216
rect 5020 101152 5036 101216
rect 5100 101152 5116 101216
rect 5180 101152 5186 101216
rect 9446 101194 10028 101222
rect 106654 101216 106970 101217
rect 4870 101151 5186 101152
rect 106654 101152 106660 101216
rect 106724 101152 106740 101216
rect 106804 101152 106820 101216
rect 106884 101152 106900 101216
rect 106964 101152 106970 101216
rect 106654 101151 106970 101152
rect 4210 100672 4526 100673
rect 4210 100608 4216 100672
rect 4280 100608 4296 100672
rect 4360 100608 4376 100672
rect 4440 100608 4456 100672
rect 4520 100608 4526 100672
rect 4210 100607 4526 100608
rect 105918 100672 106234 100673
rect 105918 100608 105924 100672
rect 105988 100608 106004 100672
rect 106068 100608 106084 100672
rect 106148 100608 106164 100672
rect 106228 100608 106234 100672
rect 105918 100607 106234 100608
rect 4870 100128 5186 100129
rect 4870 100064 4876 100128
rect 4940 100064 4956 100128
rect 5020 100064 5036 100128
rect 5100 100064 5116 100128
rect 5180 100064 5186 100128
rect 4870 100063 5186 100064
rect 106654 100128 106970 100129
rect 106654 100064 106660 100128
rect 106724 100064 106740 100128
rect 106804 100064 106820 100128
rect 106884 100064 106900 100128
rect 106964 100064 106970 100128
rect 106654 100063 106970 100064
rect 4210 99584 4526 99585
rect 4210 99520 4216 99584
rect 4280 99520 4296 99584
rect 4360 99520 4376 99584
rect 4440 99520 4456 99584
rect 4520 99520 4526 99584
rect 105918 99584 106234 99585
rect 4210 99519 4526 99520
rect 8385 99514 8451 99517
rect 9446 99514 10028 99554
rect 105918 99520 105924 99584
rect 105988 99520 106004 99584
rect 106068 99520 106084 99584
rect 106148 99520 106164 99584
rect 106228 99520 106234 99584
rect 105918 99519 106234 99520
rect 8385 99512 10028 99514
rect 8385 99456 8390 99512
rect 8446 99494 10028 99512
rect 8446 99456 9506 99494
rect 8385 99454 9506 99456
rect 8385 99451 8451 99454
rect 0 99378 800 99408
rect 1393 99378 1459 99381
rect 0 99376 1459 99378
rect 0 99320 1398 99376
rect 1454 99320 1459 99376
rect 0 99318 1459 99320
rect 0 99288 800 99318
rect 1393 99315 1459 99318
rect 4870 99040 5186 99041
rect 4870 98976 4876 99040
rect 4940 98976 4956 99040
rect 5020 98976 5036 99040
rect 5100 98976 5116 99040
rect 5180 98976 5186 99040
rect 4870 98975 5186 98976
rect 106654 99040 106970 99041
rect 106654 98976 106660 99040
rect 106724 98976 106740 99040
rect 106804 98976 106820 99040
rect 106884 98976 106900 99040
rect 106964 98976 106970 99040
rect 106654 98975 106970 98976
rect 0 98698 800 98728
rect 1301 98698 1367 98701
rect 0 98696 1367 98698
rect 0 98640 1306 98696
rect 1362 98640 1367 98696
rect 0 98638 1367 98640
rect 0 98608 800 98638
rect 1301 98635 1367 98638
rect 4210 98496 4526 98497
rect 4210 98432 4216 98496
rect 4280 98432 4296 98496
rect 4360 98432 4376 98496
rect 4440 98432 4456 98496
rect 4520 98432 4526 98496
rect 4210 98431 4526 98432
rect 105918 98496 106234 98497
rect 105918 98432 105924 98496
rect 105988 98432 106004 98496
rect 106068 98432 106084 98496
rect 106148 98432 106164 98496
rect 106228 98432 106234 98496
rect 105918 98431 106234 98432
rect 8385 98426 8451 98429
rect 8385 98424 10028 98426
rect 8385 98368 8390 98424
rect 8446 98368 10028 98424
rect 8385 98366 10028 98368
rect 8385 98363 8451 98366
rect 4870 97952 5186 97953
rect 4870 97888 4876 97952
rect 4940 97888 4956 97952
rect 5020 97888 5036 97952
rect 5100 97888 5116 97952
rect 5180 97888 5186 97952
rect 4870 97887 5186 97888
rect 106654 97952 106970 97953
rect 106654 97888 106660 97952
rect 106724 97888 106740 97952
rect 106804 97888 106820 97952
rect 106884 97888 106900 97952
rect 106964 97888 106970 97952
rect 106654 97887 106970 97888
rect 4210 97408 4526 97409
rect 4210 97344 4216 97408
rect 4280 97344 4296 97408
rect 4360 97344 4376 97408
rect 4440 97344 4456 97408
rect 4520 97344 4526 97408
rect 4210 97343 4526 97344
rect 105918 97408 106234 97409
rect 105918 97344 105924 97408
rect 105988 97344 106004 97408
rect 106068 97344 106084 97408
rect 106148 97344 106164 97408
rect 106228 97344 106234 97408
rect 105918 97343 106234 97344
rect 4870 96864 5186 96865
rect 4870 96800 4876 96864
rect 4940 96800 4956 96864
rect 5020 96800 5036 96864
rect 5100 96800 5116 96864
rect 5180 96800 5186 96864
rect 4870 96799 5186 96800
rect 106654 96864 106970 96865
rect 106654 96800 106660 96864
rect 106724 96800 106740 96864
rect 106804 96800 106820 96864
rect 106884 96800 106900 96864
rect 106964 96800 106970 96864
rect 106654 96799 106970 96800
rect 8385 96794 8451 96797
rect 8385 96792 9506 96794
rect 8385 96736 8390 96792
rect 8446 96736 9506 96792
rect 8385 96734 9506 96736
rect 8385 96731 8451 96734
rect 9446 96726 9506 96734
rect 0 96658 800 96688
rect 9446 96666 10028 96726
rect 1301 96658 1367 96661
rect 0 96656 1367 96658
rect 0 96600 1306 96656
rect 1362 96600 1367 96656
rect 0 96598 1367 96600
rect 0 96568 800 96598
rect 1301 96595 1367 96598
rect 4210 96320 4526 96321
rect 4210 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4526 96320
rect 4210 96255 4526 96256
rect 105918 96320 106234 96321
rect 105918 96256 105924 96320
rect 105988 96256 106004 96320
rect 106068 96256 106084 96320
rect 106148 96256 106164 96320
rect 106228 96256 106234 96320
rect 105918 96255 106234 96256
rect 0 95978 800 96008
rect 1209 95978 1275 95981
rect 0 95976 1275 95978
rect 0 95920 1214 95976
rect 1270 95920 1275 95976
rect 0 95918 1275 95920
rect 0 95888 800 95918
rect 1209 95915 1275 95918
rect 4870 95776 5186 95777
rect 4870 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5186 95776
rect 4870 95711 5186 95712
rect 106654 95776 106970 95777
rect 106654 95712 106660 95776
rect 106724 95712 106740 95776
rect 106804 95712 106820 95776
rect 106884 95712 106900 95776
rect 106964 95712 106970 95776
rect 106654 95711 106970 95712
rect 8385 95706 8451 95709
rect 8385 95704 9506 95706
rect 8385 95648 8390 95704
rect 8446 95648 9506 95704
rect 8385 95646 9506 95648
rect 8385 95643 8451 95646
rect 9446 95643 9506 95646
rect 9446 95583 10028 95643
rect 4210 95232 4526 95233
rect 4210 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4526 95232
rect 4210 95167 4526 95168
rect 105918 95232 106234 95233
rect 105918 95168 105924 95232
rect 105988 95168 106004 95232
rect 106068 95168 106084 95232
rect 106148 95168 106164 95232
rect 106228 95168 106234 95232
rect 105918 95167 106234 95168
rect 4870 94688 5186 94689
rect 4870 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5186 94688
rect 4870 94623 5186 94624
rect 106654 94688 106970 94689
rect 106654 94624 106660 94688
rect 106724 94624 106740 94688
rect 106804 94624 106820 94688
rect 106884 94624 106900 94688
rect 106964 94624 106970 94688
rect 106654 94623 106970 94624
rect 4210 94144 4526 94145
rect 4210 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4526 94144
rect 4210 94079 4526 94080
rect 105918 94144 106234 94145
rect 105918 94080 105924 94144
rect 105988 94080 106004 94144
rect 106068 94080 106084 94144
rect 106148 94080 106164 94144
rect 106228 94080 106234 94144
rect 105918 94079 106234 94080
rect 0 93938 800 93968
rect 1301 93938 1367 93941
rect 0 93936 1367 93938
rect 0 93880 1306 93936
rect 1362 93880 1367 93936
rect 0 93878 1367 93880
rect 0 93848 800 93878
rect 1301 93875 1367 93878
rect 8385 93938 8451 93941
rect 9446 93938 10028 93963
rect 8385 93936 10028 93938
rect 8385 93880 8390 93936
rect 8446 93903 10028 93936
rect 8446 93880 9506 93903
rect 8385 93878 9506 93880
rect 8385 93875 8451 93878
rect 4870 93600 5186 93601
rect 4870 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5186 93600
rect 4870 93535 5186 93536
rect 106654 93600 106970 93601
rect 106654 93536 106660 93600
rect 106724 93536 106740 93600
rect 106804 93536 106820 93600
rect 106884 93536 106900 93600
rect 106964 93536 106970 93600
rect 106654 93535 106970 93536
rect 4210 93056 4526 93057
rect 4210 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4526 93056
rect 4210 92991 4526 92992
rect 105918 93056 106234 93057
rect 105918 92992 105924 93056
rect 105988 92992 106004 93056
rect 106068 92992 106084 93056
rect 106148 92992 106164 93056
rect 106228 92992 106234 93056
rect 105918 92991 106234 92992
rect 4870 92512 5186 92513
rect 4870 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5186 92512
rect 4870 92447 5186 92448
rect 106654 92512 106970 92513
rect 106654 92448 106660 92512
rect 106724 92448 106740 92512
rect 106804 92448 106820 92512
rect 106884 92448 106900 92512
rect 106964 92448 106970 92512
rect 106654 92447 106970 92448
rect 4210 91968 4526 91969
rect 4210 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4526 91968
rect 4210 91903 4526 91904
rect 105918 91968 106234 91969
rect 105918 91904 105924 91968
rect 105988 91904 106004 91968
rect 106068 91904 106084 91968
rect 106148 91904 106164 91968
rect 106228 91904 106234 91968
rect 105918 91903 106234 91904
rect 4870 91424 5186 91425
rect 4870 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5186 91424
rect 4870 91359 5186 91360
rect 106654 91424 106970 91425
rect 106654 91360 106660 91424
rect 106724 91360 106740 91424
rect 106804 91360 106820 91424
rect 106884 91360 106900 91424
rect 106964 91360 106970 91424
rect 106654 91359 106970 91360
rect 4210 90880 4526 90881
rect 4210 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4526 90880
rect 4210 90815 4526 90816
rect 105918 90880 106234 90881
rect 105918 90816 105924 90880
rect 105988 90816 106004 90880
rect 106068 90816 106084 90880
rect 106148 90816 106164 90880
rect 106228 90816 106234 90880
rect 105918 90815 106234 90816
rect 4870 90336 5186 90337
rect 4870 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5186 90336
rect 4870 90271 5186 90272
rect 106654 90336 106970 90337
rect 106654 90272 106660 90336
rect 106724 90272 106740 90336
rect 106804 90272 106820 90336
rect 106884 90272 106900 90336
rect 106964 90272 106970 90336
rect 106654 90271 106970 90272
rect 4210 89792 4526 89793
rect 4210 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4526 89792
rect 4210 89727 4526 89728
rect 105918 89792 106234 89793
rect 105918 89728 105924 89792
rect 105988 89728 106004 89792
rect 106068 89728 106084 89792
rect 106148 89728 106164 89792
rect 106228 89728 106234 89792
rect 105918 89727 106234 89728
rect 4870 89248 5186 89249
rect 4870 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5186 89248
rect 4870 89183 5186 89184
rect 106654 89248 106970 89249
rect 106654 89184 106660 89248
rect 106724 89184 106740 89248
rect 106804 89184 106820 89248
rect 106884 89184 106900 89248
rect 106964 89184 106970 89248
rect 106654 89183 106970 89184
rect 4210 88704 4526 88705
rect 4210 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4526 88704
rect 4210 88639 4526 88640
rect 105918 88704 106234 88705
rect 105918 88640 105924 88704
rect 105988 88640 106004 88704
rect 106068 88640 106084 88704
rect 106148 88640 106164 88704
rect 106228 88640 106234 88704
rect 105918 88639 106234 88640
rect 4870 88160 5186 88161
rect 4870 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5186 88160
rect 4870 88095 5186 88096
rect 106654 88160 106970 88161
rect 106654 88096 106660 88160
rect 106724 88096 106740 88160
rect 106804 88096 106820 88160
rect 106884 88096 106900 88160
rect 106964 88096 106970 88160
rect 106654 88095 106970 88096
rect 4210 87616 4526 87617
rect 4210 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4526 87616
rect 4210 87551 4526 87552
rect 105918 87616 106234 87617
rect 105918 87552 105924 87616
rect 105988 87552 106004 87616
rect 106068 87552 106084 87616
rect 106148 87552 106164 87616
rect 106228 87552 106234 87616
rect 105918 87551 106234 87552
rect 4870 87072 5186 87073
rect 4870 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5186 87072
rect 4870 87007 5186 87008
rect 106654 87072 106970 87073
rect 106654 87008 106660 87072
rect 106724 87008 106740 87072
rect 106804 87008 106820 87072
rect 106884 87008 106900 87072
rect 106964 87008 106970 87072
rect 106654 87007 106970 87008
rect 4210 86528 4526 86529
rect 4210 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4526 86528
rect 4210 86463 4526 86464
rect 105918 86528 106234 86529
rect 105918 86464 105924 86528
rect 105988 86464 106004 86528
rect 106068 86464 106084 86528
rect 106148 86464 106164 86528
rect 106228 86464 106234 86528
rect 105918 86463 106234 86464
rect 4870 85984 5186 85985
rect 4870 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5186 85984
rect 4870 85919 5186 85920
rect 106654 85984 106970 85985
rect 106654 85920 106660 85984
rect 106724 85920 106740 85984
rect 106804 85920 106820 85984
rect 106884 85920 106900 85984
rect 106964 85920 106970 85984
rect 106654 85919 106970 85920
rect 4210 85440 4526 85441
rect 4210 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4526 85440
rect 4210 85375 4526 85376
rect 105918 85440 106234 85441
rect 105918 85376 105924 85440
rect 105988 85376 106004 85440
rect 106068 85376 106084 85440
rect 106148 85376 106164 85440
rect 106228 85376 106234 85440
rect 105918 85375 106234 85376
rect 104617 85098 104683 85101
rect 102550 85096 104683 85098
rect 102550 85090 104622 85096
rect 101948 85040 104622 85090
rect 104678 85040 104683 85096
rect 101948 85038 104683 85040
rect 101948 85030 102610 85038
rect 104617 85035 104683 85038
rect 4870 84896 5186 84897
rect 4870 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5186 84896
rect 4870 84831 5186 84832
rect 106654 84896 106970 84897
rect 106654 84832 106660 84896
rect 106724 84832 106740 84896
rect 106804 84832 106820 84896
rect 106884 84832 106900 84896
rect 106964 84832 106970 84896
rect 106654 84831 106970 84832
rect 4210 84352 4526 84353
rect 4210 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4526 84352
rect 4210 84287 4526 84288
rect 105918 84352 106234 84353
rect 105918 84288 105924 84352
rect 105988 84288 106004 84352
rect 106068 84288 106084 84352
rect 106148 84288 106164 84352
rect 106228 84288 106234 84352
rect 105918 84287 106234 84288
rect 4870 83808 5186 83809
rect 4870 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5186 83808
rect 4870 83743 5186 83744
rect 106654 83808 106970 83809
rect 106654 83744 106660 83808
rect 106724 83744 106740 83808
rect 106804 83744 106820 83808
rect 106884 83744 106900 83808
rect 106964 83744 106970 83808
rect 106654 83743 106970 83744
rect 102041 83390 102107 83393
rect 101948 83388 102107 83390
rect 101948 83332 102046 83388
rect 102102 83332 102107 83388
rect 101948 83330 102107 83332
rect 102041 83327 102107 83330
rect 4210 83264 4526 83265
rect 4210 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4526 83264
rect 4210 83199 4526 83200
rect 105918 83264 106234 83265
rect 105918 83200 105924 83264
rect 105988 83200 106004 83264
rect 106068 83200 106084 83264
rect 106148 83200 106164 83264
rect 106228 83200 106234 83264
rect 105918 83199 106234 83200
rect 4870 82720 5186 82721
rect 4870 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5186 82720
rect 4870 82655 5186 82656
rect 106654 82720 106970 82721
rect 106654 82656 106660 82720
rect 106724 82656 106740 82720
rect 106804 82656 106820 82720
rect 106884 82656 106900 82720
rect 106964 82656 106970 82720
rect 106654 82655 106970 82656
rect 101948 82242 102610 82262
rect 103053 82242 103119 82245
rect 101948 82240 103119 82242
rect 101948 82202 103058 82240
rect 102550 82184 103058 82202
rect 103114 82184 103119 82240
rect 102550 82182 103119 82184
rect 103053 82179 103119 82182
rect 4210 82176 4526 82177
rect 4210 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4526 82176
rect 4210 82111 4526 82112
rect 105918 82176 106234 82177
rect 105918 82112 105924 82176
rect 105988 82112 106004 82176
rect 106068 82112 106084 82176
rect 106148 82112 106164 82176
rect 106228 82112 106234 82176
rect 105918 82111 106234 82112
rect 4870 81632 5186 81633
rect 4870 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5186 81632
rect 4870 81567 5186 81568
rect 106654 81632 106970 81633
rect 106654 81568 106660 81632
rect 106724 81568 106740 81632
rect 106804 81568 106820 81632
rect 106884 81568 106900 81632
rect 106964 81568 106970 81632
rect 106654 81567 106970 81568
rect 4210 81088 4526 81089
rect 4210 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4526 81088
rect 4210 81023 4526 81024
rect 105918 81088 106234 81089
rect 105918 81024 105924 81088
rect 105988 81024 106004 81088
rect 106068 81024 106084 81088
rect 106148 81024 106164 81088
rect 106228 81024 106234 81088
rect 105918 81023 106234 81024
rect 4870 80544 5186 80545
rect 4870 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5186 80544
rect 4870 80479 5186 80480
rect 106654 80544 106970 80545
rect 106654 80480 106660 80544
rect 106724 80480 106740 80544
rect 106804 80480 106820 80544
rect 106884 80480 106900 80544
rect 106964 80480 106970 80544
rect 106654 80479 106970 80480
rect 4210 80000 4526 80001
rect 4210 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4526 80000
rect 4210 79935 4526 79936
rect 105918 80000 106234 80001
rect 105918 79936 105924 80000
rect 105988 79936 106004 80000
rect 106068 79936 106084 80000
rect 106148 79936 106164 80000
rect 106228 79936 106234 80000
rect 105918 79935 106234 79936
rect 4870 79456 5186 79457
rect 4870 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5186 79456
rect 4870 79391 5186 79392
rect 106654 79456 106970 79457
rect 106654 79392 106660 79456
rect 106724 79392 106740 79456
rect 106804 79392 106820 79456
rect 106884 79392 106900 79456
rect 106964 79392 106970 79456
rect 106654 79391 106970 79392
rect 4210 78912 4526 78913
rect 4210 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4526 78912
rect 4210 78847 4526 78848
rect 105918 78912 106234 78913
rect 105918 78848 105924 78912
rect 105988 78848 106004 78912
rect 106068 78848 106084 78912
rect 106148 78848 106164 78912
rect 106228 78848 106234 78912
rect 105918 78847 106234 78848
rect 4870 78368 5186 78369
rect 0 78298 800 78328
rect 4870 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5186 78368
rect 4870 78303 5186 78304
rect 106654 78368 106970 78369
rect 106654 78304 106660 78368
rect 106724 78304 106740 78368
rect 106804 78304 106820 78368
rect 106884 78304 106900 78368
rect 106964 78304 106970 78368
rect 106654 78303 106970 78304
rect 1301 78298 1367 78301
rect 0 78296 1367 78298
rect 0 78240 1306 78296
rect 1362 78240 1367 78296
rect 0 78238 1367 78240
rect 0 78208 800 78238
rect 1301 78235 1367 78238
rect 4210 77824 4526 77825
rect 4210 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4526 77824
rect 4210 77759 4526 77760
rect 105918 77824 106234 77825
rect 105918 77760 105924 77824
rect 105988 77760 106004 77824
rect 106068 77760 106084 77824
rect 106148 77760 106164 77824
rect 106228 77760 106234 77824
rect 105918 77759 106234 77760
rect 0 77618 800 77648
rect 1301 77618 1367 77621
rect 0 77616 1367 77618
rect 0 77560 1306 77616
rect 1362 77560 1367 77616
rect 0 77558 1367 77560
rect 0 77528 800 77558
rect 1301 77555 1367 77558
rect 4870 77280 5186 77281
rect 4870 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5186 77280
rect 4870 77215 5186 77216
rect 106654 77280 106970 77281
rect 106654 77216 106660 77280
rect 106724 77216 106740 77280
rect 106804 77216 106820 77280
rect 106884 77216 106900 77280
rect 106964 77216 106970 77280
rect 106654 77215 106970 77216
rect 0 76938 800 76968
rect 1209 76938 1275 76941
rect 0 76936 1275 76938
rect 0 76880 1214 76936
rect 1270 76880 1275 76936
rect 0 76878 1275 76880
rect 0 76848 800 76878
rect 1209 76875 1275 76878
rect 4210 76736 4526 76737
rect 4210 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4526 76736
rect 4210 76671 4526 76672
rect 105918 76736 106234 76737
rect 105918 76672 105924 76736
rect 105988 76672 106004 76736
rect 106068 76672 106084 76736
rect 106148 76672 106164 76736
rect 106228 76672 106234 76736
rect 105918 76671 106234 76672
rect 0 76258 800 76288
rect 1209 76258 1275 76261
rect 0 76256 1275 76258
rect 0 76200 1214 76256
rect 1270 76200 1275 76256
rect 0 76198 1275 76200
rect 0 76168 800 76198
rect 1209 76195 1275 76198
rect 4870 76192 5186 76193
rect 4870 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5186 76192
rect 4870 76127 5186 76128
rect 106654 76192 106970 76193
rect 106654 76128 106660 76192
rect 106724 76128 106740 76192
rect 106804 76128 106820 76192
rect 106884 76128 106900 76192
rect 106964 76128 106970 76192
rect 106654 76127 106970 76128
rect 4210 75648 4526 75649
rect 0 75578 800 75608
rect 4210 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4526 75648
rect 4210 75583 4526 75584
rect 105918 75648 106234 75649
rect 105918 75584 105924 75648
rect 105988 75584 106004 75648
rect 106068 75584 106084 75648
rect 106148 75584 106164 75648
rect 106228 75584 106234 75648
rect 105918 75583 106234 75584
rect 1393 75578 1459 75581
rect 0 75576 1459 75578
rect 0 75520 1398 75576
rect 1454 75520 1459 75576
rect 0 75518 1459 75520
rect 0 75488 800 75518
rect 1393 75515 1459 75518
rect 5533 75578 5599 75581
rect 5533 75576 9506 75578
rect 5533 75520 5538 75576
rect 5594 75520 9506 75576
rect 5533 75518 9506 75520
rect 5533 75515 5599 75518
rect 9446 75483 9506 75518
rect 9446 75423 10028 75483
rect 4870 75104 5186 75105
rect 4870 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5186 75104
rect 4870 75039 5186 75040
rect 106654 75104 106970 75105
rect 106654 75040 106660 75104
rect 106724 75040 106740 75104
rect 106804 75040 106820 75104
rect 106884 75040 106900 75104
rect 106964 75040 106970 75104
rect 106654 75039 106970 75040
rect 0 74898 800 74928
rect 1301 74898 1367 74901
rect 0 74896 1367 74898
rect 0 74840 1306 74896
rect 1362 74840 1367 74896
rect 0 74838 1367 74840
rect 0 74808 800 74838
rect 1301 74835 1367 74838
rect 4210 74560 4526 74561
rect 4210 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4526 74560
rect 4210 74495 4526 74496
rect 105918 74560 106234 74561
rect 105918 74496 105924 74560
rect 105988 74496 106004 74560
rect 106068 74496 106084 74560
rect 106148 74496 106164 74560
rect 106228 74496 106234 74560
rect 105918 74495 106234 74496
rect 0 74218 800 74248
rect 1209 74218 1275 74221
rect 0 74216 1275 74218
rect 0 74160 1214 74216
rect 1270 74160 1275 74216
rect 0 74158 1275 74160
rect 0 74128 800 74158
rect 1209 74155 1275 74158
rect 4870 74016 5186 74017
rect 4870 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5186 74016
rect 4870 73951 5186 73952
rect 106654 74016 106970 74017
rect 106654 73952 106660 74016
rect 106724 73952 106740 74016
rect 106804 73952 106820 74016
rect 106884 73952 106900 74016
rect 106964 73952 106970 74016
rect 106654 73951 106970 73952
rect 0 73538 800 73568
rect 1301 73538 1367 73541
rect 0 73536 1367 73538
rect 0 73480 1306 73536
rect 1362 73480 1367 73536
rect 0 73478 1367 73480
rect 0 73448 800 73478
rect 1301 73475 1367 73478
rect 4210 73472 4526 73473
rect 4210 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4526 73472
rect 4210 73407 4526 73408
rect 105918 73472 106234 73473
rect 105918 73408 105924 73472
rect 105988 73408 106004 73472
rect 106068 73408 106084 73472
rect 106148 73408 106164 73472
rect 106228 73408 106234 73472
rect 105918 73407 106234 73408
rect 4870 72928 5186 72929
rect 0 72858 800 72888
rect 4870 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5186 72928
rect 4870 72863 5186 72864
rect 106654 72928 106970 72929
rect 106654 72864 106660 72928
rect 106724 72864 106740 72928
rect 106804 72864 106820 72928
rect 106884 72864 106900 72928
rect 106964 72864 106970 72928
rect 106654 72863 106970 72864
rect 1485 72858 1551 72861
rect 0 72856 1551 72858
rect 0 72800 1490 72856
rect 1546 72800 1551 72856
rect 0 72798 1551 72800
rect 0 72768 800 72798
rect 1485 72795 1551 72798
rect 4210 72384 4526 72385
rect 4210 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4526 72384
rect 4210 72319 4526 72320
rect 105918 72384 106234 72385
rect 105918 72320 105924 72384
rect 105988 72320 106004 72384
rect 106068 72320 106084 72384
rect 106148 72320 106164 72384
rect 106228 72320 106234 72384
rect 105918 72319 106234 72320
rect 0 72178 800 72208
rect 1301 72178 1367 72181
rect 0 72176 1367 72178
rect 0 72120 1306 72176
rect 1362 72120 1367 72176
rect 0 72118 1367 72120
rect 0 72088 800 72118
rect 1301 72115 1367 72118
rect 4870 71840 5186 71841
rect 4870 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5186 71840
rect 4870 71775 5186 71776
rect 106654 71840 106970 71841
rect 106654 71776 106660 71840
rect 106724 71776 106740 71840
rect 106804 71776 106820 71840
rect 106884 71776 106900 71840
rect 106964 71776 106970 71840
rect 106654 71775 106970 71776
rect 0 71498 800 71528
rect 1209 71498 1275 71501
rect 0 71496 1275 71498
rect 0 71440 1214 71496
rect 1270 71440 1275 71496
rect 0 71438 1275 71440
rect 0 71408 800 71438
rect 1209 71435 1275 71438
rect 4210 71296 4526 71297
rect 4210 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4526 71296
rect 4210 71231 4526 71232
rect 105918 71296 106234 71297
rect 105918 71232 105924 71296
rect 105988 71232 106004 71296
rect 106068 71232 106084 71296
rect 106148 71232 106164 71296
rect 106228 71232 106234 71296
rect 105918 71231 106234 71232
rect 0 70818 800 70848
rect 1301 70818 1367 70821
rect 0 70816 1367 70818
rect 0 70760 1306 70816
rect 1362 70760 1367 70816
rect 0 70758 1367 70760
rect 0 70728 800 70758
rect 1301 70755 1367 70758
rect 4870 70752 5186 70753
rect 4870 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5186 70752
rect 4870 70687 5186 70688
rect 106654 70752 106970 70753
rect 106654 70688 106660 70752
rect 106724 70688 106740 70752
rect 106804 70688 106820 70752
rect 106884 70688 106900 70752
rect 106964 70688 106970 70752
rect 106654 70687 106970 70688
rect 4210 70208 4526 70209
rect 0 70138 800 70168
rect 4210 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4526 70208
rect 4210 70143 4526 70144
rect 105918 70208 106234 70209
rect 105918 70144 105924 70208
rect 105988 70144 106004 70208
rect 106068 70144 106084 70208
rect 106148 70144 106164 70208
rect 106228 70144 106234 70208
rect 105918 70143 106234 70144
rect 2221 70138 2287 70141
rect 0 70136 2287 70138
rect 0 70080 2226 70136
rect 2282 70080 2287 70136
rect 0 70078 2287 70080
rect 0 70048 800 70078
rect 2221 70075 2287 70078
rect 9213 69866 9279 69869
rect 37457 69868 37523 69869
rect 38653 69868 38719 69869
rect 33944 69866 33950 69868
rect 9213 69864 33950 69866
rect 9213 69808 9218 69864
rect 9274 69808 33950 69864
rect 9213 69806 33950 69808
rect 9213 69803 9279 69806
rect 33944 69804 33950 69806
rect 34014 69804 34020 69868
rect 37448 69866 37454 69868
rect 37366 69806 37454 69866
rect 37448 69804 37454 69806
rect 37518 69804 37524 69868
rect 38616 69866 38622 69868
rect 38562 69806 38622 69866
rect 38686 69864 38719 69868
rect 38714 69808 38719 69864
rect 38616 69804 38622 69806
rect 38686 69804 38719 69808
rect 37457 69803 37523 69804
rect 38653 69803 38719 69804
rect 39757 69868 39823 69869
rect 40953 69868 41019 69869
rect 43253 69868 43319 69869
rect 39757 69864 39790 69868
rect 39854 69866 39860 69868
rect 39757 69808 39762 69864
rect 39757 69804 39790 69808
rect 39854 69806 39914 69866
rect 39854 69804 39860 69806
rect 40952 69804 40958 69868
rect 41022 69866 41028 69868
rect 41022 69806 41110 69866
rect 43253 69864 43294 69868
rect 43358 69866 43364 69868
rect 90357 69866 90423 69869
rect 90674 69866 90680 69868
rect 43253 69808 43258 69864
rect 41022 69804 41028 69806
rect 43253 69804 43294 69808
rect 43358 69806 43410 69866
rect 90357 69864 90680 69866
rect 90357 69808 90362 69864
rect 90418 69808 90680 69864
rect 90357 69806 90680 69808
rect 43358 69804 43364 69806
rect 39757 69803 39823 69804
rect 40953 69803 41019 69804
rect 43253 69803 43319 69804
rect 90357 69803 90423 69806
rect 90674 69804 90680 69806
rect 90744 69866 90750 69868
rect 104525 69866 104591 69869
rect 90744 69864 104591 69866
rect 90744 69808 104530 69864
rect 104586 69808 104591 69864
rect 90744 69806 104591 69808
rect 90744 69804 90750 69806
rect 104525 69803 104591 69806
rect 8937 69730 9003 69733
rect 8937 69728 30666 69730
rect 8937 69672 8942 69728
rect 8998 69672 30666 69728
rect 8937 69670 30666 69672
rect 8937 69667 9003 69670
rect 4870 69664 5186 69665
rect 4870 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5186 69664
rect 4870 69599 5186 69600
rect 8845 69594 8911 69597
rect 23289 69594 23355 69597
rect 23473 69596 23539 69597
rect 24669 69596 24735 69597
rect 25773 69596 25839 69597
rect 26969 69596 27035 69597
rect 8845 69592 23355 69594
rect 8845 69536 8850 69592
rect 8906 69536 23294 69592
rect 23350 69536 23355 69592
rect 8845 69534 23355 69536
rect 8845 69531 8911 69534
rect 23289 69531 23355 69534
rect 23432 69532 23438 69596
rect 23502 69594 23539 69596
rect 23502 69592 23594 69594
rect 23534 69536 23594 69592
rect 23502 69534 23594 69536
rect 23502 69532 23539 69534
rect 24618 69532 24624 69596
rect 24688 69594 24735 69596
rect 25768 69594 25774 69596
rect 24688 69592 24780 69594
rect 24730 69536 24780 69592
rect 24688 69534 24780 69536
rect 25686 69534 25774 69594
rect 24688 69532 24735 69534
rect 25768 69532 25774 69534
rect 25838 69532 25844 69596
rect 26936 69594 26942 69596
rect 26878 69534 26942 69594
rect 27006 69592 27035 69596
rect 27030 69536 27035 69592
rect 26936 69532 26942 69534
rect 27006 69532 27035 69536
rect 23473 69531 23539 69532
rect 24669 69531 24735 69532
rect 25773 69531 25839 69532
rect 26944 69531 27035 69532
rect 28073 69596 28139 69597
rect 30465 69596 30531 69597
rect 28073 69592 28110 69596
rect 28174 69594 28180 69596
rect 30440 69594 30446 69596
rect 28073 69536 28078 69592
rect 28073 69532 28110 69536
rect 28174 69534 28230 69594
rect 30374 69534 30446 69594
rect 30510 69592 30531 69596
rect 30526 69536 30531 69592
rect 28174 69532 28180 69534
rect 30440 69532 30446 69534
rect 30510 69532 30531 69536
rect 30606 69594 30666 69670
rect 106654 69664 106970 69665
rect 106654 69600 106660 69664
rect 106724 69600 106740 69664
rect 106804 69600 106820 69664
rect 106884 69600 106900 69664
rect 106964 69600 106970 69664
rect 106654 69599 106970 69600
rect 31608 69594 31614 69596
rect 30606 69534 31614 69594
rect 31608 69532 31614 69534
rect 31678 69594 31684 69596
rect 31753 69594 31819 69597
rect 32857 69596 32923 69597
rect 33961 69596 34027 69597
rect 35157 69596 35223 69597
rect 36353 69596 36419 69597
rect 42149 69596 42215 69597
rect 32806 69594 32812 69596
rect 31678 69592 31819 69594
rect 31678 69536 31758 69592
rect 31814 69536 31819 69592
rect 31678 69534 31819 69536
rect 32766 69534 32812 69594
rect 32876 69592 32923 69596
rect 33944 69594 33950 69596
rect 32918 69536 32923 69592
rect 31678 69532 31684 69534
rect 28073 69531 28139 69532
rect 30465 69531 30531 69532
rect 31753 69531 31819 69534
rect 32806 69532 32812 69534
rect 32876 69532 32923 69536
rect 33870 69534 33950 69594
rect 34014 69592 34027 69596
rect 35112 69594 35118 69596
rect 34022 69536 34027 69592
rect 33944 69532 33950 69534
rect 34014 69532 34027 69536
rect 35066 69534 35118 69594
rect 35182 69592 35223 69596
rect 36302 69594 36308 69596
rect 35218 69536 35223 69592
rect 35112 69532 35118 69534
rect 35182 69532 35223 69536
rect 36262 69534 36308 69594
rect 36372 69592 36419 69596
rect 42120 69594 42126 69596
rect 36414 69536 36419 69592
rect 36302 69532 36308 69534
rect 36372 69532 36419 69536
rect 42058 69534 42126 69594
rect 42190 69592 42215 69596
rect 42210 69536 42215 69592
rect 42120 69532 42126 69534
rect 42190 69532 42215 69536
rect 90521 69532 90527 69596
rect 90591 69594 90597 69596
rect 96889 69594 96955 69597
rect 90591 69592 96955 69594
rect 90591 69536 96894 69592
rect 96950 69536 96955 69592
rect 90591 69534 96955 69536
rect 90591 69532 90597 69534
rect 32857 69531 32923 69532
rect 33961 69531 34027 69532
rect 35157 69531 35223 69532
rect 36353 69531 36419 69532
rect 42149 69531 42215 69532
rect 96889 69531 96955 69534
rect 0 69458 800 69488
rect 1301 69458 1367 69461
rect 0 69456 1367 69458
rect 0 69400 1306 69456
rect 1362 69400 1367 69456
rect 0 69398 1367 69400
rect 0 69368 800 69398
rect 1301 69395 1367 69398
rect 9397 69458 9463 69461
rect 26944 69458 27004 69531
rect 9397 69456 27004 69458
rect 9397 69400 9402 69456
rect 9458 69400 27004 69456
rect 9397 69398 27004 69400
rect 108481 69458 108547 69461
rect 109200 69458 110000 69488
rect 108481 69456 110000 69458
rect 108481 69400 108486 69456
rect 108542 69400 110000 69456
rect 108481 69398 110000 69400
rect 9397 69395 9463 69398
rect 108481 69395 108547 69398
rect 109200 69368 110000 69398
rect 23289 69322 23355 69325
rect 29310 69322 29316 69324
rect 23289 69320 29316 69322
rect 23289 69264 23294 69320
rect 23350 69264 29316 69320
rect 23289 69262 29316 69264
rect 23289 69259 23355 69262
rect 29310 69260 29316 69262
rect 29380 69322 29386 69324
rect 29545 69322 29611 69325
rect 29380 69320 29611 69322
rect 29380 69264 29550 69320
rect 29606 69264 29611 69320
rect 29380 69262 29611 69264
rect 29380 69260 29386 69262
rect 29545 69259 29611 69262
rect 4210 69120 4526 69121
rect 4210 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4526 69120
rect 4210 69055 4526 69056
rect 105918 69120 106234 69121
rect 105918 69056 105924 69120
rect 105988 69056 106004 69120
rect 106068 69056 106084 69120
rect 106148 69056 106164 69120
rect 106228 69056 106234 69120
rect 105918 69055 106234 69056
rect 0 68778 800 68808
rect 1209 68778 1275 68781
rect 90817 68780 90883 68781
rect 90766 68778 90772 68780
rect 0 68776 1275 68778
rect 0 68720 1214 68776
rect 1270 68720 1275 68776
rect 0 68718 1275 68720
rect 90726 68718 90772 68778
rect 90836 68776 90883 68780
rect 90878 68720 90883 68776
rect 0 68688 800 68718
rect 1209 68715 1275 68718
rect 90766 68716 90772 68718
rect 90836 68716 90883 68720
rect 90817 68715 90883 68716
rect 108481 68778 108547 68781
rect 109200 68778 110000 68808
rect 108481 68776 110000 68778
rect 108481 68720 108486 68776
rect 108542 68720 110000 68776
rect 108481 68718 110000 68720
rect 108481 68715 108547 68718
rect 109200 68688 110000 68718
rect 4870 68576 5186 68577
rect 4870 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5186 68576
rect 4870 68511 5186 68512
rect 106654 68576 106970 68577
rect 106654 68512 106660 68576
rect 106724 68512 106740 68576
rect 106804 68512 106820 68576
rect 106884 68512 106900 68576
rect 106964 68512 106970 68576
rect 106654 68511 106970 68512
rect 69749 68234 69815 68237
rect 102409 68234 102475 68237
rect 69749 68232 102475 68234
rect 69749 68176 69754 68232
rect 69810 68176 102414 68232
rect 102470 68176 102475 68232
rect 69749 68174 102475 68176
rect 69749 68171 69815 68174
rect 102409 68171 102475 68174
rect 0 68098 800 68128
rect 1301 68098 1367 68101
rect 0 68096 1367 68098
rect 0 68040 1306 68096
rect 1362 68040 1367 68096
rect 0 68038 1367 68040
rect 0 68008 800 68038
rect 1301 68035 1367 68038
rect 108481 68098 108547 68101
rect 109200 68098 110000 68128
rect 108481 68096 110000 68098
rect 108481 68040 108486 68096
rect 108542 68040 110000 68096
rect 108481 68038 110000 68040
rect 108481 68035 108547 68038
rect 4210 68032 4526 68033
rect 4210 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4526 68032
rect 4210 67967 4526 67968
rect 65650 68032 65966 68033
rect 65650 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65966 68032
rect 65650 67967 65966 67968
rect 96370 68032 96686 68033
rect 96370 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96686 68032
rect 96370 67967 96686 67968
rect 105918 68032 106234 68033
rect 105918 67968 105924 68032
rect 105988 67968 106004 68032
rect 106068 67968 106084 68032
rect 106148 67968 106164 68032
rect 106228 67968 106234 68032
rect 109200 68008 110000 68038
rect 105918 67967 106234 67968
rect 95601 67826 95667 67829
rect 96981 67826 97047 67829
rect 95601 67824 97047 67826
rect 95601 67768 95606 67824
rect 95662 67768 96986 67824
rect 97042 67768 97047 67824
rect 95601 67766 97047 67768
rect 95601 67763 95667 67766
rect 96981 67763 97047 67766
rect 16062 67628 16068 67692
rect 16132 67690 16138 67692
rect 16389 67690 16455 67693
rect 16132 67688 16455 67690
rect 16132 67632 16394 67688
rect 16450 67632 16455 67688
rect 16132 67630 16455 67632
rect 16132 67628 16138 67630
rect 16389 67627 16455 67630
rect 35390 67630 36137 67690
rect 35390 67554 35450 67630
rect 22050 67494 35450 67554
rect 36077 67554 36137 67630
rect 86166 67628 86172 67692
rect 86236 67690 86242 67692
rect 90909 67690 90975 67693
rect 86236 67688 90975 67690
rect 86236 67632 90914 67688
rect 90970 67632 90975 67688
rect 86236 67630 90975 67632
rect 86236 67628 86242 67630
rect 90909 67627 90975 67630
rect 95325 67690 95391 67693
rect 96613 67690 96679 67693
rect 95325 67688 96679 67690
rect 95325 67632 95330 67688
rect 95386 67632 96618 67688
rect 96674 67632 96679 67688
rect 95325 67630 96679 67632
rect 95325 67627 95391 67630
rect 96613 67627 96679 67630
rect 96846 67630 97642 67690
rect 40401 67554 40467 67557
rect 36077 67552 40467 67554
rect 36077 67496 40406 67552
rect 40462 67496 40467 67552
rect 36077 67494 40467 67496
rect 4870 67488 5186 67489
rect 0 67418 800 67448
rect 4870 67424 4876 67488
rect 4940 67424 4956 67488
rect 5020 67424 5036 67488
rect 5100 67424 5116 67488
rect 5180 67424 5186 67488
rect 4870 67423 5186 67424
rect 1117 67418 1183 67421
rect 0 67416 1183 67418
rect 0 67360 1122 67416
rect 1178 67360 1183 67416
rect 0 67358 1183 67360
rect 0 67328 800 67358
rect 1117 67355 1183 67358
rect 8201 67418 8267 67421
rect 22050 67418 22110 67494
rect 40401 67491 40467 67494
rect 69013 67554 69079 67557
rect 79961 67554 80027 67557
rect 69013 67552 80027 67554
rect 69013 67496 69018 67552
rect 69074 67496 79966 67552
rect 80022 67496 80027 67552
rect 69013 67494 80027 67496
rect 69013 67491 69079 67494
rect 79961 67491 80027 67494
rect 90817 67554 90883 67557
rect 94773 67554 94839 67557
rect 90817 67552 94839 67554
rect 90817 67496 90822 67552
rect 90878 67496 94778 67552
rect 94834 67496 94839 67552
rect 90817 67494 94839 67496
rect 90817 67491 90883 67494
rect 94773 67491 94839 67494
rect 95785 67554 95851 67557
rect 96705 67554 96771 67557
rect 95785 67552 96771 67554
rect 95785 67496 95790 67552
rect 95846 67496 96710 67552
rect 96766 67496 96771 67552
rect 95785 67494 96771 67496
rect 95785 67491 95851 67494
rect 96705 67491 96771 67494
rect 35590 67488 35906 67489
rect 35590 67424 35596 67488
rect 35660 67424 35676 67488
rect 35740 67424 35756 67488
rect 35820 67424 35836 67488
rect 35900 67424 35906 67488
rect 35590 67423 35906 67424
rect 66310 67488 66626 67489
rect 66310 67424 66316 67488
rect 66380 67424 66396 67488
rect 66460 67424 66476 67488
rect 66540 67424 66556 67488
rect 66620 67424 66626 67488
rect 66310 67423 66626 67424
rect 8201 67416 22110 67418
rect 8201 67360 8206 67416
rect 8262 67360 22110 67416
rect 8201 67358 22110 67360
rect 75361 67418 75427 67421
rect 96846 67418 96906 67630
rect 97582 67554 97642 67630
rect 102225 67554 102291 67557
rect 97582 67552 102291 67554
rect 97582 67496 102230 67552
rect 102286 67496 102291 67552
rect 97582 67494 102291 67496
rect 102225 67491 102291 67494
rect 97030 67488 97346 67489
rect 97030 67424 97036 67488
rect 97100 67424 97116 67488
rect 97180 67424 97196 67488
rect 97260 67424 97276 67488
rect 97340 67424 97346 67488
rect 97030 67423 97346 67424
rect 106654 67488 106970 67489
rect 106654 67424 106660 67488
rect 106724 67424 106740 67488
rect 106804 67424 106820 67488
rect 106884 67424 106900 67488
rect 106964 67424 106970 67488
rect 106654 67423 106970 67424
rect 75361 67416 96906 67418
rect 75361 67360 75366 67416
rect 75422 67360 96906 67416
rect 75361 67358 96906 67360
rect 108481 67418 108547 67421
rect 109200 67418 110000 67448
rect 108481 67416 110000 67418
rect 108481 67360 108486 67416
rect 108542 67360 110000 67416
rect 108481 67358 110000 67360
rect 8201 67355 8267 67358
rect 75361 67355 75427 67358
rect 108481 67355 108547 67358
rect 109200 67328 110000 67358
rect 8017 67282 8083 67285
rect 46657 67282 46723 67285
rect 8017 67280 46723 67282
rect 8017 67224 8022 67280
rect 8078 67224 46662 67280
rect 46718 67224 46723 67280
rect 8017 67222 46723 67224
rect 8017 67219 8083 67222
rect 46657 67219 46723 67222
rect 62389 67282 62455 67285
rect 102133 67282 102199 67285
rect 62389 67280 102199 67282
rect 62389 67224 62394 67280
rect 62450 67224 102138 67280
rect 102194 67224 102199 67280
rect 62389 67222 102199 67224
rect 62389 67219 62455 67222
rect 102133 67219 102199 67222
rect 9121 67146 9187 67149
rect 44449 67146 44515 67149
rect 9121 67144 44515 67146
rect 9121 67088 9126 67144
rect 9182 67088 44454 67144
rect 44510 67088 44515 67144
rect 9121 67086 44515 67088
rect 9121 67083 9187 67086
rect 44449 67083 44515 67086
rect 62205 67146 62271 67149
rect 104341 67146 104407 67149
rect 62205 67144 104407 67146
rect 62205 67088 62210 67144
rect 62266 67088 104346 67144
rect 104402 67088 104407 67144
rect 62205 67086 104407 67088
rect 62205 67083 62271 67086
rect 104341 67083 104407 67086
rect 19333 67010 19399 67013
rect 28993 67010 29059 67013
rect 19333 67008 29059 67010
rect 19333 66952 19338 67008
rect 19394 66952 28998 67008
rect 29054 66952 29059 67008
rect 19333 66950 29059 66952
rect 19333 66947 19399 66950
rect 28993 66947 29059 66950
rect 70393 67010 70459 67013
rect 85573 67010 85639 67013
rect 70393 67008 85639 67010
rect 70393 66952 70398 67008
rect 70454 66952 85578 67008
rect 85634 66952 85639 67008
rect 70393 66950 85639 66952
rect 70393 66947 70459 66950
rect 85573 66947 85639 66950
rect 4210 66944 4526 66945
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 34930 66944 35246 66945
rect 34930 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35246 66944
rect 34930 66879 35246 66880
rect 65650 66944 65966 66945
rect 65650 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65966 66944
rect 65650 66879 65966 66880
rect 96370 66944 96686 66945
rect 96370 66880 96376 66944
rect 96440 66880 96456 66944
rect 96520 66880 96536 66944
rect 96600 66880 96616 66944
rect 96680 66880 96686 66944
rect 96370 66879 96686 66880
rect 841 66874 907 66877
rect 798 66872 907 66874
rect 798 66816 846 66872
rect 902 66816 907 66872
rect 798 66811 907 66816
rect 20345 66874 20411 66877
rect 27061 66874 27127 66877
rect 29729 66874 29795 66877
rect 20345 66872 29795 66874
rect 20345 66816 20350 66872
rect 20406 66816 27066 66872
rect 27122 66816 29734 66872
rect 29790 66816 29795 66872
rect 20345 66814 29795 66816
rect 20345 66811 20411 66814
rect 27061 66811 27127 66814
rect 29729 66811 29795 66814
rect 798 66768 858 66811
rect 0 66678 858 66768
rect 8109 66738 8175 66741
rect 39113 66738 39179 66741
rect 8109 66736 39179 66738
rect 8109 66680 8114 66736
rect 8170 66680 39118 66736
rect 39174 66680 39179 66736
rect 8109 66678 39179 66680
rect 0 66648 800 66678
rect 8109 66675 8175 66678
rect 39113 66675 39179 66678
rect 63534 66676 63540 66740
rect 63604 66738 63610 66740
rect 67541 66738 67607 66741
rect 63604 66736 67607 66738
rect 63604 66680 67546 66736
rect 67602 66680 67607 66736
rect 63604 66678 67607 66680
rect 63604 66676 63610 66678
rect 67541 66675 67607 66678
rect 84837 66738 84903 66741
rect 85389 66738 85455 66741
rect 102317 66738 102383 66741
rect 84837 66736 102383 66738
rect 84837 66680 84842 66736
rect 84898 66680 85394 66736
rect 85450 66680 102322 66736
rect 102378 66680 102383 66736
rect 84837 66678 102383 66680
rect 84837 66675 84903 66678
rect 85389 66675 85455 66678
rect 102317 66675 102383 66678
rect 108481 66738 108547 66741
rect 109200 66738 110000 66768
rect 108481 66736 110000 66738
rect 108481 66680 108486 66736
rect 108542 66680 110000 66736
rect 108481 66678 110000 66680
rect 108481 66675 108547 66678
rect 109200 66648 110000 66678
rect 33041 66602 33107 66605
rect 33869 66602 33935 66605
rect 33041 66600 33935 66602
rect 33041 66544 33046 66600
rect 33102 66544 33874 66600
rect 33930 66544 33935 66600
rect 33041 66542 33935 66544
rect 33041 66539 33107 66542
rect 33869 66539 33935 66542
rect 35341 66602 35407 66605
rect 36118 66602 36124 66604
rect 35341 66600 36124 66602
rect 35341 66544 35346 66600
rect 35402 66544 36124 66600
rect 35341 66542 36124 66544
rect 35341 66539 35407 66542
rect 36118 66540 36124 66542
rect 36188 66540 36194 66604
rect 47853 66602 47919 66605
rect 51022 66602 51028 66604
rect 47853 66600 51028 66602
rect 47853 66544 47858 66600
rect 47914 66544 51028 66600
rect 47853 66542 51028 66544
rect 47853 66539 47919 66542
rect 51022 66540 51028 66542
rect 51092 66540 51098 66604
rect 66110 66540 66116 66604
rect 66180 66602 66186 66604
rect 67633 66602 67699 66605
rect 66180 66600 67699 66602
rect 66180 66544 67638 66600
rect 67694 66544 67699 66600
rect 66180 66542 67699 66544
rect 66180 66540 66186 66542
rect 67633 66539 67699 66542
rect 84653 66602 84719 66605
rect 106181 66602 106247 66605
rect 84653 66600 106247 66602
rect 84653 66544 84658 66600
rect 84714 66544 106186 66600
rect 106242 66544 106247 66600
rect 84653 66542 106247 66544
rect 84653 66539 84719 66542
rect 106181 66539 106247 66542
rect 87965 66466 88031 66469
rect 88517 66466 88583 66469
rect 87965 66464 88583 66466
rect 87965 66408 87970 66464
rect 88026 66408 88522 66464
rect 88578 66408 88583 66464
rect 87965 66406 88583 66408
rect 87965 66403 88031 66406
rect 88517 66403 88583 66406
rect 4870 66400 5186 66401
rect 4870 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5186 66400
rect 4870 66335 5186 66336
rect 35590 66400 35906 66401
rect 35590 66336 35596 66400
rect 35660 66336 35676 66400
rect 35740 66336 35756 66400
rect 35820 66336 35836 66400
rect 35900 66336 35906 66400
rect 35590 66335 35906 66336
rect 66310 66400 66626 66401
rect 66310 66336 66316 66400
rect 66380 66336 66396 66400
rect 66460 66336 66476 66400
rect 66540 66336 66556 66400
rect 66620 66336 66626 66400
rect 66310 66335 66626 66336
rect 97030 66400 97346 66401
rect 97030 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97346 66400
rect 97030 66335 97346 66336
rect 106654 66400 106970 66401
rect 106654 66336 106660 66400
rect 106724 66336 106740 66400
rect 106804 66336 106820 66400
rect 106884 66336 106900 66400
rect 106964 66336 106970 66400
rect 106654 66335 106970 66336
rect 39021 66330 39087 66333
rect 41086 66330 41092 66332
rect 39021 66328 41092 66330
rect 39021 66272 39026 66328
rect 39082 66272 41092 66328
rect 39021 66270 41092 66272
rect 39021 66267 39087 66270
rect 41086 66268 41092 66270
rect 41156 66268 41162 66332
rect 71078 66268 71084 66332
rect 71148 66330 71154 66332
rect 73705 66330 73771 66333
rect 71148 66328 73771 66330
rect 71148 66272 73710 66328
rect 73766 66272 73771 66328
rect 71148 66270 73771 66272
rect 71148 66268 71154 66270
rect 73705 66267 73771 66270
rect 87270 66268 87276 66332
rect 87340 66330 87346 66332
rect 91001 66330 91067 66333
rect 87340 66328 91067 66330
rect 87340 66272 91006 66328
rect 91062 66272 91067 66328
rect 87340 66270 91067 66272
rect 87340 66268 87346 66270
rect 91001 66267 91067 66270
rect 45737 66194 45803 66197
rect 46054 66194 46060 66196
rect 45737 66192 46060 66194
rect 45737 66136 45742 66192
rect 45798 66136 46060 66192
rect 45737 66134 46060 66136
rect 45737 66131 45803 66134
rect 46054 66132 46060 66134
rect 46124 66132 46130 66196
rect 0 66058 800 66088
rect 108481 66058 108547 66061
rect 109200 66058 110000 66088
rect 0 65968 858 66058
rect 108481 66056 110000 66058
rect 108481 66000 108486 66056
rect 108542 66000 110000 66056
rect 108481 65998 110000 66000
rect 108481 65995 108547 65998
rect 109200 65968 110000 65998
rect 798 65925 858 65968
rect 798 65920 907 65925
rect 53649 65924 53715 65925
rect 798 65864 846 65920
rect 902 65864 907 65920
rect 798 65862 907 65864
rect 841 65859 907 65862
rect 53598 65860 53604 65924
rect 53668 65922 53715 65924
rect 53668 65920 53760 65922
rect 53710 65864 53760 65920
rect 53668 65862 53760 65864
rect 53668 65860 53715 65862
rect 53649 65859 53715 65860
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 34930 65856 35246 65857
rect 34930 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35246 65856
rect 34930 65791 35246 65792
rect 65650 65856 65966 65857
rect 65650 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65966 65856
rect 65650 65791 65966 65792
rect 96370 65856 96686 65857
rect 96370 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96686 65856
rect 96370 65791 96686 65792
rect 105918 65856 106234 65857
rect 105918 65792 105924 65856
rect 105988 65792 106004 65856
rect 106068 65792 106084 65856
rect 106148 65792 106164 65856
rect 106228 65792 106234 65856
rect 105918 65791 106234 65792
rect 841 65514 907 65517
rect 798 65512 907 65514
rect 798 65456 846 65512
rect 902 65456 907 65512
rect 798 65451 907 65456
rect 33501 65514 33567 65517
rect 43478 65514 43484 65516
rect 33501 65512 43484 65514
rect 33501 65456 33506 65512
rect 33562 65456 43484 65512
rect 33501 65454 43484 65456
rect 33501 65451 33567 65454
rect 43478 65452 43484 65454
rect 43548 65452 43554 65516
rect 73470 65452 73476 65516
rect 73540 65514 73546 65516
rect 84929 65514 84995 65517
rect 73540 65512 84995 65514
rect 73540 65456 84934 65512
rect 84990 65456 84995 65512
rect 73540 65454 84995 65456
rect 73540 65452 73546 65454
rect 84929 65451 84995 65454
rect 798 65408 858 65451
rect 0 65318 858 65408
rect 108481 65378 108547 65381
rect 109200 65378 110000 65408
rect 108481 65376 110000 65378
rect 108481 65320 108486 65376
rect 108542 65320 110000 65376
rect 108481 65318 110000 65320
rect 0 65288 800 65318
rect 108481 65315 108547 65318
rect 4870 65312 5186 65313
rect 4870 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5186 65312
rect 4870 65247 5186 65248
rect 106654 65312 106970 65313
rect 106654 65248 106660 65312
rect 106724 65248 106740 65312
rect 106804 65248 106820 65312
rect 106884 65248 106900 65312
rect 106964 65248 106970 65312
rect 109200 65288 110000 65318
rect 106654 65247 106970 65248
rect 4210 64768 4526 64769
rect 0 64698 800 64728
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 105918 64768 106234 64769
rect 105918 64704 105924 64768
rect 105988 64704 106004 64768
rect 106068 64704 106084 64768
rect 106148 64704 106164 64768
rect 106228 64704 106234 64768
rect 105918 64703 106234 64704
rect 1393 64698 1459 64701
rect 0 64696 1459 64698
rect 0 64640 1398 64696
rect 1454 64640 1459 64696
rect 0 64638 1459 64640
rect 0 64608 800 64638
rect 1393 64635 1459 64638
rect 108481 64698 108547 64701
rect 109200 64698 110000 64728
rect 108481 64696 110000 64698
rect 108481 64640 108486 64696
rect 108542 64640 110000 64696
rect 108481 64638 110000 64640
rect 108481 64635 108547 64638
rect 109200 64608 110000 64638
rect 4870 64224 5186 64225
rect 4870 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5186 64224
rect 4870 64159 5186 64160
rect 106654 64224 106970 64225
rect 106654 64160 106660 64224
rect 106724 64160 106740 64224
rect 106804 64160 106820 64224
rect 106884 64160 106900 64224
rect 106964 64160 106970 64224
rect 106654 64159 106970 64160
rect 841 64154 907 64157
rect 798 64152 907 64154
rect 798 64096 846 64152
rect 902 64096 907 64152
rect 798 64091 907 64096
rect 35985 64154 36051 64157
rect 38565 64154 38571 64156
rect 35985 64152 38571 64154
rect 35985 64096 35990 64152
rect 36046 64096 38571 64152
rect 35985 64094 38571 64096
rect 35985 64091 36051 64094
rect 38565 64092 38571 64094
rect 38635 64092 38641 64156
rect 47485 64154 47551 64157
rect 48538 64154 48544 64156
rect 47485 64152 48544 64154
rect 47485 64096 47490 64152
rect 47546 64096 48544 64152
rect 47485 64094 48544 64096
rect 47485 64091 47551 64094
rect 48538 64092 48544 64094
rect 48608 64092 48614 64156
rect 56037 64092 56043 64156
rect 56107 64154 56113 64156
rect 63401 64154 63467 64157
rect 56107 64152 63467 64154
rect 56107 64096 63406 64152
rect 63462 64096 63467 64152
rect 56107 64094 63467 64096
rect 56107 64092 56113 64094
rect 63401 64091 63467 64094
rect 68517 64092 68523 64156
rect 68587 64154 68593 64156
rect 75453 64154 75519 64157
rect 68587 64152 75519 64154
rect 68587 64096 75458 64152
rect 75514 64096 75519 64152
rect 68587 64094 75519 64096
rect 68587 64092 68593 64094
rect 75453 64091 75519 64094
rect 798 64048 858 64091
rect 0 63958 858 64048
rect 0 63928 800 63958
rect 58533 63956 58539 64020
rect 58603 64018 58609 64020
rect 66161 64018 66227 64021
rect 58603 64016 66227 64018
rect 58603 63960 66166 64016
rect 66222 63960 66227 64016
rect 58603 63958 66227 63960
rect 58603 63956 58609 63958
rect 66161 63955 66227 63958
rect 108481 64018 108547 64021
rect 109200 64018 110000 64048
rect 108481 64016 110000 64018
rect 108481 63960 108486 64016
rect 108542 63960 110000 64016
rect 108481 63958 110000 63960
rect 108481 63955 108547 63958
rect 109200 63928 110000 63958
rect 61050 63820 61056 63884
rect 61120 63882 61126 63884
rect 71865 63882 71931 63885
rect 61120 63880 71931 63882
rect 61120 63824 71870 63880
rect 71926 63824 71931 63880
rect 61120 63822 71931 63824
rect 61120 63820 61126 63822
rect 71865 63819 71931 63822
rect 95852 63820 95858 63884
rect 95922 63882 95928 63884
rect 96153 63882 96219 63885
rect 105629 63882 105695 63885
rect 95922 63880 105695 63882
rect 95922 63824 96158 63880
rect 96214 63824 105634 63880
rect 105690 63824 105695 63880
rect 95922 63822 105695 63824
rect 95922 63820 95928 63822
rect 96153 63819 96219 63822
rect 105629 63819 105695 63822
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 105918 63680 106234 63681
rect 105918 63616 105924 63680
rect 105988 63616 106004 63680
rect 106068 63616 106084 63680
rect 106148 63616 106164 63680
rect 106228 63616 106234 63680
rect 105918 63615 106234 63616
rect 841 63474 907 63477
rect 798 63472 907 63474
rect 798 63416 846 63472
rect 902 63416 907 63472
rect 798 63411 907 63416
rect 798 63368 858 63411
rect 0 63278 858 63368
rect 0 63248 800 63278
rect 4870 63136 5186 63137
rect 4870 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5186 63136
rect 4870 63071 5186 63072
rect 106654 63136 106970 63137
rect 106654 63072 106660 63136
rect 106724 63072 106740 63136
rect 106804 63072 106820 63136
rect 106884 63072 106900 63136
rect 106964 63072 106970 63136
rect 106654 63071 106970 63072
rect 841 62794 907 62797
rect 798 62792 907 62794
rect 798 62736 846 62792
rect 902 62736 907 62792
rect 798 62731 907 62736
rect 798 62688 858 62731
rect 0 62598 858 62688
rect 0 62568 800 62598
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 4210 62527 4526 62528
rect 105918 62592 106234 62593
rect 105918 62528 105924 62592
rect 105988 62528 106004 62592
rect 106068 62528 106084 62592
rect 106148 62528 106164 62592
rect 106228 62528 106234 62592
rect 105918 62527 106234 62528
rect 4870 62048 5186 62049
rect 0 61978 800 62008
rect 4870 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5186 62048
rect 4870 61983 5186 61984
rect 106654 62048 106970 62049
rect 106654 61984 106660 62048
rect 106724 61984 106740 62048
rect 106804 61984 106820 62048
rect 106884 61984 106900 62048
rect 106964 61984 106970 62048
rect 106654 61983 106970 61984
rect 1485 61978 1551 61981
rect 0 61976 1551 61978
rect 0 61920 1490 61976
rect 1546 61920 1551 61976
rect 0 61918 1551 61920
rect 0 61888 800 61918
rect 1485 61915 1551 61918
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 105918 61504 106234 61505
rect 105918 61440 105924 61504
rect 105988 61440 106004 61504
rect 106068 61440 106084 61504
rect 106148 61440 106164 61504
rect 106228 61440 106234 61504
rect 105918 61439 106234 61440
rect 0 61298 800 61328
rect 1301 61298 1367 61301
rect 0 61296 1367 61298
rect 0 61240 1306 61296
rect 1362 61240 1367 61296
rect 0 61238 1367 61240
rect 0 61208 800 61238
rect 1301 61235 1367 61238
rect 4870 60960 5186 60961
rect 4870 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5186 60960
rect 4870 60895 5186 60896
rect 106654 60960 106970 60961
rect 106654 60896 106660 60960
rect 106724 60896 106740 60960
rect 106804 60896 106820 60960
rect 106884 60896 106900 60960
rect 106964 60896 106970 60960
rect 106654 60895 106970 60896
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 105918 60416 106234 60417
rect 105918 60352 105924 60416
rect 105988 60352 106004 60416
rect 106068 60352 106084 60416
rect 106148 60352 106164 60416
rect 106228 60352 106234 60416
rect 105918 60351 106234 60352
rect 4870 59872 5186 59873
rect 4870 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5186 59872
rect 4870 59807 5186 59808
rect 106654 59872 106970 59873
rect 106654 59808 106660 59872
rect 106724 59808 106740 59872
rect 106804 59808 106820 59872
rect 106884 59808 106900 59872
rect 106964 59808 106970 59872
rect 106654 59807 106970 59808
rect 103973 59802 104039 59805
rect 102550 59800 104039 59802
rect 102550 59768 103978 59800
rect 101948 59744 103978 59768
rect 104034 59744 104039 59800
rect 101948 59742 104039 59744
rect 101948 59708 102610 59742
rect 103973 59739 104039 59742
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 105918 59328 106234 59329
rect 105918 59264 105924 59328
rect 105988 59264 106004 59328
rect 106068 59264 106084 59328
rect 106148 59264 106164 59328
rect 106228 59264 106234 59328
rect 105918 59263 106234 59264
rect 4870 58784 5186 58785
rect 4870 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5186 58784
rect 4870 58719 5186 58720
rect 106654 58784 106970 58785
rect 106654 58720 106660 58784
rect 106724 58720 106740 58784
rect 106804 58720 106820 58784
rect 106884 58720 106900 58784
rect 106964 58720 106970 58784
rect 106654 58719 106970 58720
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 105918 58240 106234 58241
rect 105918 58176 105924 58240
rect 105988 58176 106004 58240
rect 106068 58176 106084 58240
rect 106148 58176 106164 58240
rect 106228 58176 106234 58240
rect 105918 58175 106234 58176
rect 4870 57696 5186 57697
rect 4870 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5186 57696
rect 4870 57631 5186 57632
rect 106654 57696 106970 57697
rect 106654 57632 106660 57696
rect 106724 57632 106740 57696
rect 106804 57632 106820 57696
rect 106884 57632 106900 57696
rect 106964 57632 106970 57696
rect 106654 57631 106970 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 105918 57152 106234 57153
rect 105918 57088 105924 57152
rect 105988 57088 106004 57152
rect 106068 57088 106084 57152
rect 106148 57088 106164 57152
rect 106228 57088 106234 57152
rect 105918 57087 106234 57088
rect 4870 56608 5186 56609
rect 4870 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5186 56608
rect 4870 56543 5186 56544
rect 106654 56608 106970 56609
rect 106654 56544 106660 56608
rect 106724 56544 106740 56608
rect 106804 56544 106820 56608
rect 106884 56544 106900 56608
rect 106964 56544 106970 56608
rect 106654 56543 106970 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 105918 56064 106234 56065
rect 105918 56000 105924 56064
rect 105988 56000 106004 56064
rect 106068 56000 106084 56064
rect 106148 56000 106164 56064
rect 106228 56000 106234 56064
rect 105918 55999 106234 56000
rect 4870 55520 5186 55521
rect 4870 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5186 55520
rect 4870 55455 5186 55456
rect 106654 55520 106970 55521
rect 106654 55456 106660 55520
rect 106724 55456 106740 55520
rect 106804 55456 106820 55520
rect 106884 55456 106900 55520
rect 106964 55456 106970 55520
rect 106654 55455 106970 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 105918 54976 106234 54977
rect 105918 54912 105924 54976
rect 105988 54912 106004 54976
rect 106068 54912 106084 54976
rect 106148 54912 106164 54976
rect 106228 54912 106234 54976
rect 105918 54911 106234 54912
rect 4870 54432 5186 54433
rect 4870 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5186 54432
rect 4870 54367 5186 54368
rect 106654 54432 106970 54433
rect 106654 54368 106660 54432
rect 106724 54368 106740 54432
rect 106804 54368 106820 54432
rect 106884 54368 106900 54432
rect 106964 54368 106970 54432
rect 106654 54367 106970 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 105918 53888 106234 53889
rect 105918 53824 105924 53888
rect 105988 53824 106004 53888
rect 106068 53824 106084 53888
rect 106148 53824 106164 53888
rect 106228 53824 106234 53888
rect 105918 53823 106234 53824
rect 4870 53344 5186 53345
rect 4870 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5186 53344
rect 4870 53279 5186 53280
rect 106654 53344 106970 53345
rect 106654 53280 106660 53344
rect 106724 53280 106740 53344
rect 106804 53280 106820 53344
rect 106884 53280 106900 53344
rect 106964 53280 106970 53344
rect 106654 53279 106970 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 105918 52800 106234 52801
rect 105918 52736 105924 52800
rect 105988 52736 106004 52800
rect 106068 52736 106084 52800
rect 106148 52736 106164 52800
rect 106228 52736 106234 52800
rect 105918 52735 106234 52736
rect 4870 52256 5186 52257
rect 4870 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5186 52256
rect 4870 52191 5186 52192
rect 106654 52256 106970 52257
rect 106654 52192 106660 52256
rect 106724 52192 106740 52256
rect 106804 52192 106820 52256
rect 106884 52192 106900 52256
rect 106964 52192 106970 52256
rect 106654 52191 106970 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 105918 51712 106234 51713
rect 105918 51648 105924 51712
rect 105988 51648 106004 51712
rect 106068 51648 106084 51712
rect 106148 51648 106164 51712
rect 106228 51648 106234 51712
rect 105918 51647 106234 51648
rect 4870 51168 5186 51169
rect 4870 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5186 51168
rect 4870 51103 5186 51104
rect 106654 51168 106970 51169
rect 106654 51104 106660 51168
rect 106724 51104 106740 51168
rect 106804 51104 106820 51168
rect 106884 51104 106900 51168
rect 106964 51104 106970 51168
rect 106654 51103 106970 51104
rect 108481 51098 108547 51101
rect 109200 51098 110000 51128
rect 108481 51096 110000 51098
rect 108481 51040 108486 51096
rect 108542 51040 110000 51096
rect 108481 51038 110000 51040
rect 108481 51035 108547 51038
rect 109200 51008 110000 51038
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 105918 50624 106234 50625
rect 105918 50560 105924 50624
rect 105988 50560 106004 50624
rect 106068 50560 106084 50624
rect 106148 50560 106164 50624
rect 106228 50560 106234 50624
rect 105918 50559 106234 50560
rect 4870 50080 5186 50081
rect 4870 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5186 50080
rect 4870 50015 5186 50016
rect 106654 50080 106970 50081
rect 106654 50016 106660 50080
rect 106724 50016 106740 50080
rect 106804 50016 106820 50080
rect 106884 50016 106900 50080
rect 106964 50016 106970 50080
rect 106654 50015 106970 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 105918 49536 106234 49537
rect 105918 49472 105924 49536
rect 105988 49472 106004 49536
rect 106068 49472 106084 49536
rect 106148 49472 106164 49536
rect 106228 49472 106234 49536
rect 105918 49471 106234 49472
rect 4870 48992 5186 48993
rect 4870 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5186 48992
rect 4870 48927 5186 48928
rect 106654 48992 106970 48993
rect 106654 48928 106660 48992
rect 106724 48928 106740 48992
rect 106804 48928 106820 48992
rect 106884 48928 106900 48992
rect 106964 48928 106970 48992
rect 106654 48927 106970 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 105918 48448 106234 48449
rect 105918 48384 105924 48448
rect 105988 48384 106004 48448
rect 106068 48384 106084 48448
rect 106148 48384 106164 48448
rect 106228 48384 106234 48448
rect 105918 48383 106234 48384
rect 4870 47904 5186 47905
rect 4870 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5186 47904
rect 4870 47839 5186 47840
rect 106654 47904 106970 47905
rect 106654 47840 106660 47904
rect 106724 47840 106740 47904
rect 106804 47840 106820 47904
rect 106884 47840 106900 47904
rect 106964 47840 106970 47904
rect 106654 47839 106970 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 105918 47360 106234 47361
rect 105918 47296 105924 47360
rect 105988 47296 106004 47360
rect 106068 47296 106084 47360
rect 106148 47296 106164 47360
rect 106228 47296 106234 47360
rect 105918 47295 106234 47296
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 106654 46816 106970 46817
rect 106654 46752 106660 46816
rect 106724 46752 106740 46816
rect 106804 46752 106820 46816
rect 106884 46752 106900 46816
rect 106964 46752 106970 46816
rect 106654 46751 106970 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 105918 46272 106234 46273
rect 105918 46208 105924 46272
rect 105988 46208 106004 46272
rect 106068 46208 106084 46272
rect 106148 46208 106164 46272
rect 106228 46208 106234 46272
rect 105918 46207 106234 46208
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 106654 45728 106970 45729
rect 106654 45664 106660 45728
rect 106724 45664 106740 45728
rect 106804 45664 106820 45728
rect 106884 45664 106900 45728
rect 106964 45664 106970 45728
rect 106654 45663 106970 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 105918 45184 106234 45185
rect 105918 45120 105924 45184
rect 105988 45120 106004 45184
rect 106068 45120 106084 45184
rect 106148 45120 106164 45184
rect 106228 45120 106234 45184
rect 105918 45119 106234 45120
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 106654 44640 106970 44641
rect 106654 44576 106660 44640
rect 106724 44576 106740 44640
rect 106804 44576 106820 44640
rect 106884 44576 106900 44640
rect 106964 44576 106970 44640
rect 106654 44575 106970 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 105918 44096 106234 44097
rect 105918 44032 105924 44096
rect 105988 44032 106004 44096
rect 106068 44032 106084 44096
rect 106148 44032 106164 44096
rect 106228 44032 106234 44096
rect 105918 44031 106234 44032
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 106654 43552 106970 43553
rect 106654 43488 106660 43552
rect 106724 43488 106740 43552
rect 106804 43488 106820 43552
rect 106884 43488 106900 43552
rect 106964 43488 106970 43552
rect 106654 43487 106970 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 105918 43008 106234 43009
rect 105918 42944 105924 43008
rect 105988 42944 106004 43008
rect 106068 42944 106084 43008
rect 106148 42944 106164 43008
rect 106228 42944 106234 43008
rect 105918 42943 106234 42944
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 106654 42464 106970 42465
rect 106654 42400 106660 42464
rect 106724 42400 106740 42464
rect 106804 42400 106820 42464
rect 106884 42400 106900 42464
rect 106964 42400 106970 42464
rect 106654 42399 106970 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 105918 41920 106234 41921
rect 105918 41856 105924 41920
rect 105988 41856 106004 41920
rect 106068 41856 106084 41920
rect 106148 41856 106164 41920
rect 106228 41856 106234 41920
rect 105918 41855 106234 41856
rect 0 41578 800 41608
rect 1209 41578 1275 41581
rect 0 41576 1275 41578
rect 0 41520 1214 41576
rect 1270 41520 1275 41576
rect 0 41518 1275 41520
rect 0 41488 800 41518
rect 1209 41515 1275 41518
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 106654 41376 106970 41377
rect 106654 41312 106660 41376
rect 106724 41312 106740 41376
rect 106804 41312 106820 41376
rect 106884 41312 106900 41376
rect 106964 41312 106970 41376
rect 106654 41311 106970 41312
rect 5533 41306 5599 41309
rect 5533 41304 9506 41306
rect 5533 41248 5538 41304
rect 5594 41254 9506 41304
rect 5594 41248 10028 41254
rect 5533 41246 10028 41248
rect 5533 41243 5599 41246
rect 9446 41194 10028 41246
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 105918 40832 106234 40833
rect 105918 40768 105924 40832
rect 105988 40768 106004 40832
rect 106068 40768 106084 40832
rect 106148 40768 106164 40832
rect 106228 40768 106234 40832
rect 105918 40767 106234 40768
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 106654 40288 106970 40289
rect 106654 40224 106660 40288
rect 106724 40224 106740 40288
rect 106804 40224 106820 40288
rect 106884 40224 106900 40288
rect 106964 40224 106970 40288
rect 106654 40223 106970 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 105918 39744 106234 39745
rect 105918 39680 105924 39744
rect 105988 39680 106004 39744
rect 106068 39680 106084 39744
rect 106148 39680 106164 39744
rect 106228 39680 106234 39744
rect 105918 39679 106234 39680
rect 5533 39674 5599 39677
rect 5533 39672 9506 39674
rect 5533 39616 5538 39672
rect 5594 39616 9506 39672
rect 5533 39614 9506 39616
rect 5533 39611 5599 39614
rect 0 39538 800 39568
rect 9446 39554 9506 39614
rect 1393 39538 1459 39541
rect 0 39536 1459 39538
rect 0 39480 1398 39536
rect 1454 39480 1459 39536
rect 9446 39494 10028 39554
rect 0 39478 1459 39480
rect 0 39448 800 39478
rect 1393 39475 1459 39478
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 106654 39200 106970 39201
rect 106654 39136 106660 39200
rect 106724 39136 106740 39200
rect 106804 39136 106820 39200
rect 106884 39136 106900 39200
rect 106964 39136 106970 39200
rect 106654 39135 106970 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 105918 38656 106234 38657
rect 105918 38592 105924 38656
rect 105988 38592 106004 38656
rect 106068 38592 106084 38656
rect 106148 38592 106164 38656
rect 106228 38592 106234 38656
rect 105918 38591 106234 38592
rect 8385 38450 8451 38453
rect 8385 38448 9506 38450
rect 8385 38392 8390 38448
rect 8446 38426 9506 38448
rect 8446 38392 10028 38426
rect 8385 38390 10028 38392
rect 8385 38387 8451 38390
rect 9446 38366 10028 38390
rect 0 38178 800 38208
rect 1209 38178 1275 38181
rect 0 38176 1275 38178
rect 0 38120 1214 38176
rect 1270 38120 1275 38176
rect 0 38118 1275 38120
rect 0 38088 800 38118
rect 1209 38115 1275 38118
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 106654 38112 106970 38113
rect 106654 38048 106660 38112
rect 106724 38048 106740 38112
rect 106804 38048 106820 38112
rect 106884 38048 106900 38112
rect 106964 38048 106970 38112
rect 106654 38047 106970 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 105918 37568 106234 37569
rect 105918 37504 105924 37568
rect 105988 37504 106004 37568
rect 106068 37504 106084 37568
rect 106148 37504 106164 37568
rect 106228 37504 106234 37568
rect 105918 37503 106234 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 106654 37024 106970 37025
rect 106654 36960 106660 37024
rect 106724 36960 106740 37024
rect 106804 36960 106820 37024
rect 106884 36960 106900 37024
rect 106964 36960 106970 37024
rect 106654 36959 106970 36960
rect 0 36818 800 36848
rect 1393 36818 1459 36821
rect 0 36816 1459 36818
rect 0 36760 1398 36816
rect 1454 36760 1459 36816
rect 0 36758 1459 36760
rect 0 36728 800 36758
rect 1393 36755 1459 36758
rect 9489 36726 9555 36729
rect 9489 36724 10028 36726
rect 9489 36668 9494 36724
rect 9550 36668 10028 36724
rect 9489 36666 10028 36668
rect 9489 36663 9555 36666
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 105918 36480 106234 36481
rect 105918 36416 105924 36480
rect 105988 36416 106004 36480
rect 106068 36416 106084 36480
rect 106148 36416 106164 36480
rect 106228 36416 106234 36480
rect 105918 36415 106234 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 106654 35936 106970 35937
rect 106654 35872 106660 35936
rect 106724 35872 106740 35936
rect 106804 35872 106820 35936
rect 106884 35872 106900 35936
rect 106964 35872 106970 35936
rect 106654 35871 106970 35872
rect 9489 35643 9555 35646
rect 9489 35641 10028 35643
rect 9489 35585 9494 35641
rect 9550 35585 10028 35641
rect 9489 35583 10028 35585
rect 9489 35580 9555 35583
rect 0 35458 800 35488
rect 1301 35458 1367 35461
rect 0 35456 1367 35458
rect 0 35400 1306 35456
rect 1362 35400 1367 35456
rect 0 35398 1367 35400
rect 0 35368 800 35398
rect 1301 35395 1367 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 105918 35392 106234 35393
rect 105918 35328 105924 35392
rect 105988 35328 106004 35392
rect 106068 35328 106084 35392
rect 106148 35328 106164 35392
rect 106228 35328 106234 35392
rect 105918 35327 106234 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 106654 34848 106970 34849
rect 106654 34784 106660 34848
rect 106724 34784 106740 34848
rect 106804 34784 106820 34848
rect 106884 34784 106900 34848
rect 106964 34784 106970 34848
rect 106654 34783 106970 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 105918 34304 106234 34305
rect 105918 34240 105924 34304
rect 105988 34240 106004 34304
rect 106068 34240 106084 34304
rect 106148 34240 106164 34304
rect 106228 34240 106234 34304
rect 105918 34239 106234 34240
rect 0 34098 800 34128
rect 1393 34098 1459 34101
rect 0 34096 1459 34098
rect 0 34040 1398 34096
rect 1454 34040 1459 34096
rect 0 34038 1459 34040
rect 0 34008 800 34038
rect 1393 34035 1459 34038
rect 5533 33962 5599 33965
rect 9446 33962 10028 33963
rect 5533 33960 10028 33962
rect 5533 33904 5538 33960
rect 5594 33904 10028 33960
rect 5533 33903 10028 33904
rect 5533 33902 9506 33903
rect 5533 33899 5599 33902
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 106654 33760 106970 33761
rect 106654 33696 106660 33760
rect 106724 33696 106740 33760
rect 106804 33696 106820 33760
rect 106884 33696 106900 33760
rect 106964 33696 106970 33760
rect 106654 33695 106970 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 105918 33216 106234 33217
rect 105918 33152 105924 33216
rect 105988 33152 106004 33216
rect 106068 33152 106084 33216
rect 106148 33152 106164 33216
rect 106228 33152 106234 33216
rect 105918 33151 106234 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 106654 32672 106970 32673
rect 106654 32608 106660 32672
rect 106724 32608 106740 32672
rect 106804 32608 106820 32672
rect 106884 32608 106900 32672
rect 106964 32608 106970 32672
rect 106654 32607 106970 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 105918 32128 106234 32129
rect 105918 32064 105924 32128
rect 105988 32064 106004 32128
rect 106068 32064 106084 32128
rect 106148 32064 106164 32128
rect 106228 32064 106234 32128
rect 105918 32063 106234 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 106654 31584 106970 31585
rect 106654 31520 106660 31584
rect 106724 31520 106740 31584
rect 106804 31520 106820 31584
rect 106884 31520 106900 31584
rect 106964 31520 106970 31584
rect 106654 31519 106970 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 105918 31040 106234 31041
rect 105918 30976 105924 31040
rect 105988 30976 106004 31040
rect 106068 30976 106084 31040
rect 106148 30976 106164 31040
rect 106228 30976 106234 31040
rect 105918 30975 106234 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 106654 30496 106970 30497
rect 106654 30432 106660 30496
rect 106724 30432 106740 30496
rect 106804 30432 106820 30496
rect 106884 30432 106900 30496
rect 106964 30432 106970 30496
rect 106654 30431 106970 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 105918 29952 106234 29953
rect 105918 29888 105924 29952
rect 105988 29888 106004 29952
rect 106068 29888 106084 29952
rect 106148 29888 106164 29952
rect 106228 29888 106234 29952
rect 105918 29887 106234 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 106654 29408 106970 29409
rect 106654 29344 106660 29408
rect 106724 29344 106740 29408
rect 106804 29344 106820 29408
rect 106884 29344 106900 29408
rect 106964 29344 106970 29408
rect 106654 29343 106970 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 105918 28864 106234 28865
rect 105918 28800 105924 28864
rect 105988 28800 106004 28864
rect 106068 28800 106084 28864
rect 106148 28800 106164 28864
rect 106228 28800 106234 28864
rect 105918 28799 106234 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 106654 28320 106970 28321
rect 106654 28256 106660 28320
rect 106724 28256 106740 28320
rect 106804 28256 106820 28320
rect 106884 28256 106900 28320
rect 106964 28256 106970 28320
rect 106654 28255 106970 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 105918 27776 106234 27777
rect 105918 27712 105924 27776
rect 105988 27712 106004 27776
rect 106068 27712 106084 27776
rect 106148 27712 106164 27776
rect 106228 27712 106234 27776
rect 105918 27711 106234 27712
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 106654 27232 106970 27233
rect 106654 27168 106660 27232
rect 106724 27168 106740 27232
rect 106804 27168 106820 27232
rect 106884 27168 106900 27232
rect 106964 27168 106970 27232
rect 106654 27167 106970 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 105918 26688 106234 26689
rect 105918 26624 105924 26688
rect 105988 26624 106004 26688
rect 106068 26624 106084 26688
rect 106148 26624 106164 26688
rect 106228 26624 106234 26688
rect 105918 26623 106234 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 106654 26144 106970 26145
rect 106654 26080 106660 26144
rect 106724 26080 106740 26144
rect 106804 26080 106820 26144
rect 106884 26080 106900 26144
rect 106964 26080 106970 26144
rect 106654 26079 106970 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 105918 25600 106234 25601
rect 105918 25536 105924 25600
rect 105988 25536 106004 25600
rect 106068 25536 106084 25600
rect 106148 25536 106164 25600
rect 106228 25536 106234 25600
rect 105918 25535 106234 25536
rect 102593 25122 102659 25125
rect 102550 25120 102659 25122
rect 102317 25090 102383 25093
rect 102550 25090 102598 25120
rect 101948 25088 102598 25090
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 101948 25032 102322 25088
rect 102378 25064 102598 25088
rect 102654 25064 102659 25120
rect 102378 25059 102659 25064
rect 102378 25032 102610 25059
rect 101948 25030 102610 25032
rect 106654 25056 106970 25057
rect 102317 25027 102383 25030
rect 4870 24991 5186 24992
rect 106654 24992 106660 25056
rect 106724 24992 106740 25056
rect 106804 24992 106820 25056
rect 106884 24992 106900 25056
rect 106964 24992 106970 25056
rect 106654 24991 106970 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 105918 24512 106234 24513
rect 105918 24448 105924 24512
rect 105988 24448 106004 24512
rect 106068 24448 106084 24512
rect 106148 24448 106164 24512
rect 106228 24448 106234 24512
rect 105918 24447 106234 24448
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 106654 23968 106970 23969
rect 106654 23904 106660 23968
rect 106724 23904 106740 23968
rect 106804 23904 106820 23968
rect 106884 23904 106900 23968
rect 106964 23904 106970 23968
rect 106654 23903 106970 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 105918 23424 106234 23425
rect 102041 23390 102107 23393
rect 4210 23359 4526 23360
rect 101948 23388 102107 23390
rect 101948 23332 102046 23388
rect 102102 23332 102107 23388
rect 105918 23360 105924 23424
rect 105988 23360 106004 23424
rect 106068 23360 106084 23424
rect 106148 23360 106164 23424
rect 106228 23360 106234 23424
rect 105918 23359 106234 23360
rect 101948 23330 102107 23332
rect 102041 23327 102107 23330
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 106654 22880 106970 22881
rect 106654 22816 106660 22880
rect 106724 22816 106740 22880
rect 106804 22816 106820 22880
rect 106884 22816 106900 22880
rect 106964 22816 106970 22880
rect 106654 22815 106970 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 105918 22336 106234 22337
rect 105918 22272 105924 22336
rect 105988 22272 106004 22336
rect 106068 22272 106084 22336
rect 106148 22272 106164 22336
rect 106228 22272 106234 22336
rect 105918 22271 106234 22272
rect 104341 22266 104407 22269
rect 102550 22264 104407 22266
rect 102550 22262 104346 22264
rect 101948 22208 104346 22262
rect 104402 22208 104407 22264
rect 101948 22206 104407 22208
rect 101948 22202 102610 22206
rect 104341 22203 104407 22206
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 106654 21792 106970 21793
rect 106654 21728 106660 21792
rect 106724 21728 106740 21792
rect 106804 21728 106820 21792
rect 106884 21728 106900 21792
rect 106964 21728 106970 21792
rect 106654 21727 106970 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 105918 21248 106234 21249
rect 105918 21184 105924 21248
rect 105988 21184 106004 21248
rect 106068 21184 106084 21248
rect 106148 21184 106164 21248
rect 106228 21184 106234 21248
rect 105918 21183 106234 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 106654 20704 106970 20705
rect 106654 20640 106660 20704
rect 106724 20640 106740 20704
rect 106804 20640 106820 20704
rect 106884 20640 106900 20704
rect 106964 20640 106970 20704
rect 106654 20639 106970 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 105918 20160 106234 20161
rect 105918 20096 105924 20160
rect 105988 20096 106004 20160
rect 106068 20096 106084 20160
rect 106148 20096 106164 20160
rect 106228 20096 106234 20160
rect 105918 20095 106234 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 106654 19616 106970 19617
rect 106654 19552 106660 19616
rect 106724 19552 106740 19616
rect 106804 19552 106820 19616
rect 106884 19552 106900 19616
rect 106964 19552 106970 19616
rect 106654 19551 106970 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 105918 19072 106234 19073
rect 105918 19008 105924 19072
rect 105988 19008 106004 19072
rect 106068 19008 106084 19072
rect 106148 19008 106164 19072
rect 106228 19008 106234 19072
rect 105918 19007 106234 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 106654 18528 106970 18529
rect 106654 18464 106660 18528
rect 106724 18464 106740 18528
rect 106804 18464 106820 18528
rect 106884 18464 106900 18528
rect 106964 18464 106970 18528
rect 106654 18463 106970 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 105918 17984 106234 17985
rect 105918 17920 105924 17984
rect 105988 17920 106004 17984
rect 106068 17920 106084 17984
rect 106148 17920 106164 17984
rect 106228 17920 106234 17984
rect 105918 17919 106234 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 106654 17440 106970 17441
rect 106654 17376 106660 17440
rect 106724 17376 106740 17440
rect 106804 17376 106820 17440
rect 106884 17376 106900 17440
rect 106964 17376 106970 17440
rect 106654 17375 106970 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 105918 16896 106234 16897
rect 105918 16832 105924 16896
rect 105988 16832 106004 16896
rect 106068 16832 106084 16896
rect 106148 16832 106164 16896
rect 106228 16832 106234 16896
rect 105918 16831 106234 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 106654 16352 106970 16353
rect 106654 16288 106660 16352
rect 106724 16288 106740 16352
rect 106804 16288 106820 16352
rect 106884 16288 106900 16352
rect 106964 16288 106970 16352
rect 106654 16287 106970 16288
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 105918 15808 106234 15809
rect 105918 15744 105924 15808
rect 105988 15744 106004 15808
rect 106068 15744 106084 15808
rect 106148 15744 106164 15808
rect 106228 15744 106234 15808
rect 105918 15743 106234 15744
rect 1301 15738 1367 15741
rect 0 15736 1367 15738
rect 0 15680 1306 15736
rect 1362 15680 1367 15736
rect 0 15678 1367 15680
rect 0 15648 800 15678
rect 1301 15675 1367 15678
rect 9489 15483 9555 15486
rect 9489 15481 10028 15483
rect 9489 15425 9494 15481
rect 9550 15425 10028 15481
rect 9489 15423 10028 15425
rect 9489 15420 9555 15423
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 106654 15264 106970 15265
rect 106654 15200 106660 15264
rect 106724 15200 106740 15264
rect 106804 15200 106820 15264
rect 106884 15200 106900 15264
rect 106964 15200 106970 15264
rect 106654 15199 106970 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 105918 14720 106234 14721
rect 105918 14656 105924 14720
rect 105988 14656 106004 14720
rect 106068 14656 106084 14720
rect 106148 14656 106164 14720
rect 106228 14656 106234 14720
rect 105918 14655 106234 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 106654 14176 106970 14177
rect 106654 14112 106660 14176
rect 106724 14112 106740 14176
rect 106804 14112 106820 14176
rect 106884 14112 106900 14176
rect 106964 14112 106970 14176
rect 106654 14111 106970 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 105918 13632 106234 13633
rect 105918 13568 105924 13632
rect 105988 13568 106004 13632
rect 106068 13568 106084 13632
rect 106148 13568 106164 13632
rect 106228 13568 106234 13632
rect 105918 13567 106234 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 106654 13088 106970 13089
rect 106654 13024 106660 13088
rect 106724 13024 106740 13088
rect 106804 13024 106820 13088
rect 106884 13024 106900 13088
rect 106964 13024 106970 13088
rect 106654 13023 106970 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 105918 12544 106234 12545
rect 105918 12480 105924 12544
rect 105988 12480 106004 12544
rect 106068 12480 106084 12544
rect 106148 12480 106164 12544
rect 106228 12480 106234 12544
rect 105918 12479 106234 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 106654 12000 106970 12001
rect 106654 11936 106660 12000
rect 106724 11936 106740 12000
rect 106804 11936 106820 12000
rect 106884 11936 106900 12000
rect 106964 11936 106970 12000
rect 106654 11935 106970 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 105918 11456 106234 11457
rect 105918 11392 105924 11456
rect 105988 11392 106004 11456
rect 106068 11392 106084 11456
rect 106148 11392 106164 11456
rect 106228 11392 106234 11456
rect 105918 11391 106234 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 106654 10912 106970 10913
rect 106654 10848 106660 10912
rect 106724 10848 106740 10912
rect 106804 10848 106820 10912
rect 106884 10848 106900 10912
rect 106964 10848 106970 10912
rect 106654 10847 106970 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 105918 10368 106234 10369
rect 105918 10304 105924 10368
rect 105988 10304 106004 10368
rect 106068 10304 106084 10368
rect 106148 10304 106164 10368
rect 106228 10304 106234 10368
rect 105918 10303 106234 10304
rect 9581 9890 9647 9893
rect 16113 9892 16179 9893
rect 16052 9890 16058 9892
rect 9581 9888 16058 9890
rect 16122 9890 16179 9892
rect 16122 9888 16250 9890
rect 9581 9832 9586 9888
rect 9642 9832 16058 9888
rect 16174 9832 16250 9888
rect 9581 9830 16058 9832
rect 9581 9827 9647 9830
rect 16052 9828 16058 9830
rect 16122 9830 16250 9832
rect 16122 9828 16179 9830
rect 90521 9828 90527 9892
rect 90591 9890 90597 9892
rect 90817 9890 90883 9893
rect 90591 9888 90883 9890
rect 90591 9832 90822 9888
rect 90878 9832 90883 9888
rect 90591 9830 90883 9832
rect 90591 9828 90597 9830
rect 16113 9827 16179 9828
rect 90817 9827 90883 9830
rect 90950 9828 90956 9892
rect 91020 9890 91026 9892
rect 104801 9890 104867 9893
rect 91020 9888 104867 9890
rect 91020 9832 104806 9888
rect 104862 9832 104867 9888
rect 91020 9830 104867 9832
rect 91020 9828 91026 9830
rect 104801 9827 104867 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 106654 9824 106970 9825
rect 106654 9760 106660 9824
rect 106724 9760 106740 9824
rect 106804 9760 106820 9824
rect 106884 9760 106900 9824
rect 106964 9760 106970 9824
rect 106654 9759 106970 9760
rect 90725 9756 90791 9757
rect 90674 9754 90680 9756
rect 90634 9694 90680 9754
rect 90744 9752 90791 9756
rect 90786 9696 90791 9752
rect 90674 9692 90680 9694
rect 90744 9692 90791 9696
rect 90725 9691 90791 9692
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 105918 9280 106234 9281
rect 105918 9216 105924 9280
rect 105988 9216 106004 9280
rect 106068 9216 106084 9280
rect 106148 9216 106164 9280
rect 106228 9216 106234 9280
rect 105918 9215 106234 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 106654 8736 106970 8737
rect 106654 8672 106660 8736
rect 106724 8672 106740 8736
rect 106804 8672 106820 8736
rect 106884 8672 106900 8736
rect 106964 8672 106970 8736
rect 106654 8671 106970 8672
rect 23473 8260 23539 8261
rect 24761 8260 24827 8261
rect 25865 8260 25931 8261
rect 23422 8258 23428 8260
rect 23382 8198 23428 8258
rect 23492 8256 23539 8260
rect 23534 8200 23539 8256
rect 23422 8196 23428 8198
rect 23492 8196 23539 8200
rect 24710 8196 24716 8260
rect 24780 8258 24827 8260
rect 25814 8258 25820 8260
rect 24780 8256 24872 8258
rect 24822 8200 24872 8256
rect 24780 8198 24872 8200
rect 25774 8198 25820 8258
rect 25884 8256 25931 8260
rect 25926 8200 25931 8256
rect 24780 8196 24827 8198
rect 25814 8196 25820 8198
rect 25884 8196 25931 8200
rect 26918 8196 26924 8260
rect 26988 8258 26994 8260
rect 27153 8258 27219 8261
rect 26988 8256 27219 8258
rect 26988 8200 27158 8256
rect 27214 8200 27219 8256
rect 26988 8198 27219 8200
rect 26988 8196 26994 8198
rect 23473 8195 23539 8196
rect 24761 8195 24827 8196
rect 25865 8195 25931 8196
rect 27153 8195 27219 8198
rect 28206 8196 28212 8260
rect 28276 8258 28282 8260
rect 28441 8258 28507 8261
rect 28276 8256 28507 8258
rect 28276 8200 28446 8256
rect 28502 8200 28507 8256
rect 28276 8198 28507 8200
rect 28276 8196 28282 8198
rect 28441 8195 28507 8198
rect 29269 8260 29335 8261
rect 29269 8256 29316 8260
rect 29380 8258 29386 8260
rect 29269 8200 29274 8256
rect 29269 8196 29316 8200
rect 29380 8198 29426 8258
rect 29380 8196 29386 8198
rect 30414 8196 30420 8260
rect 30484 8258 30490 8260
rect 30557 8258 30623 8261
rect 31661 8260 31727 8261
rect 31661 8258 31708 8260
rect 30484 8256 30623 8258
rect 30484 8200 30562 8256
rect 30618 8200 30623 8256
rect 30484 8198 30623 8200
rect 31616 8256 31708 8258
rect 31616 8200 31666 8256
rect 31616 8198 31708 8200
rect 30484 8196 30490 8198
rect 29269 8195 29335 8196
rect 30557 8195 30623 8198
rect 31661 8196 31708 8198
rect 31772 8196 31778 8260
rect 32806 8196 32812 8260
rect 32876 8258 32882 8260
rect 32949 8258 33015 8261
rect 32876 8256 33015 8258
rect 32876 8200 32954 8256
rect 33010 8200 33015 8256
rect 32876 8198 33015 8200
rect 32876 8196 32882 8198
rect 31661 8195 31727 8196
rect 32949 8195 33015 8198
rect 33910 8196 33916 8260
rect 33980 8258 33986 8260
rect 34237 8258 34303 8261
rect 33980 8256 34303 8258
rect 33980 8200 34242 8256
rect 34298 8200 34303 8256
rect 33980 8198 34303 8200
rect 33980 8196 33986 8198
rect 34237 8195 34303 8198
rect 35198 8196 35204 8260
rect 35268 8258 35274 8260
rect 35433 8258 35499 8261
rect 36353 8260 36419 8261
rect 37457 8260 37523 8261
rect 38745 8260 38811 8261
rect 36302 8258 36308 8260
rect 35268 8256 35499 8258
rect 35268 8200 35438 8256
rect 35494 8200 35499 8256
rect 35268 8198 35499 8200
rect 36262 8198 36308 8258
rect 36372 8256 36419 8260
rect 37406 8258 37412 8260
rect 36414 8200 36419 8256
rect 35268 8196 35274 8198
rect 35433 8195 35499 8198
rect 36302 8196 36308 8198
rect 36372 8196 36419 8200
rect 37366 8198 37412 8258
rect 37476 8256 37523 8260
rect 38694 8258 38700 8260
rect 37518 8200 37523 8256
rect 37406 8196 37412 8198
rect 37476 8196 37523 8200
rect 38654 8198 38700 8258
rect 38764 8256 38811 8260
rect 38806 8200 38811 8256
rect 38694 8196 38700 8198
rect 38764 8196 38811 8200
rect 40902 8196 40908 8260
rect 40972 8258 40978 8260
rect 41321 8258 41387 8261
rect 40972 8256 41387 8258
rect 40972 8200 41326 8256
rect 41382 8200 41387 8256
rect 40972 8198 41387 8200
rect 40972 8196 40978 8198
rect 36353 8195 36419 8196
rect 37457 8195 37523 8196
rect 38745 8195 38811 8196
rect 41321 8195 41387 8198
rect 42149 8260 42215 8261
rect 42149 8256 42196 8260
rect 42260 8258 42266 8260
rect 42149 8200 42154 8256
rect 42149 8196 42196 8200
rect 42260 8198 42306 8258
rect 42260 8196 42266 8198
rect 43294 8196 43300 8260
rect 43364 8258 43370 8260
rect 43437 8258 43503 8261
rect 90633 8260 90699 8261
rect 91001 8260 91067 8261
rect 90582 8258 90588 8260
rect 43364 8256 43503 8258
rect 43364 8200 43442 8256
rect 43498 8200 43503 8256
rect 43364 8198 43503 8200
rect 90542 8198 90588 8258
rect 90652 8256 90699 8260
rect 90950 8258 90956 8260
rect 90694 8200 90699 8256
rect 43364 8196 43370 8198
rect 42149 8195 42215 8196
rect 43437 8195 43503 8198
rect 90582 8196 90588 8198
rect 90652 8196 90699 8200
rect 90910 8198 90956 8258
rect 91020 8256 91067 8260
rect 91062 8200 91067 8256
rect 90950 8196 90956 8198
rect 91020 8196 91067 8200
rect 90633 8195 90699 8196
rect 91001 8195 91067 8196
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 105918 8192 106234 8193
rect 105918 8128 105924 8192
rect 105988 8128 106004 8192
rect 106068 8128 106084 8192
rect 106148 8128 106164 8192
rect 106228 8128 106234 8192
rect 105918 8127 106234 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 66310 7648 66626 7649
rect 66310 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66626 7648
rect 66310 7583 66626 7584
rect 97030 7648 97346 7649
rect 97030 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97346 7648
rect 97030 7583 97346 7584
rect 106654 7648 106970 7649
rect 106654 7584 106660 7648
rect 106724 7584 106740 7648
rect 106804 7584 106820 7648
rect 106884 7584 106900 7648
rect 106964 7584 106970 7648
rect 106654 7583 106970 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 96370 7104 96686 7105
rect 96370 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96686 7104
rect 96370 7039 96686 7040
rect 105918 7104 106234 7105
rect 105918 7040 105924 7104
rect 105988 7040 106004 7104
rect 106068 7040 106084 7104
rect 106148 7040 106164 7104
rect 106228 7040 106234 7104
rect 105918 7039 106234 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 66310 6560 66626 6561
rect 66310 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66626 6560
rect 66310 6495 66626 6496
rect 97030 6560 97346 6561
rect 97030 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97346 6560
rect 97030 6495 97346 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 96370 6016 96686 6017
rect 96370 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96686 6016
rect 96370 5951 96686 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 66310 5472 66626 5473
rect 66310 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66626 5472
rect 66310 5407 66626 5408
rect 97030 5472 97346 5473
rect 97030 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97346 5472
rect 97030 5407 97346 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 96370 4928 96686 4929
rect 96370 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96686 4928
rect 96370 4863 96686 4864
rect 39798 4524 39804 4588
rect 39868 4586 39874 4588
rect 39941 4586 40007 4589
rect 39868 4584 40007 4586
rect 39868 4528 39946 4584
rect 40002 4528 40007 4584
rect 39868 4526 40007 4528
rect 39868 4524 39874 4526
rect 39941 4523 40007 4526
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 66310 4384 66626 4385
rect 66310 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66626 4384
rect 66310 4319 66626 4320
rect 97030 4384 97346 4385
rect 97030 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97346 4384
rect 97030 4319 97346 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 96370 3840 96686 3841
rect 96370 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96686 3840
rect 96370 3775 96686 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 66310 3296 66626 3297
rect 66310 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66626 3296
rect 66310 3231 66626 3232
rect 97030 3296 97346 3297
rect 97030 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97346 3296
rect 97030 3231 97346 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 96370 2752 96686 2753
rect 96370 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96686 2752
rect 96370 2687 96686 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 66310 2208 66626 2209
rect 66310 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66626 2208
rect 66310 2143 66626 2144
rect 97030 2208 97346 2209
rect 97030 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97346 2208
rect 97030 2143 97346 2144
<< via3 >>
rect 4876 127324 4940 127328
rect 4876 127268 4880 127324
rect 4880 127268 4936 127324
rect 4936 127268 4940 127324
rect 4876 127264 4940 127268
rect 4956 127324 5020 127328
rect 4956 127268 4960 127324
rect 4960 127268 5016 127324
rect 5016 127268 5020 127324
rect 4956 127264 5020 127268
rect 5036 127324 5100 127328
rect 5036 127268 5040 127324
rect 5040 127268 5096 127324
rect 5096 127268 5100 127324
rect 5036 127264 5100 127268
rect 5116 127324 5180 127328
rect 5116 127268 5120 127324
rect 5120 127268 5176 127324
rect 5176 127268 5180 127324
rect 5116 127264 5180 127268
rect 35596 127324 35660 127328
rect 35596 127268 35600 127324
rect 35600 127268 35656 127324
rect 35656 127268 35660 127324
rect 35596 127264 35660 127268
rect 35676 127324 35740 127328
rect 35676 127268 35680 127324
rect 35680 127268 35736 127324
rect 35736 127268 35740 127324
rect 35676 127264 35740 127268
rect 35756 127324 35820 127328
rect 35756 127268 35760 127324
rect 35760 127268 35816 127324
rect 35816 127268 35820 127324
rect 35756 127264 35820 127268
rect 35836 127324 35900 127328
rect 35836 127268 35840 127324
rect 35840 127268 35896 127324
rect 35896 127268 35900 127324
rect 35836 127264 35900 127268
rect 66316 127324 66380 127328
rect 66316 127268 66320 127324
rect 66320 127268 66376 127324
rect 66376 127268 66380 127324
rect 66316 127264 66380 127268
rect 66396 127324 66460 127328
rect 66396 127268 66400 127324
rect 66400 127268 66456 127324
rect 66456 127268 66460 127324
rect 66396 127264 66460 127268
rect 66476 127324 66540 127328
rect 66476 127268 66480 127324
rect 66480 127268 66536 127324
rect 66536 127268 66540 127324
rect 66476 127264 66540 127268
rect 66556 127324 66620 127328
rect 66556 127268 66560 127324
rect 66560 127268 66616 127324
rect 66616 127268 66620 127324
rect 66556 127264 66620 127268
rect 97036 127324 97100 127328
rect 97036 127268 97040 127324
rect 97040 127268 97096 127324
rect 97096 127268 97100 127324
rect 97036 127264 97100 127268
rect 97116 127324 97180 127328
rect 97116 127268 97120 127324
rect 97120 127268 97176 127324
rect 97176 127268 97180 127324
rect 97116 127264 97180 127268
rect 97196 127324 97260 127328
rect 97196 127268 97200 127324
rect 97200 127268 97256 127324
rect 97256 127268 97260 127324
rect 97196 127264 97260 127268
rect 97276 127324 97340 127328
rect 97276 127268 97280 127324
rect 97280 127268 97336 127324
rect 97336 127268 97340 127324
rect 97276 127264 97340 127268
rect 4216 126780 4280 126784
rect 4216 126724 4220 126780
rect 4220 126724 4276 126780
rect 4276 126724 4280 126780
rect 4216 126720 4280 126724
rect 4296 126780 4360 126784
rect 4296 126724 4300 126780
rect 4300 126724 4356 126780
rect 4356 126724 4360 126780
rect 4296 126720 4360 126724
rect 4376 126780 4440 126784
rect 4376 126724 4380 126780
rect 4380 126724 4436 126780
rect 4436 126724 4440 126780
rect 4376 126720 4440 126724
rect 4456 126780 4520 126784
rect 4456 126724 4460 126780
rect 4460 126724 4516 126780
rect 4516 126724 4520 126780
rect 4456 126720 4520 126724
rect 34936 126780 35000 126784
rect 34936 126724 34940 126780
rect 34940 126724 34996 126780
rect 34996 126724 35000 126780
rect 34936 126720 35000 126724
rect 35016 126780 35080 126784
rect 35016 126724 35020 126780
rect 35020 126724 35076 126780
rect 35076 126724 35080 126780
rect 35016 126720 35080 126724
rect 35096 126780 35160 126784
rect 35096 126724 35100 126780
rect 35100 126724 35156 126780
rect 35156 126724 35160 126780
rect 35096 126720 35160 126724
rect 35176 126780 35240 126784
rect 35176 126724 35180 126780
rect 35180 126724 35236 126780
rect 35236 126724 35240 126780
rect 35176 126720 35240 126724
rect 65656 126780 65720 126784
rect 65656 126724 65660 126780
rect 65660 126724 65716 126780
rect 65716 126724 65720 126780
rect 65656 126720 65720 126724
rect 65736 126780 65800 126784
rect 65736 126724 65740 126780
rect 65740 126724 65796 126780
rect 65796 126724 65800 126780
rect 65736 126720 65800 126724
rect 65816 126780 65880 126784
rect 65816 126724 65820 126780
rect 65820 126724 65876 126780
rect 65876 126724 65880 126780
rect 65816 126720 65880 126724
rect 65896 126780 65960 126784
rect 65896 126724 65900 126780
rect 65900 126724 65956 126780
rect 65956 126724 65960 126780
rect 65896 126720 65960 126724
rect 96376 126780 96440 126784
rect 96376 126724 96380 126780
rect 96380 126724 96436 126780
rect 96436 126724 96440 126780
rect 96376 126720 96440 126724
rect 96456 126780 96520 126784
rect 96456 126724 96460 126780
rect 96460 126724 96516 126780
rect 96516 126724 96520 126780
rect 96456 126720 96520 126724
rect 96536 126780 96600 126784
rect 96536 126724 96540 126780
rect 96540 126724 96596 126780
rect 96596 126724 96600 126780
rect 96536 126720 96600 126724
rect 96616 126780 96680 126784
rect 96616 126724 96620 126780
rect 96620 126724 96676 126780
rect 96676 126724 96680 126780
rect 96616 126720 96680 126724
rect 105924 126780 105988 126784
rect 105924 126724 105928 126780
rect 105928 126724 105984 126780
rect 105984 126724 105988 126780
rect 105924 126720 105988 126724
rect 106004 126780 106068 126784
rect 106004 126724 106008 126780
rect 106008 126724 106064 126780
rect 106064 126724 106068 126780
rect 106004 126720 106068 126724
rect 106084 126780 106148 126784
rect 106084 126724 106088 126780
rect 106088 126724 106144 126780
rect 106144 126724 106148 126780
rect 106084 126720 106148 126724
rect 106164 126780 106228 126784
rect 106164 126724 106168 126780
rect 106168 126724 106224 126780
rect 106224 126724 106228 126780
rect 106164 126720 106228 126724
rect 73476 126380 73540 126444
rect 4876 126236 4940 126240
rect 4876 126180 4880 126236
rect 4880 126180 4936 126236
rect 4936 126180 4940 126236
rect 4876 126176 4940 126180
rect 4956 126236 5020 126240
rect 4956 126180 4960 126236
rect 4960 126180 5016 126236
rect 5016 126180 5020 126236
rect 4956 126176 5020 126180
rect 5036 126236 5100 126240
rect 5036 126180 5040 126236
rect 5040 126180 5096 126236
rect 5096 126180 5100 126236
rect 5036 126176 5100 126180
rect 5116 126236 5180 126240
rect 5116 126180 5120 126236
rect 5120 126180 5176 126236
rect 5176 126180 5180 126236
rect 5116 126176 5180 126180
rect 35596 126236 35660 126240
rect 35596 126180 35600 126236
rect 35600 126180 35656 126236
rect 35656 126180 35660 126236
rect 35596 126176 35660 126180
rect 35676 126236 35740 126240
rect 35676 126180 35680 126236
rect 35680 126180 35736 126236
rect 35736 126180 35740 126236
rect 35676 126176 35740 126180
rect 35756 126236 35820 126240
rect 35756 126180 35760 126236
rect 35760 126180 35816 126236
rect 35816 126180 35820 126236
rect 35756 126176 35820 126180
rect 35836 126236 35900 126240
rect 35836 126180 35840 126236
rect 35840 126180 35896 126236
rect 35896 126180 35900 126236
rect 35836 126176 35900 126180
rect 66316 126236 66380 126240
rect 66316 126180 66320 126236
rect 66320 126180 66376 126236
rect 66376 126180 66380 126236
rect 66316 126176 66380 126180
rect 66396 126236 66460 126240
rect 66396 126180 66400 126236
rect 66400 126180 66456 126236
rect 66456 126180 66460 126236
rect 66396 126176 66460 126180
rect 66476 126236 66540 126240
rect 66476 126180 66480 126236
rect 66480 126180 66536 126236
rect 66536 126180 66540 126236
rect 66476 126176 66540 126180
rect 66556 126236 66620 126240
rect 66556 126180 66560 126236
rect 66560 126180 66616 126236
rect 66616 126180 66620 126236
rect 66556 126176 66620 126180
rect 97036 126236 97100 126240
rect 97036 126180 97040 126236
rect 97040 126180 97096 126236
rect 97096 126180 97100 126236
rect 97036 126176 97100 126180
rect 97116 126236 97180 126240
rect 97116 126180 97120 126236
rect 97120 126180 97176 126236
rect 97176 126180 97180 126236
rect 97116 126176 97180 126180
rect 97196 126236 97260 126240
rect 97196 126180 97200 126236
rect 97200 126180 97256 126236
rect 97256 126180 97260 126236
rect 97196 126176 97260 126180
rect 97276 126236 97340 126240
rect 97276 126180 97280 126236
rect 97280 126180 97336 126236
rect 97336 126180 97340 126236
rect 97276 126176 97340 126180
rect 106660 126236 106724 126240
rect 106660 126180 106664 126236
rect 106664 126180 106720 126236
rect 106720 126180 106724 126236
rect 106660 126176 106724 126180
rect 106740 126236 106804 126240
rect 106740 126180 106744 126236
rect 106744 126180 106800 126236
rect 106800 126180 106804 126236
rect 106740 126176 106804 126180
rect 106820 126236 106884 126240
rect 106820 126180 106824 126236
rect 106824 126180 106880 126236
rect 106880 126180 106884 126236
rect 106820 126176 106884 126180
rect 106900 126236 106964 126240
rect 106900 126180 106904 126236
rect 106904 126180 106960 126236
rect 106960 126180 106964 126236
rect 106900 126176 106964 126180
rect 46060 125972 46124 126036
rect 53604 125972 53668 126036
rect 58572 125700 58636 125764
rect 4216 125692 4280 125696
rect 4216 125636 4220 125692
rect 4220 125636 4276 125692
rect 4276 125636 4280 125692
rect 4216 125632 4280 125636
rect 4296 125692 4360 125696
rect 4296 125636 4300 125692
rect 4300 125636 4356 125692
rect 4356 125636 4360 125692
rect 4296 125632 4360 125636
rect 4376 125692 4440 125696
rect 4376 125636 4380 125692
rect 4380 125636 4436 125692
rect 4436 125636 4440 125692
rect 4376 125632 4440 125636
rect 4456 125692 4520 125696
rect 4456 125636 4460 125692
rect 4460 125636 4516 125692
rect 4516 125636 4520 125692
rect 4456 125632 4520 125636
rect 105924 125692 105988 125696
rect 105924 125636 105928 125692
rect 105928 125636 105984 125692
rect 105984 125636 105988 125692
rect 105924 125632 105988 125636
rect 106004 125692 106068 125696
rect 106004 125636 106008 125692
rect 106008 125636 106064 125692
rect 106064 125636 106068 125692
rect 106004 125632 106068 125636
rect 106084 125692 106148 125696
rect 106084 125636 106088 125692
rect 106088 125636 106144 125692
rect 106144 125636 106148 125692
rect 106084 125632 106148 125636
rect 106164 125692 106228 125696
rect 106164 125636 106168 125692
rect 106168 125636 106224 125692
rect 106224 125636 106228 125692
rect 106164 125632 106228 125636
rect 51028 125564 51092 125628
rect 55996 125564 56060 125628
rect 61148 125564 61212 125628
rect 63540 125156 63604 125220
rect 4876 125148 4940 125152
rect 4876 125092 4880 125148
rect 4880 125092 4936 125148
rect 4936 125092 4940 125148
rect 4876 125088 4940 125092
rect 4956 125148 5020 125152
rect 4956 125092 4960 125148
rect 4960 125092 5016 125148
rect 5016 125092 5020 125148
rect 4956 125088 5020 125092
rect 5036 125148 5100 125152
rect 5036 125092 5040 125148
rect 5040 125092 5096 125148
rect 5096 125092 5100 125148
rect 5036 125088 5100 125092
rect 5116 125148 5180 125152
rect 5116 125092 5120 125148
rect 5120 125092 5176 125148
rect 5176 125092 5180 125148
rect 5116 125088 5180 125092
rect 106660 125148 106724 125152
rect 106660 125092 106664 125148
rect 106664 125092 106720 125148
rect 106720 125092 106724 125148
rect 106660 125088 106724 125092
rect 106740 125148 106804 125152
rect 106740 125092 106744 125148
rect 106744 125092 106800 125148
rect 106800 125092 106804 125148
rect 106740 125088 106804 125092
rect 106820 125148 106884 125152
rect 106820 125092 106824 125148
rect 106824 125092 106880 125148
rect 106880 125092 106884 125148
rect 106820 125088 106884 125092
rect 106900 125148 106964 125152
rect 106900 125092 106904 125148
rect 106904 125092 106960 125148
rect 106960 125092 106964 125148
rect 106900 125088 106964 125092
rect 4216 124604 4280 124608
rect 4216 124548 4220 124604
rect 4220 124548 4276 124604
rect 4276 124548 4280 124604
rect 4216 124544 4280 124548
rect 4296 124604 4360 124608
rect 4296 124548 4300 124604
rect 4300 124548 4356 124604
rect 4356 124548 4360 124604
rect 4296 124544 4360 124548
rect 4376 124604 4440 124608
rect 4376 124548 4380 124604
rect 4380 124548 4436 124604
rect 4436 124548 4440 124604
rect 4376 124544 4440 124548
rect 4456 124604 4520 124608
rect 4456 124548 4460 124604
rect 4460 124548 4516 124604
rect 4516 124548 4520 124604
rect 4456 124544 4520 124548
rect 105924 124604 105988 124608
rect 105924 124548 105928 124604
rect 105928 124548 105984 124604
rect 105984 124548 105988 124604
rect 105924 124544 105988 124548
rect 106004 124604 106068 124608
rect 106004 124548 106008 124604
rect 106008 124548 106064 124604
rect 106064 124548 106068 124604
rect 106004 124544 106068 124548
rect 106084 124604 106148 124608
rect 106084 124548 106088 124604
rect 106088 124548 106144 124604
rect 106144 124548 106148 124604
rect 106084 124544 106148 124548
rect 106164 124604 106228 124608
rect 106164 124548 106168 124604
rect 106168 124548 106224 124604
rect 106224 124548 106228 124604
rect 106164 124544 106228 124548
rect 36075 124264 36139 124268
rect 36075 124208 36082 124264
rect 36082 124208 36138 124264
rect 36138 124208 36139 124264
rect 36075 124204 36139 124208
rect 38571 124204 38635 124268
rect 41067 124204 41131 124268
rect 48544 124264 48608 124268
rect 48544 124208 48558 124264
rect 48558 124208 48608 124264
rect 48544 124204 48608 124208
rect 66027 124264 66091 124268
rect 66027 124208 66074 124264
rect 66074 124208 66091 124264
rect 66027 124204 66091 124208
rect 68523 124264 68587 124268
rect 68523 124208 68558 124264
rect 68558 124208 68587 124264
rect 68523 124204 68587 124208
rect 71019 124204 71083 124268
rect 43563 124068 43627 124132
rect 4876 124060 4940 124064
rect 4876 124004 4880 124060
rect 4880 124004 4936 124060
rect 4936 124004 4940 124060
rect 4876 124000 4940 124004
rect 4956 124060 5020 124064
rect 4956 124004 4960 124060
rect 4960 124004 5016 124060
rect 5016 124004 5020 124060
rect 4956 124000 5020 124004
rect 5036 124060 5100 124064
rect 5036 124004 5040 124060
rect 5040 124004 5096 124060
rect 5096 124004 5100 124060
rect 5036 124000 5100 124004
rect 5116 124060 5180 124064
rect 5116 124004 5120 124060
rect 5120 124004 5176 124060
rect 5176 124004 5180 124060
rect 5116 124000 5180 124004
rect 106660 124060 106724 124064
rect 106660 124004 106664 124060
rect 106664 124004 106720 124060
rect 106720 124004 106724 124060
rect 106660 124000 106724 124004
rect 106740 124060 106804 124064
rect 106740 124004 106744 124060
rect 106744 124004 106800 124060
rect 106800 124004 106804 124060
rect 106740 124000 106804 124004
rect 106820 124060 106884 124064
rect 106820 124004 106824 124060
rect 106824 124004 106880 124060
rect 106880 124004 106884 124060
rect 106820 124000 106884 124004
rect 106900 124060 106964 124064
rect 106900 124004 106904 124060
rect 106904 124004 106960 124060
rect 106960 124004 106964 124060
rect 106900 124000 106964 124004
rect 86142 123932 86206 123996
rect 87310 123856 87374 123860
rect 87310 123800 87326 123856
rect 87326 123800 87374 123856
rect 87310 123796 87374 123800
rect 96108 123856 96172 123860
rect 96108 123800 96122 123856
rect 96122 123800 96172 123856
rect 96108 123796 96172 123800
rect 4216 123516 4280 123520
rect 4216 123460 4220 123516
rect 4220 123460 4276 123516
rect 4276 123460 4280 123516
rect 4216 123456 4280 123460
rect 4296 123516 4360 123520
rect 4296 123460 4300 123516
rect 4300 123460 4356 123516
rect 4356 123460 4360 123516
rect 4296 123456 4360 123460
rect 4376 123516 4440 123520
rect 4376 123460 4380 123516
rect 4380 123460 4436 123516
rect 4436 123460 4440 123516
rect 4376 123456 4440 123460
rect 4456 123516 4520 123520
rect 4456 123460 4460 123516
rect 4460 123460 4516 123516
rect 4516 123460 4520 123516
rect 4456 123456 4520 123460
rect 105924 123516 105988 123520
rect 105924 123460 105928 123516
rect 105928 123460 105984 123516
rect 105984 123460 105988 123516
rect 105924 123456 105988 123460
rect 106004 123516 106068 123520
rect 106004 123460 106008 123516
rect 106008 123460 106064 123516
rect 106064 123460 106068 123516
rect 106004 123456 106068 123460
rect 106084 123516 106148 123520
rect 106084 123460 106088 123516
rect 106088 123460 106144 123516
rect 106144 123460 106148 123516
rect 106084 123456 106148 123460
rect 106164 123516 106228 123520
rect 106164 123460 106168 123516
rect 106168 123460 106224 123516
rect 106224 123460 106228 123516
rect 106164 123456 106228 123460
rect 4876 122972 4940 122976
rect 4876 122916 4880 122972
rect 4880 122916 4936 122972
rect 4936 122916 4940 122972
rect 4876 122912 4940 122916
rect 4956 122972 5020 122976
rect 4956 122916 4960 122972
rect 4960 122916 5016 122972
rect 5016 122916 5020 122972
rect 4956 122912 5020 122916
rect 5036 122972 5100 122976
rect 5036 122916 5040 122972
rect 5040 122916 5096 122972
rect 5096 122916 5100 122972
rect 5036 122912 5100 122916
rect 5116 122972 5180 122976
rect 5116 122916 5120 122972
rect 5120 122916 5176 122972
rect 5176 122916 5180 122972
rect 5116 122912 5180 122916
rect 106660 122972 106724 122976
rect 106660 122916 106664 122972
rect 106664 122916 106720 122972
rect 106720 122916 106724 122972
rect 106660 122912 106724 122916
rect 106740 122972 106804 122976
rect 106740 122916 106744 122972
rect 106744 122916 106800 122972
rect 106800 122916 106804 122972
rect 106740 122912 106804 122916
rect 106820 122972 106884 122976
rect 106820 122916 106824 122972
rect 106824 122916 106880 122972
rect 106880 122916 106884 122972
rect 106820 122912 106884 122916
rect 106900 122972 106964 122976
rect 106900 122916 106904 122972
rect 106904 122916 106960 122972
rect 106960 122916 106964 122972
rect 106900 122912 106964 122916
rect 4216 122428 4280 122432
rect 4216 122372 4220 122428
rect 4220 122372 4276 122428
rect 4276 122372 4280 122428
rect 4216 122368 4280 122372
rect 4296 122428 4360 122432
rect 4296 122372 4300 122428
rect 4300 122372 4356 122428
rect 4356 122372 4360 122428
rect 4296 122368 4360 122372
rect 4376 122428 4440 122432
rect 4376 122372 4380 122428
rect 4380 122372 4436 122428
rect 4436 122372 4440 122428
rect 4376 122368 4440 122372
rect 4456 122428 4520 122432
rect 4456 122372 4460 122428
rect 4460 122372 4516 122428
rect 4516 122372 4520 122428
rect 4456 122368 4520 122372
rect 105924 122428 105988 122432
rect 105924 122372 105928 122428
rect 105928 122372 105984 122428
rect 105984 122372 105988 122428
rect 105924 122368 105988 122372
rect 106004 122428 106068 122432
rect 106004 122372 106008 122428
rect 106008 122372 106064 122428
rect 106064 122372 106068 122428
rect 106004 122368 106068 122372
rect 106084 122428 106148 122432
rect 106084 122372 106088 122428
rect 106088 122372 106144 122428
rect 106144 122372 106148 122428
rect 106084 122368 106148 122372
rect 106164 122428 106228 122432
rect 106164 122372 106168 122428
rect 106168 122372 106224 122428
rect 106224 122372 106228 122428
rect 106164 122368 106228 122372
rect 4876 121884 4940 121888
rect 4876 121828 4880 121884
rect 4880 121828 4936 121884
rect 4936 121828 4940 121884
rect 4876 121824 4940 121828
rect 4956 121884 5020 121888
rect 4956 121828 4960 121884
rect 4960 121828 5016 121884
rect 5016 121828 5020 121884
rect 4956 121824 5020 121828
rect 5036 121884 5100 121888
rect 5036 121828 5040 121884
rect 5040 121828 5096 121884
rect 5096 121828 5100 121884
rect 5036 121824 5100 121828
rect 5116 121884 5180 121888
rect 5116 121828 5120 121884
rect 5120 121828 5176 121884
rect 5176 121828 5180 121884
rect 5116 121824 5180 121828
rect 106660 121884 106724 121888
rect 106660 121828 106664 121884
rect 106664 121828 106720 121884
rect 106720 121828 106724 121884
rect 106660 121824 106724 121828
rect 106740 121884 106804 121888
rect 106740 121828 106744 121884
rect 106744 121828 106800 121884
rect 106800 121828 106804 121884
rect 106740 121824 106804 121828
rect 106820 121884 106884 121888
rect 106820 121828 106824 121884
rect 106824 121828 106880 121884
rect 106880 121828 106884 121884
rect 106820 121824 106884 121828
rect 106900 121884 106964 121888
rect 106900 121828 106904 121884
rect 106904 121828 106960 121884
rect 106960 121828 106964 121884
rect 106900 121824 106964 121828
rect 4216 121340 4280 121344
rect 4216 121284 4220 121340
rect 4220 121284 4276 121340
rect 4276 121284 4280 121340
rect 4216 121280 4280 121284
rect 4296 121340 4360 121344
rect 4296 121284 4300 121340
rect 4300 121284 4356 121340
rect 4356 121284 4360 121340
rect 4296 121280 4360 121284
rect 4376 121340 4440 121344
rect 4376 121284 4380 121340
rect 4380 121284 4436 121340
rect 4436 121284 4440 121340
rect 4376 121280 4440 121284
rect 4456 121340 4520 121344
rect 4456 121284 4460 121340
rect 4460 121284 4516 121340
rect 4516 121284 4520 121340
rect 4456 121280 4520 121284
rect 105924 121340 105988 121344
rect 105924 121284 105928 121340
rect 105928 121284 105984 121340
rect 105984 121284 105988 121340
rect 105924 121280 105988 121284
rect 106004 121340 106068 121344
rect 106004 121284 106008 121340
rect 106008 121284 106064 121340
rect 106064 121284 106068 121340
rect 106004 121280 106068 121284
rect 106084 121340 106148 121344
rect 106084 121284 106088 121340
rect 106088 121284 106144 121340
rect 106144 121284 106148 121340
rect 106084 121280 106148 121284
rect 106164 121340 106228 121344
rect 106164 121284 106168 121340
rect 106168 121284 106224 121340
rect 106224 121284 106228 121340
rect 106164 121280 106228 121284
rect 4876 120796 4940 120800
rect 4876 120740 4880 120796
rect 4880 120740 4936 120796
rect 4936 120740 4940 120796
rect 4876 120736 4940 120740
rect 4956 120796 5020 120800
rect 4956 120740 4960 120796
rect 4960 120740 5016 120796
rect 5016 120740 5020 120796
rect 4956 120736 5020 120740
rect 5036 120796 5100 120800
rect 5036 120740 5040 120796
rect 5040 120740 5096 120796
rect 5096 120740 5100 120796
rect 5036 120736 5100 120740
rect 5116 120796 5180 120800
rect 5116 120740 5120 120796
rect 5120 120740 5176 120796
rect 5176 120740 5180 120796
rect 5116 120736 5180 120740
rect 106660 120796 106724 120800
rect 106660 120740 106664 120796
rect 106664 120740 106720 120796
rect 106720 120740 106724 120796
rect 106660 120736 106724 120740
rect 106740 120796 106804 120800
rect 106740 120740 106744 120796
rect 106744 120740 106800 120796
rect 106800 120740 106804 120796
rect 106740 120736 106804 120740
rect 106820 120796 106884 120800
rect 106820 120740 106824 120796
rect 106824 120740 106880 120796
rect 106880 120740 106884 120796
rect 106820 120736 106884 120740
rect 106900 120796 106964 120800
rect 106900 120740 106904 120796
rect 106904 120740 106960 120796
rect 106960 120740 106964 120796
rect 106900 120736 106964 120740
rect 4216 120252 4280 120256
rect 4216 120196 4220 120252
rect 4220 120196 4276 120252
rect 4276 120196 4280 120252
rect 4216 120192 4280 120196
rect 4296 120252 4360 120256
rect 4296 120196 4300 120252
rect 4300 120196 4356 120252
rect 4356 120196 4360 120252
rect 4296 120192 4360 120196
rect 4376 120252 4440 120256
rect 4376 120196 4380 120252
rect 4380 120196 4436 120252
rect 4436 120196 4440 120252
rect 4376 120192 4440 120196
rect 4456 120252 4520 120256
rect 4456 120196 4460 120252
rect 4460 120196 4516 120252
rect 4516 120196 4520 120252
rect 4456 120192 4520 120196
rect 105924 120252 105988 120256
rect 105924 120196 105928 120252
rect 105928 120196 105984 120252
rect 105984 120196 105988 120252
rect 105924 120192 105988 120196
rect 106004 120252 106068 120256
rect 106004 120196 106008 120252
rect 106008 120196 106064 120252
rect 106064 120196 106068 120252
rect 106004 120192 106068 120196
rect 106084 120252 106148 120256
rect 106084 120196 106088 120252
rect 106088 120196 106144 120252
rect 106144 120196 106148 120252
rect 106084 120192 106148 120196
rect 106164 120252 106228 120256
rect 106164 120196 106168 120252
rect 106168 120196 106224 120252
rect 106224 120196 106228 120252
rect 106164 120192 106228 120196
rect 4876 119708 4940 119712
rect 4876 119652 4880 119708
rect 4880 119652 4936 119708
rect 4936 119652 4940 119708
rect 4876 119648 4940 119652
rect 4956 119708 5020 119712
rect 4956 119652 4960 119708
rect 4960 119652 5016 119708
rect 5016 119652 5020 119708
rect 4956 119648 5020 119652
rect 5036 119708 5100 119712
rect 5036 119652 5040 119708
rect 5040 119652 5096 119708
rect 5096 119652 5100 119708
rect 5036 119648 5100 119652
rect 5116 119708 5180 119712
rect 5116 119652 5120 119708
rect 5120 119652 5176 119708
rect 5176 119652 5180 119708
rect 5116 119648 5180 119652
rect 106660 119708 106724 119712
rect 106660 119652 106664 119708
rect 106664 119652 106720 119708
rect 106720 119652 106724 119708
rect 106660 119648 106724 119652
rect 106740 119708 106804 119712
rect 106740 119652 106744 119708
rect 106744 119652 106800 119708
rect 106800 119652 106804 119708
rect 106740 119648 106804 119652
rect 106820 119708 106884 119712
rect 106820 119652 106824 119708
rect 106824 119652 106880 119708
rect 106880 119652 106884 119708
rect 106820 119648 106884 119652
rect 106900 119708 106964 119712
rect 106900 119652 106904 119708
rect 106904 119652 106960 119708
rect 106960 119652 106964 119708
rect 106900 119648 106964 119652
rect 4216 119164 4280 119168
rect 4216 119108 4220 119164
rect 4220 119108 4276 119164
rect 4276 119108 4280 119164
rect 4216 119104 4280 119108
rect 4296 119164 4360 119168
rect 4296 119108 4300 119164
rect 4300 119108 4356 119164
rect 4356 119108 4360 119164
rect 4296 119104 4360 119108
rect 4376 119164 4440 119168
rect 4376 119108 4380 119164
rect 4380 119108 4436 119164
rect 4436 119108 4440 119164
rect 4376 119104 4440 119108
rect 4456 119164 4520 119168
rect 4456 119108 4460 119164
rect 4460 119108 4516 119164
rect 4516 119108 4520 119164
rect 4456 119104 4520 119108
rect 105924 119164 105988 119168
rect 105924 119108 105928 119164
rect 105928 119108 105984 119164
rect 105984 119108 105988 119164
rect 105924 119104 105988 119108
rect 106004 119164 106068 119168
rect 106004 119108 106008 119164
rect 106008 119108 106064 119164
rect 106064 119108 106068 119164
rect 106004 119104 106068 119108
rect 106084 119164 106148 119168
rect 106084 119108 106088 119164
rect 106088 119108 106144 119164
rect 106144 119108 106148 119164
rect 106084 119104 106148 119108
rect 106164 119164 106228 119168
rect 106164 119108 106168 119164
rect 106168 119108 106224 119164
rect 106224 119108 106228 119164
rect 106164 119104 106228 119108
rect 4876 118620 4940 118624
rect 4876 118564 4880 118620
rect 4880 118564 4936 118620
rect 4936 118564 4940 118620
rect 4876 118560 4940 118564
rect 4956 118620 5020 118624
rect 4956 118564 4960 118620
rect 4960 118564 5016 118620
rect 5016 118564 5020 118620
rect 4956 118560 5020 118564
rect 5036 118620 5100 118624
rect 5036 118564 5040 118620
rect 5040 118564 5096 118620
rect 5096 118564 5100 118620
rect 5036 118560 5100 118564
rect 5116 118620 5180 118624
rect 5116 118564 5120 118620
rect 5120 118564 5176 118620
rect 5176 118564 5180 118620
rect 5116 118560 5180 118564
rect 106660 118620 106724 118624
rect 106660 118564 106664 118620
rect 106664 118564 106720 118620
rect 106720 118564 106724 118620
rect 106660 118560 106724 118564
rect 106740 118620 106804 118624
rect 106740 118564 106744 118620
rect 106744 118564 106800 118620
rect 106800 118564 106804 118620
rect 106740 118560 106804 118564
rect 106820 118620 106884 118624
rect 106820 118564 106824 118620
rect 106824 118564 106880 118620
rect 106880 118564 106884 118620
rect 106820 118560 106884 118564
rect 106900 118620 106964 118624
rect 106900 118564 106904 118620
rect 106904 118564 106960 118620
rect 106960 118564 106964 118620
rect 106900 118560 106964 118564
rect 4216 118076 4280 118080
rect 4216 118020 4220 118076
rect 4220 118020 4276 118076
rect 4276 118020 4280 118076
rect 4216 118016 4280 118020
rect 4296 118076 4360 118080
rect 4296 118020 4300 118076
rect 4300 118020 4356 118076
rect 4356 118020 4360 118076
rect 4296 118016 4360 118020
rect 4376 118076 4440 118080
rect 4376 118020 4380 118076
rect 4380 118020 4436 118076
rect 4436 118020 4440 118076
rect 4376 118016 4440 118020
rect 4456 118076 4520 118080
rect 4456 118020 4460 118076
rect 4460 118020 4516 118076
rect 4516 118020 4520 118076
rect 4456 118016 4520 118020
rect 105924 118076 105988 118080
rect 105924 118020 105928 118076
rect 105928 118020 105984 118076
rect 105984 118020 105988 118076
rect 105924 118016 105988 118020
rect 106004 118076 106068 118080
rect 106004 118020 106008 118076
rect 106008 118020 106064 118076
rect 106064 118020 106068 118076
rect 106004 118016 106068 118020
rect 106084 118076 106148 118080
rect 106084 118020 106088 118076
rect 106088 118020 106144 118076
rect 106144 118020 106148 118076
rect 106084 118016 106148 118020
rect 106164 118076 106228 118080
rect 106164 118020 106168 118076
rect 106168 118020 106224 118076
rect 106224 118020 106228 118076
rect 106164 118016 106228 118020
rect 4876 117532 4940 117536
rect 4876 117476 4880 117532
rect 4880 117476 4936 117532
rect 4936 117476 4940 117532
rect 4876 117472 4940 117476
rect 4956 117532 5020 117536
rect 4956 117476 4960 117532
rect 4960 117476 5016 117532
rect 5016 117476 5020 117532
rect 4956 117472 5020 117476
rect 5036 117532 5100 117536
rect 5036 117476 5040 117532
rect 5040 117476 5096 117532
rect 5096 117476 5100 117532
rect 5036 117472 5100 117476
rect 5116 117532 5180 117536
rect 5116 117476 5120 117532
rect 5120 117476 5176 117532
rect 5176 117476 5180 117532
rect 5116 117472 5180 117476
rect 106660 117532 106724 117536
rect 106660 117476 106664 117532
rect 106664 117476 106720 117532
rect 106720 117476 106724 117532
rect 106660 117472 106724 117476
rect 106740 117532 106804 117536
rect 106740 117476 106744 117532
rect 106744 117476 106800 117532
rect 106800 117476 106804 117532
rect 106740 117472 106804 117476
rect 106820 117532 106884 117536
rect 106820 117476 106824 117532
rect 106824 117476 106880 117532
rect 106880 117476 106884 117532
rect 106820 117472 106884 117476
rect 106900 117532 106964 117536
rect 106900 117476 106904 117532
rect 106904 117476 106960 117532
rect 106960 117476 106964 117532
rect 106900 117472 106964 117476
rect 4216 116988 4280 116992
rect 4216 116932 4220 116988
rect 4220 116932 4276 116988
rect 4276 116932 4280 116988
rect 4216 116928 4280 116932
rect 4296 116988 4360 116992
rect 4296 116932 4300 116988
rect 4300 116932 4356 116988
rect 4356 116932 4360 116988
rect 4296 116928 4360 116932
rect 4376 116988 4440 116992
rect 4376 116932 4380 116988
rect 4380 116932 4436 116988
rect 4436 116932 4440 116988
rect 4376 116928 4440 116932
rect 4456 116988 4520 116992
rect 4456 116932 4460 116988
rect 4460 116932 4516 116988
rect 4516 116932 4520 116988
rect 4456 116928 4520 116932
rect 105924 116988 105988 116992
rect 105924 116932 105928 116988
rect 105928 116932 105984 116988
rect 105984 116932 105988 116988
rect 105924 116928 105988 116932
rect 106004 116988 106068 116992
rect 106004 116932 106008 116988
rect 106008 116932 106064 116988
rect 106064 116932 106068 116988
rect 106004 116928 106068 116932
rect 106084 116988 106148 116992
rect 106084 116932 106088 116988
rect 106088 116932 106144 116988
rect 106144 116932 106148 116988
rect 106084 116928 106148 116932
rect 106164 116988 106228 116992
rect 106164 116932 106168 116988
rect 106168 116932 106224 116988
rect 106224 116932 106228 116988
rect 106164 116928 106228 116932
rect 4876 116444 4940 116448
rect 4876 116388 4880 116444
rect 4880 116388 4936 116444
rect 4936 116388 4940 116444
rect 4876 116384 4940 116388
rect 4956 116444 5020 116448
rect 4956 116388 4960 116444
rect 4960 116388 5016 116444
rect 5016 116388 5020 116444
rect 4956 116384 5020 116388
rect 5036 116444 5100 116448
rect 5036 116388 5040 116444
rect 5040 116388 5096 116444
rect 5096 116388 5100 116444
rect 5036 116384 5100 116388
rect 5116 116444 5180 116448
rect 5116 116388 5120 116444
rect 5120 116388 5176 116444
rect 5176 116388 5180 116444
rect 5116 116384 5180 116388
rect 106660 116444 106724 116448
rect 106660 116388 106664 116444
rect 106664 116388 106720 116444
rect 106720 116388 106724 116444
rect 106660 116384 106724 116388
rect 106740 116444 106804 116448
rect 106740 116388 106744 116444
rect 106744 116388 106800 116444
rect 106800 116388 106804 116444
rect 106740 116384 106804 116388
rect 106820 116444 106884 116448
rect 106820 116388 106824 116444
rect 106824 116388 106880 116444
rect 106880 116388 106884 116444
rect 106820 116384 106884 116388
rect 106900 116444 106964 116448
rect 106900 116388 106904 116444
rect 106904 116388 106960 116444
rect 106960 116388 106964 116444
rect 106900 116384 106964 116388
rect 4216 115900 4280 115904
rect 4216 115844 4220 115900
rect 4220 115844 4276 115900
rect 4276 115844 4280 115900
rect 4216 115840 4280 115844
rect 4296 115900 4360 115904
rect 4296 115844 4300 115900
rect 4300 115844 4356 115900
rect 4356 115844 4360 115900
rect 4296 115840 4360 115844
rect 4376 115900 4440 115904
rect 4376 115844 4380 115900
rect 4380 115844 4436 115900
rect 4436 115844 4440 115900
rect 4376 115840 4440 115844
rect 4456 115900 4520 115904
rect 4456 115844 4460 115900
rect 4460 115844 4516 115900
rect 4516 115844 4520 115900
rect 4456 115840 4520 115844
rect 105924 115900 105988 115904
rect 105924 115844 105928 115900
rect 105928 115844 105984 115900
rect 105984 115844 105988 115900
rect 105924 115840 105988 115844
rect 106004 115900 106068 115904
rect 106004 115844 106008 115900
rect 106008 115844 106064 115900
rect 106064 115844 106068 115900
rect 106004 115840 106068 115844
rect 106084 115900 106148 115904
rect 106084 115844 106088 115900
rect 106088 115844 106144 115900
rect 106144 115844 106148 115900
rect 106084 115840 106148 115844
rect 106164 115900 106228 115904
rect 106164 115844 106168 115900
rect 106168 115844 106224 115900
rect 106224 115844 106228 115900
rect 106164 115840 106228 115844
rect 4876 115356 4940 115360
rect 4876 115300 4880 115356
rect 4880 115300 4936 115356
rect 4936 115300 4940 115356
rect 4876 115296 4940 115300
rect 4956 115356 5020 115360
rect 4956 115300 4960 115356
rect 4960 115300 5016 115356
rect 5016 115300 5020 115356
rect 4956 115296 5020 115300
rect 5036 115356 5100 115360
rect 5036 115300 5040 115356
rect 5040 115300 5096 115356
rect 5096 115300 5100 115356
rect 5036 115296 5100 115300
rect 5116 115356 5180 115360
rect 5116 115300 5120 115356
rect 5120 115300 5176 115356
rect 5176 115300 5180 115356
rect 5116 115296 5180 115300
rect 106660 115356 106724 115360
rect 106660 115300 106664 115356
rect 106664 115300 106720 115356
rect 106720 115300 106724 115356
rect 106660 115296 106724 115300
rect 106740 115356 106804 115360
rect 106740 115300 106744 115356
rect 106744 115300 106800 115356
rect 106800 115300 106804 115356
rect 106740 115296 106804 115300
rect 106820 115356 106884 115360
rect 106820 115300 106824 115356
rect 106824 115300 106880 115356
rect 106880 115300 106884 115356
rect 106820 115296 106884 115300
rect 106900 115356 106964 115360
rect 106900 115300 106904 115356
rect 106904 115300 106960 115356
rect 106960 115300 106964 115356
rect 106900 115296 106964 115300
rect 4216 114812 4280 114816
rect 4216 114756 4220 114812
rect 4220 114756 4276 114812
rect 4276 114756 4280 114812
rect 4216 114752 4280 114756
rect 4296 114812 4360 114816
rect 4296 114756 4300 114812
rect 4300 114756 4356 114812
rect 4356 114756 4360 114812
rect 4296 114752 4360 114756
rect 4376 114812 4440 114816
rect 4376 114756 4380 114812
rect 4380 114756 4436 114812
rect 4436 114756 4440 114812
rect 4376 114752 4440 114756
rect 4456 114812 4520 114816
rect 4456 114756 4460 114812
rect 4460 114756 4516 114812
rect 4516 114756 4520 114812
rect 4456 114752 4520 114756
rect 105924 114812 105988 114816
rect 105924 114756 105928 114812
rect 105928 114756 105984 114812
rect 105984 114756 105988 114812
rect 105924 114752 105988 114756
rect 106004 114812 106068 114816
rect 106004 114756 106008 114812
rect 106008 114756 106064 114812
rect 106064 114756 106068 114812
rect 106004 114752 106068 114756
rect 106084 114812 106148 114816
rect 106084 114756 106088 114812
rect 106088 114756 106144 114812
rect 106144 114756 106148 114812
rect 106084 114752 106148 114756
rect 106164 114812 106228 114816
rect 106164 114756 106168 114812
rect 106168 114756 106224 114812
rect 106224 114756 106228 114812
rect 106164 114752 106228 114756
rect 4876 114268 4940 114272
rect 4876 114212 4880 114268
rect 4880 114212 4936 114268
rect 4936 114212 4940 114268
rect 4876 114208 4940 114212
rect 4956 114268 5020 114272
rect 4956 114212 4960 114268
rect 4960 114212 5016 114268
rect 5016 114212 5020 114268
rect 4956 114208 5020 114212
rect 5036 114268 5100 114272
rect 5036 114212 5040 114268
rect 5040 114212 5096 114268
rect 5096 114212 5100 114268
rect 5036 114208 5100 114212
rect 5116 114268 5180 114272
rect 5116 114212 5120 114268
rect 5120 114212 5176 114268
rect 5176 114212 5180 114268
rect 5116 114208 5180 114212
rect 106660 114268 106724 114272
rect 106660 114212 106664 114268
rect 106664 114212 106720 114268
rect 106720 114212 106724 114268
rect 106660 114208 106724 114212
rect 106740 114268 106804 114272
rect 106740 114212 106744 114268
rect 106744 114212 106800 114268
rect 106800 114212 106804 114268
rect 106740 114208 106804 114212
rect 106820 114268 106884 114272
rect 106820 114212 106824 114268
rect 106824 114212 106880 114268
rect 106880 114212 106884 114268
rect 106820 114208 106884 114212
rect 106900 114268 106964 114272
rect 106900 114212 106904 114268
rect 106904 114212 106960 114268
rect 106960 114212 106964 114268
rect 106900 114208 106964 114212
rect 4216 113724 4280 113728
rect 4216 113668 4220 113724
rect 4220 113668 4276 113724
rect 4276 113668 4280 113724
rect 4216 113664 4280 113668
rect 4296 113724 4360 113728
rect 4296 113668 4300 113724
rect 4300 113668 4356 113724
rect 4356 113668 4360 113724
rect 4296 113664 4360 113668
rect 4376 113724 4440 113728
rect 4376 113668 4380 113724
rect 4380 113668 4436 113724
rect 4436 113668 4440 113724
rect 4376 113664 4440 113668
rect 4456 113724 4520 113728
rect 4456 113668 4460 113724
rect 4460 113668 4516 113724
rect 4516 113668 4520 113724
rect 4456 113664 4520 113668
rect 105924 113724 105988 113728
rect 105924 113668 105928 113724
rect 105928 113668 105984 113724
rect 105984 113668 105988 113724
rect 105924 113664 105988 113668
rect 106004 113724 106068 113728
rect 106004 113668 106008 113724
rect 106008 113668 106064 113724
rect 106064 113668 106068 113724
rect 106004 113664 106068 113668
rect 106084 113724 106148 113728
rect 106084 113668 106088 113724
rect 106088 113668 106144 113724
rect 106144 113668 106148 113724
rect 106084 113664 106148 113668
rect 106164 113724 106228 113728
rect 106164 113668 106168 113724
rect 106168 113668 106224 113724
rect 106224 113668 106228 113724
rect 106164 113664 106228 113668
rect 4876 113180 4940 113184
rect 4876 113124 4880 113180
rect 4880 113124 4936 113180
rect 4936 113124 4940 113180
rect 4876 113120 4940 113124
rect 4956 113180 5020 113184
rect 4956 113124 4960 113180
rect 4960 113124 5016 113180
rect 5016 113124 5020 113180
rect 4956 113120 5020 113124
rect 5036 113180 5100 113184
rect 5036 113124 5040 113180
rect 5040 113124 5096 113180
rect 5096 113124 5100 113180
rect 5036 113120 5100 113124
rect 5116 113180 5180 113184
rect 5116 113124 5120 113180
rect 5120 113124 5176 113180
rect 5176 113124 5180 113180
rect 5116 113120 5180 113124
rect 106660 113180 106724 113184
rect 106660 113124 106664 113180
rect 106664 113124 106720 113180
rect 106720 113124 106724 113180
rect 106660 113120 106724 113124
rect 106740 113180 106804 113184
rect 106740 113124 106744 113180
rect 106744 113124 106800 113180
rect 106800 113124 106804 113180
rect 106740 113120 106804 113124
rect 106820 113180 106884 113184
rect 106820 113124 106824 113180
rect 106824 113124 106880 113180
rect 106880 113124 106884 113180
rect 106820 113120 106884 113124
rect 106900 113180 106964 113184
rect 106900 113124 106904 113180
rect 106904 113124 106960 113180
rect 106960 113124 106964 113180
rect 106900 113120 106964 113124
rect 4216 112636 4280 112640
rect 4216 112580 4220 112636
rect 4220 112580 4276 112636
rect 4276 112580 4280 112636
rect 4216 112576 4280 112580
rect 4296 112636 4360 112640
rect 4296 112580 4300 112636
rect 4300 112580 4356 112636
rect 4356 112580 4360 112636
rect 4296 112576 4360 112580
rect 4376 112636 4440 112640
rect 4376 112580 4380 112636
rect 4380 112580 4436 112636
rect 4436 112580 4440 112636
rect 4376 112576 4440 112580
rect 4456 112636 4520 112640
rect 4456 112580 4460 112636
rect 4460 112580 4516 112636
rect 4516 112580 4520 112636
rect 4456 112576 4520 112580
rect 105924 112636 105988 112640
rect 105924 112580 105928 112636
rect 105928 112580 105984 112636
rect 105984 112580 105988 112636
rect 105924 112576 105988 112580
rect 106004 112636 106068 112640
rect 106004 112580 106008 112636
rect 106008 112580 106064 112636
rect 106064 112580 106068 112636
rect 106004 112576 106068 112580
rect 106084 112636 106148 112640
rect 106084 112580 106088 112636
rect 106088 112580 106144 112636
rect 106144 112580 106148 112636
rect 106084 112576 106148 112580
rect 106164 112636 106228 112640
rect 106164 112580 106168 112636
rect 106168 112580 106224 112636
rect 106224 112580 106228 112636
rect 106164 112576 106228 112580
rect 4876 112092 4940 112096
rect 4876 112036 4880 112092
rect 4880 112036 4936 112092
rect 4936 112036 4940 112092
rect 4876 112032 4940 112036
rect 4956 112092 5020 112096
rect 4956 112036 4960 112092
rect 4960 112036 5016 112092
rect 5016 112036 5020 112092
rect 4956 112032 5020 112036
rect 5036 112092 5100 112096
rect 5036 112036 5040 112092
rect 5040 112036 5096 112092
rect 5096 112036 5100 112092
rect 5036 112032 5100 112036
rect 5116 112092 5180 112096
rect 5116 112036 5120 112092
rect 5120 112036 5176 112092
rect 5176 112036 5180 112092
rect 5116 112032 5180 112036
rect 106660 112092 106724 112096
rect 106660 112036 106664 112092
rect 106664 112036 106720 112092
rect 106720 112036 106724 112092
rect 106660 112032 106724 112036
rect 106740 112092 106804 112096
rect 106740 112036 106744 112092
rect 106744 112036 106800 112092
rect 106800 112036 106804 112092
rect 106740 112032 106804 112036
rect 106820 112092 106884 112096
rect 106820 112036 106824 112092
rect 106824 112036 106880 112092
rect 106880 112036 106884 112092
rect 106820 112032 106884 112036
rect 106900 112092 106964 112096
rect 106900 112036 106904 112092
rect 106904 112036 106960 112092
rect 106960 112036 106964 112092
rect 106900 112032 106964 112036
rect 4216 111548 4280 111552
rect 4216 111492 4220 111548
rect 4220 111492 4276 111548
rect 4276 111492 4280 111548
rect 4216 111488 4280 111492
rect 4296 111548 4360 111552
rect 4296 111492 4300 111548
rect 4300 111492 4356 111548
rect 4356 111492 4360 111548
rect 4296 111488 4360 111492
rect 4376 111548 4440 111552
rect 4376 111492 4380 111548
rect 4380 111492 4436 111548
rect 4436 111492 4440 111548
rect 4376 111488 4440 111492
rect 4456 111548 4520 111552
rect 4456 111492 4460 111548
rect 4460 111492 4516 111548
rect 4516 111492 4520 111548
rect 4456 111488 4520 111492
rect 105924 111548 105988 111552
rect 105924 111492 105928 111548
rect 105928 111492 105984 111548
rect 105984 111492 105988 111548
rect 105924 111488 105988 111492
rect 106004 111548 106068 111552
rect 106004 111492 106008 111548
rect 106008 111492 106064 111548
rect 106064 111492 106068 111548
rect 106004 111488 106068 111492
rect 106084 111548 106148 111552
rect 106084 111492 106088 111548
rect 106088 111492 106144 111548
rect 106144 111492 106148 111548
rect 106084 111488 106148 111492
rect 106164 111548 106228 111552
rect 106164 111492 106168 111548
rect 106168 111492 106224 111548
rect 106224 111492 106228 111548
rect 106164 111488 106228 111492
rect 4876 111004 4940 111008
rect 4876 110948 4880 111004
rect 4880 110948 4936 111004
rect 4936 110948 4940 111004
rect 4876 110944 4940 110948
rect 4956 111004 5020 111008
rect 4956 110948 4960 111004
rect 4960 110948 5016 111004
rect 5016 110948 5020 111004
rect 4956 110944 5020 110948
rect 5036 111004 5100 111008
rect 5036 110948 5040 111004
rect 5040 110948 5096 111004
rect 5096 110948 5100 111004
rect 5036 110944 5100 110948
rect 5116 111004 5180 111008
rect 5116 110948 5120 111004
rect 5120 110948 5176 111004
rect 5176 110948 5180 111004
rect 5116 110944 5180 110948
rect 106660 111004 106724 111008
rect 106660 110948 106664 111004
rect 106664 110948 106720 111004
rect 106720 110948 106724 111004
rect 106660 110944 106724 110948
rect 106740 111004 106804 111008
rect 106740 110948 106744 111004
rect 106744 110948 106800 111004
rect 106800 110948 106804 111004
rect 106740 110944 106804 110948
rect 106820 111004 106884 111008
rect 106820 110948 106824 111004
rect 106824 110948 106880 111004
rect 106880 110948 106884 111004
rect 106820 110944 106884 110948
rect 106900 111004 106964 111008
rect 106900 110948 106904 111004
rect 106904 110948 106960 111004
rect 106960 110948 106964 111004
rect 106900 110944 106964 110948
rect 4216 110460 4280 110464
rect 4216 110404 4220 110460
rect 4220 110404 4276 110460
rect 4276 110404 4280 110460
rect 4216 110400 4280 110404
rect 4296 110460 4360 110464
rect 4296 110404 4300 110460
rect 4300 110404 4356 110460
rect 4356 110404 4360 110460
rect 4296 110400 4360 110404
rect 4376 110460 4440 110464
rect 4376 110404 4380 110460
rect 4380 110404 4436 110460
rect 4436 110404 4440 110460
rect 4376 110400 4440 110404
rect 4456 110460 4520 110464
rect 4456 110404 4460 110460
rect 4460 110404 4516 110460
rect 4516 110404 4520 110460
rect 4456 110400 4520 110404
rect 105924 110460 105988 110464
rect 105924 110404 105928 110460
rect 105928 110404 105984 110460
rect 105984 110404 105988 110460
rect 105924 110400 105988 110404
rect 106004 110460 106068 110464
rect 106004 110404 106008 110460
rect 106008 110404 106064 110460
rect 106064 110404 106068 110460
rect 106004 110400 106068 110404
rect 106084 110460 106148 110464
rect 106084 110404 106088 110460
rect 106088 110404 106144 110460
rect 106144 110404 106148 110460
rect 106084 110400 106148 110404
rect 106164 110460 106228 110464
rect 106164 110404 106168 110460
rect 106168 110404 106224 110460
rect 106224 110404 106228 110460
rect 106164 110400 106228 110404
rect 4876 109916 4940 109920
rect 4876 109860 4880 109916
rect 4880 109860 4936 109916
rect 4936 109860 4940 109916
rect 4876 109856 4940 109860
rect 4956 109916 5020 109920
rect 4956 109860 4960 109916
rect 4960 109860 5016 109916
rect 5016 109860 5020 109916
rect 4956 109856 5020 109860
rect 5036 109916 5100 109920
rect 5036 109860 5040 109916
rect 5040 109860 5096 109916
rect 5096 109860 5100 109916
rect 5036 109856 5100 109860
rect 5116 109916 5180 109920
rect 5116 109860 5120 109916
rect 5120 109860 5176 109916
rect 5176 109860 5180 109916
rect 5116 109856 5180 109860
rect 106660 109916 106724 109920
rect 106660 109860 106664 109916
rect 106664 109860 106720 109916
rect 106720 109860 106724 109916
rect 106660 109856 106724 109860
rect 106740 109916 106804 109920
rect 106740 109860 106744 109916
rect 106744 109860 106800 109916
rect 106800 109860 106804 109916
rect 106740 109856 106804 109860
rect 106820 109916 106884 109920
rect 106820 109860 106824 109916
rect 106824 109860 106880 109916
rect 106880 109860 106884 109916
rect 106820 109856 106884 109860
rect 106900 109916 106964 109920
rect 106900 109860 106904 109916
rect 106904 109860 106960 109916
rect 106960 109860 106964 109916
rect 106900 109856 106964 109860
rect 4216 109372 4280 109376
rect 4216 109316 4220 109372
rect 4220 109316 4276 109372
rect 4276 109316 4280 109372
rect 4216 109312 4280 109316
rect 4296 109372 4360 109376
rect 4296 109316 4300 109372
rect 4300 109316 4356 109372
rect 4356 109316 4360 109372
rect 4296 109312 4360 109316
rect 4376 109372 4440 109376
rect 4376 109316 4380 109372
rect 4380 109316 4436 109372
rect 4436 109316 4440 109372
rect 4376 109312 4440 109316
rect 4456 109372 4520 109376
rect 4456 109316 4460 109372
rect 4460 109316 4516 109372
rect 4516 109316 4520 109372
rect 4456 109312 4520 109316
rect 105924 109372 105988 109376
rect 105924 109316 105928 109372
rect 105928 109316 105984 109372
rect 105984 109316 105988 109372
rect 105924 109312 105988 109316
rect 106004 109372 106068 109376
rect 106004 109316 106008 109372
rect 106008 109316 106064 109372
rect 106064 109316 106068 109372
rect 106004 109312 106068 109316
rect 106084 109372 106148 109376
rect 106084 109316 106088 109372
rect 106088 109316 106144 109372
rect 106144 109316 106148 109372
rect 106084 109312 106148 109316
rect 106164 109372 106228 109376
rect 106164 109316 106168 109372
rect 106168 109316 106224 109372
rect 106224 109316 106228 109372
rect 106164 109312 106228 109316
rect 4876 108828 4940 108832
rect 4876 108772 4880 108828
rect 4880 108772 4936 108828
rect 4936 108772 4940 108828
rect 4876 108768 4940 108772
rect 4956 108828 5020 108832
rect 4956 108772 4960 108828
rect 4960 108772 5016 108828
rect 5016 108772 5020 108828
rect 4956 108768 5020 108772
rect 5036 108828 5100 108832
rect 5036 108772 5040 108828
rect 5040 108772 5096 108828
rect 5096 108772 5100 108828
rect 5036 108768 5100 108772
rect 5116 108828 5180 108832
rect 5116 108772 5120 108828
rect 5120 108772 5176 108828
rect 5176 108772 5180 108828
rect 5116 108768 5180 108772
rect 106660 108828 106724 108832
rect 106660 108772 106664 108828
rect 106664 108772 106720 108828
rect 106720 108772 106724 108828
rect 106660 108768 106724 108772
rect 106740 108828 106804 108832
rect 106740 108772 106744 108828
rect 106744 108772 106800 108828
rect 106800 108772 106804 108828
rect 106740 108768 106804 108772
rect 106820 108828 106884 108832
rect 106820 108772 106824 108828
rect 106824 108772 106880 108828
rect 106880 108772 106884 108828
rect 106820 108768 106884 108772
rect 106900 108828 106964 108832
rect 106900 108772 106904 108828
rect 106904 108772 106960 108828
rect 106960 108772 106964 108828
rect 106900 108768 106964 108772
rect 4216 108284 4280 108288
rect 4216 108228 4220 108284
rect 4220 108228 4276 108284
rect 4276 108228 4280 108284
rect 4216 108224 4280 108228
rect 4296 108284 4360 108288
rect 4296 108228 4300 108284
rect 4300 108228 4356 108284
rect 4356 108228 4360 108284
rect 4296 108224 4360 108228
rect 4376 108284 4440 108288
rect 4376 108228 4380 108284
rect 4380 108228 4436 108284
rect 4436 108228 4440 108284
rect 4376 108224 4440 108228
rect 4456 108284 4520 108288
rect 4456 108228 4460 108284
rect 4460 108228 4516 108284
rect 4516 108228 4520 108284
rect 4456 108224 4520 108228
rect 105924 108284 105988 108288
rect 105924 108228 105928 108284
rect 105928 108228 105984 108284
rect 105984 108228 105988 108284
rect 105924 108224 105988 108228
rect 106004 108284 106068 108288
rect 106004 108228 106008 108284
rect 106008 108228 106064 108284
rect 106064 108228 106068 108284
rect 106004 108224 106068 108228
rect 106084 108284 106148 108288
rect 106084 108228 106088 108284
rect 106088 108228 106144 108284
rect 106144 108228 106148 108284
rect 106084 108224 106148 108228
rect 106164 108284 106228 108288
rect 106164 108228 106168 108284
rect 106168 108228 106224 108284
rect 106224 108228 106228 108284
rect 106164 108224 106228 108228
rect 4876 107740 4940 107744
rect 4876 107684 4880 107740
rect 4880 107684 4936 107740
rect 4936 107684 4940 107740
rect 4876 107680 4940 107684
rect 4956 107740 5020 107744
rect 4956 107684 4960 107740
rect 4960 107684 5016 107740
rect 5016 107684 5020 107740
rect 4956 107680 5020 107684
rect 5036 107740 5100 107744
rect 5036 107684 5040 107740
rect 5040 107684 5096 107740
rect 5096 107684 5100 107740
rect 5036 107680 5100 107684
rect 5116 107740 5180 107744
rect 5116 107684 5120 107740
rect 5120 107684 5176 107740
rect 5176 107684 5180 107740
rect 5116 107680 5180 107684
rect 106660 107740 106724 107744
rect 106660 107684 106664 107740
rect 106664 107684 106720 107740
rect 106720 107684 106724 107740
rect 106660 107680 106724 107684
rect 106740 107740 106804 107744
rect 106740 107684 106744 107740
rect 106744 107684 106800 107740
rect 106800 107684 106804 107740
rect 106740 107680 106804 107684
rect 106820 107740 106884 107744
rect 106820 107684 106824 107740
rect 106824 107684 106880 107740
rect 106880 107684 106884 107740
rect 106820 107680 106884 107684
rect 106900 107740 106964 107744
rect 106900 107684 106904 107740
rect 106904 107684 106960 107740
rect 106960 107684 106964 107740
rect 106900 107680 106964 107684
rect 4216 107196 4280 107200
rect 4216 107140 4220 107196
rect 4220 107140 4276 107196
rect 4276 107140 4280 107196
rect 4216 107136 4280 107140
rect 4296 107196 4360 107200
rect 4296 107140 4300 107196
rect 4300 107140 4356 107196
rect 4356 107140 4360 107196
rect 4296 107136 4360 107140
rect 4376 107196 4440 107200
rect 4376 107140 4380 107196
rect 4380 107140 4436 107196
rect 4436 107140 4440 107196
rect 4376 107136 4440 107140
rect 4456 107196 4520 107200
rect 4456 107140 4460 107196
rect 4460 107140 4516 107196
rect 4516 107140 4520 107196
rect 4456 107136 4520 107140
rect 105924 107196 105988 107200
rect 105924 107140 105928 107196
rect 105928 107140 105984 107196
rect 105984 107140 105988 107196
rect 105924 107136 105988 107140
rect 106004 107196 106068 107200
rect 106004 107140 106008 107196
rect 106008 107140 106064 107196
rect 106064 107140 106068 107196
rect 106004 107136 106068 107140
rect 106084 107196 106148 107200
rect 106084 107140 106088 107196
rect 106088 107140 106144 107196
rect 106144 107140 106148 107196
rect 106084 107136 106148 107140
rect 106164 107196 106228 107200
rect 106164 107140 106168 107196
rect 106168 107140 106224 107196
rect 106224 107140 106228 107196
rect 106164 107136 106228 107140
rect 4876 106652 4940 106656
rect 4876 106596 4880 106652
rect 4880 106596 4936 106652
rect 4936 106596 4940 106652
rect 4876 106592 4940 106596
rect 4956 106652 5020 106656
rect 4956 106596 4960 106652
rect 4960 106596 5016 106652
rect 5016 106596 5020 106652
rect 4956 106592 5020 106596
rect 5036 106652 5100 106656
rect 5036 106596 5040 106652
rect 5040 106596 5096 106652
rect 5096 106596 5100 106652
rect 5036 106592 5100 106596
rect 5116 106652 5180 106656
rect 5116 106596 5120 106652
rect 5120 106596 5176 106652
rect 5176 106596 5180 106652
rect 5116 106592 5180 106596
rect 106660 106652 106724 106656
rect 106660 106596 106664 106652
rect 106664 106596 106720 106652
rect 106720 106596 106724 106652
rect 106660 106592 106724 106596
rect 106740 106652 106804 106656
rect 106740 106596 106744 106652
rect 106744 106596 106800 106652
rect 106800 106596 106804 106652
rect 106740 106592 106804 106596
rect 106820 106652 106884 106656
rect 106820 106596 106824 106652
rect 106824 106596 106880 106652
rect 106880 106596 106884 106652
rect 106820 106592 106884 106596
rect 106900 106652 106964 106656
rect 106900 106596 106904 106652
rect 106904 106596 106960 106652
rect 106960 106596 106964 106652
rect 106900 106592 106964 106596
rect 4216 106108 4280 106112
rect 4216 106052 4220 106108
rect 4220 106052 4276 106108
rect 4276 106052 4280 106108
rect 4216 106048 4280 106052
rect 4296 106108 4360 106112
rect 4296 106052 4300 106108
rect 4300 106052 4356 106108
rect 4356 106052 4360 106108
rect 4296 106048 4360 106052
rect 4376 106108 4440 106112
rect 4376 106052 4380 106108
rect 4380 106052 4436 106108
rect 4436 106052 4440 106108
rect 4376 106048 4440 106052
rect 4456 106108 4520 106112
rect 4456 106052 4460 106108
rect 4460 106052 4516 106108
rect 4516 106052 4520 106108
rect 4456 106048 4520 106052
rect 105924 106108 105988 106112
rect 105924 106052 105928 106108
rect 105928 106052 105984 106108
rect 105984 106052 105988 106108
rect 105924 106048 105988 106052
rect 106004 106108 106068 106112
rect 106004 106052 106008 106108
rect 106008 106052 106064 106108
rect 106064 106052 106068 106108
rect 106004 106048 106068 106052
rect 106084 106108 106148 106112
rect 106084 106052 106088 106108
rect 106088 106052 106144 106108
rect 106144 106052 106148 106108
rect 106084 106048 106148 106052
rect 106164 106108 106228 106112
rect 106164 106052 106168 106108
rect 106168 106052 106224 106108
rect 106224 106052 106228 106108
rect 106164 106048 106228 106052
rect 4876 105564 4940 105568
rect 4876 105508 4880 105564
rect 4880 105508 4936 105564
rect 4936 105508 4940 105564
rect 4876 105504 4940 105508
rect 4956 105564 5020 105568
rect 4956 105508 4960 105564
rect 4960 105508 5016 105564
rect 5016 105508 5020 105564
rect 4956 105504 5020 105508
rect 5036 105564 5100 105568
rect 5036 105508 5040 105564
rect 5040 105508 5096 105564
rect 5096 105508 5100 105564
rect 5036 105504 5100 105508
rect 5116 105564 5180 105568
rect 5116 105508 5120 105564
rect 5120 105508 5176 105564
rect 5176 105508 5180 105564
rect 5116 105504 5180 105508
rect 106660 105564 106724 105568
rect 106660 105508 106664 105564
rect 106664 105508 106720 105564
rect 106720 105508 106724 105564
rect 106660 105504 106724 105508
rect 106740 105564 106804 105568
rect 106740 105508 106744 105564
rect 106744 105508 106800 105564
rect 106800 105508 106804 105564
rect 106740 105504 106804 105508
rect 106820 105564 106884 105568
rect 106820 105508 106824 105564
rect 106824 105508 106880 105564
rect 106880 105508 106884 105564
rect 106820 105504 106884 105508
rect 106900 105564 106964 105568
rect 106900 105508 106904 105564
rect 106904 105508 106960 105564
rect 106960 105508 106964 105564
rect 106900 105504 106964 105508
rect 4216 105020 4280 105024
rect 4216 104964 4220 105020
rect 4220 104964 4276 105020
rect 4276 104964 4280 105020
rect 4216 104960 4280 104964
rect 4296 105020 4360 105024
rect 4296 104964 4300 105020
rect 4300 104964 4356 105020
rect 4356 104964 4360 105020
rect 4296 104960 4360 104964
rect 4376 105020 4440 105024
rect 4376 104964 4380 105020
rect 4380 104964 4436 105020
rect 4436 104964 4440 105020
rect 4376 104960 4440 104964
rect 4456 105020 4520 105024
rect 4456 104964 4460 105020
rect 4460 104964 4516 105020
rect 4516 104964 4520 105020
rect 4456 104960 4520 104964
rect 105924 105020 105988 105024
rect 105924 104964 105928 105020
rect 105928 104964 105984 105020
rect 105984 104964 105988 105020
rect 105924 104960 105988 104964
rect 106004 105020 106068 105024
rect 106004 104964 106008 105020
rect 106008 104964 106064 105020
rect 106064 104964 106068 105020
rect 106004 104960 106068 104964
rect 106084 105020 106148 105024
rect 106084 104964 106088 105020
rect 106088 104964 106144 105020
rect 106144 104964 106148 105020
rect 106084 104960 106148 104964
rect 106164 105020 106228 105024
rect 106164 104964 106168 105020
rect 106168 104964 106224 105020
rect 106224 104964 106228 105020
rect 106164 104960 106228 104964
rect 4876 104476 4940 104480
rect 4876 104420 4880 104476
rect 4880 104420 4936 104476
rect 4936 104420 4940 104476
rect 4876 104416 4940 104420
rect 4956 104476 5020 104480
rect 4956 104420 4960 104476
rect 4960 104420 5016 104476
rect 5016 104420 5020 104476
rect 4956 104416 5020 104420
rect 5036 104476 5100 104480
rect 5036 104420 5040 104476
rect 5040 104420 5096 104476
rect 5096 104420 5100 104476
rect 5036 104416 5100 104420
rect 5116 104476 5180 104480
rect 5116 104420 5120 104476
rect 5120 104420 5176 104476
rect 5176 104420 5180 104476
rect 5116 104416 5180 104420
rect 106660 104476 106724 104480
rect 106660 104420 106664 104476
rect 106664 104420 106720 104476
rect 106720 104420 106724 104476
rect 106660 104416 106724 104420
rect 106740 104476 106804 104480
rect 106740 104420 106744 104476
rect 106744 104420 106800 104476
rect 106800 104420 106804 104476
rect 106740 104416 106804 104420
rect 106820 104476 106884 104480
rect 106820 104420 106824 104476
rect 106824 104420 106880 104476
rect 106880 104420 106884 104476
rect 106820 104416 106884 104420
rect 106900 104476 106964 104480
rect 106900 104420 106904 104476
rect 106904 104420 106960 104476
rect 106960 104420 106964 104476
rect 106900 104416 106964 104420
rect 4216 103932 4280 103936
rect 4216 103876 4220 103932
rect 4220 103876 4276 103932
rect 4276 103876 4280 103932
rect 4216 103872 4280 103876
rect 4296 103932 4360 103936
rect 4296 103876 4300 103932
rect 4300 103876 4356 103932
rect 4356 103876 4360 103932
rect 4296 103872 4360 103876
rect 4376 103932 4440 103936
rect 4376 103876 4380 103932
rect 4380 103876 4436 103932
rect 4436 103876 4440 103932
rect 4376 103872 4440 103876
rect 4456 103932 4520 103936
rect 4456 103876 4460 103932
rect 4460 103876 4516 103932
rect 4516 103876 4520 103932
rect 4456 103872 4520 103876
rect 105924 103932 105988 103936
rect 105924 103876 105928 103932
rect 105928 103876 105984 103932
rect 105984 103876 105988 103932
rect 105924 103872 105988 103876
rect 106004 103932 106068 103936
rect 106004 103876 106008 103932
rect 106008 103876 106064 103932
rect 106064 103876 106068 103932
rect 106004 103872 106068 103876
rect 106084 103932 106148 103936
rect 106084 103876 106088 103932
rect 106088 103876 106144 103932
rect 106144 103876 106148 103932
rect 106084 103872 106148 103876
rect 106164 103932 106228 103936
rect 106164 103876 106168 103932
rect 106168 103876 106224 103932
rect 106224 103876 106228 103932
rect 106164 103872 106228 103876
rect 4876 103388 4940 103392
rect 4876 103332 4880 103388
rect 4880 103332 4936 103388
rect 4936 103332 4940 103388
rect 4876 103328 4940 103332
rect 4956 103388 5020 103392
rect 4956 103332 4960 103388
rect 4960 103332 5016 103388
rect 5016 103332 5020 103388
rect 4956 103328 5020 103332
rect 5036 103388 5100 103392
rect 5036 103332 5040 103388
rect 5040 103332 5096 103388
rect 5096 103332 5100 103388
rect 5036 103328 5100 103332
rect 5116 103388 5180 103392
rect 5116 103332 5120 103388
rect 5120 103332 5176 103388
rect 5176 103332 5180 103388
rect 5116 103328 5180 103332
rect 106660 103388 106724 103392
rect 106660 103332 106664 103388
rect 106664 103332 106720 103388
rect 106720 103332 106724 103388
rect 106660 103328 106724 103332
rect 106740 103388 106804 103392
rect 106740 103332 106744 103388
rect 106744 103332 106800 103388
rect 106800 103332 106804 103388
rect 106740 103328 106804 103332
rect 106820 103388 106884 103392
rect 106820 103332 106824 103388
rect 106824 103332 106880 103388
rect 106880 103332 106884 103388
rect 106820 103328 106884 103332
rect 106900 103388 106964 103392
rect 106900 103332 106904 103388
rect 106904 103332 106960 103388
rect 106960 103332 106964 103388
rect 106900 103328 106964 103332
rect 4216 102844 4280 102848
rect 4216 102788 4220 102844
rect 4220 102788 4276 102844
rect 4276 102788 4280 102844
rect 4216 102784 4280 102788
rect 4296 102844 4360 102848
rect 4296 102788 4300 102844
rect 4300 102788 4356 102844
rect 4356 102788 4360 102844
rect 4296 102784 4360 102788
rect 4376 102844 4440 102848
rect 4376 102788 4380 102844
rect 4380 102788 4436 102844
rect 4436 102788 4440 102844
rect 4376 102784 4440 102788
rect 4456 102844 4520 102848
rect 4456 102788 4460 102844
rect 4460 102788 4516 102844
rect 4516 102788 4520 102844
rect 4456 102784 4520 102788
rect 105924 102844 105988 102848
rect 105924 102788 105928 102844
rect 105928 102788 105984 102844
rect 105984 102788 105988 102844
rect 105924 102784 105988 102788
rect 106004 102844 106068 102848
rect 106004 102788 106008 102844
rect 106008 102788 106064 102844
rect 106064 102788 106068 102844
rect 106004 102784 106068 102788
rect 106084 102844 106148 102848
rect 106084 102788 106088 102844
rect 106088 102788 106144 102844
rect 106144 102788 106148 102844
rect 106084 102784 106148 102788
rect 106164 102844 106228 102848
rect 106164 102788 106168 102844
rect 106168 102788 106224 102844
rect 106224 102788 106228 102844
rect 106164 102784 106228 102788
rect 4876 102300 4940 102304
rect 4876 102244 4880 102300
rect 4880 102244 4936 102300
rect 4936 102244 4940 102300
rect 4876 102240 4940 102244
rect 4956 102300 5020 102304
rect 4956 102244 4960 102300
rect 4960 102244 5016 102300
rect 5016 102244 5020 102300
rect 4956 102240 5020 102244
rect 5036 102300 5100 102304
rect 5036 102244 5040 102300
rect 5040 102244 5096 102300
rect 5096 102244 5100 102300
rect 5036 102240 5100 102244
rect 5116 102300 5180 102304
rect 5116 102244 5120 102300
rect 5120 102244 5176 102300
rect 5176 102244 5180 102300
rect 5116 102240 5180 102244
rect 106660 102300 106724 102304
rect 106660 102244 106664 102300
rect 106664 102244 106720 102300
rect 106720 102244 106724 102300
rect 106660 102240 106724 102244
rect 106740 102300 106804 102304
rect 106740 102244 106744 102300
rect 106744 102244 106800 102300
rect 106800 102244 106804 102300
rect 106740 102240 106804 102244
rect 106820 102300 106884 102304
rect 106820 102244 106824 102300
rect 106824 102244 106880 102300
rect 106880 102244 106884 102300
rect 106820 102240 106884 102244
rect 106900 102300 106964 102304
rect 106900 102244 106904 102300
rect 106904 102244 106960 102300
rect 106960 102244 106964 102300
rect 106900 102240 106964 102244
rect 4216 101756 4280 101760
rect 4216 101700 4220 101756
rect 4220 101700 4276 101756
rect 4276 101700 4280 101756
rect 4216 101696 4280 101700
rect 4296 101756 4360 101760
rect 4296 101700 4300 101756
rect 4300 101700 4356 101756
rect 4356 101700 4360 101756
rect 4296 101696 4360 101700
rect 4376 101756 4440 101760
rect 4376 101700 4380 101756
rect 4380 101700 4436 101756
rect 4436 101700 4440 101756
rect 4376 101696 4440 101700
rect 4456 101756 4520 101760
rect 4456 101700 4460 101756
rect 4460 101700 4516 101756
rect 4516 101700 4520 101756
rect 4456 101696 4520 101700
rect 105924 101756 105988 101760
rect 105924 101700 105928 101756
rect 105928 101700 105984 101756
rect 105984 101700 105988 101756
rect 105924 101696 105988 101700
rect 106004 101756 106068 101760
rect 106004 101700 106008 101756
rect 106008 101700 106064 101756
rect 106064 101700 106068 101756
rect 106004 101696 106068 101700
rect 106084 101756 106148 101760
rect 106084 101700 106088 101756
rect 106088 101700 106144 101756
rect 106144 101700 106148 101756
rect 106084 101696 106148 101700
rect 106164 101756 106228 101760
rect 106164 101700 106168 101756
rect 106168 101700 106224 101756
rect 106224 101700 106228 101756
rect 106164 101696 106228 101700
rect 4876 101212 4940 101216
rect 4876 101156 4880 101212
rect 4880 101156 4936 101212
rect 4936 101156 4940 101212
rect 4876 101152 4940 101156
rect 4956 101212 5020 101216
rect 4956 101156 4960 101212
rect 4960 101156 5016 101212
rect 5016 101156 5020 101212
rect 4956 101152 5020 101156
rect 5036 101212 5100 101216
rect 5036 101156 5040 101212
rect 5040 101156 5096 101212
rect 5096 101156 5100 101212
rect 5036 101152 5100 101156
rect 5116 101212 5180 101216
rect 5116 101156 5120 101212
rect 5120 101156 5176 101212
rect 5176 101156 5180 101212
rect 5116 101152 5180 101156
rect 106660 101212 106724 101216
rect 106660 101156 106664 101212
rect 106664 101156 106720 101212
rect 106720 101156 106724 101212
rect 106660 101152 106724 101156
rect 106740 101212 106804 101216
rect 106740 101156 106744 101212
rect 106744 101156 106800 101212
rect 106800 101156 106804 101212
rect 106740 101152 106804 101156
rect 106820 101212 106884 101216
rect 106820 101156 106824 101212
rect 106824 101156 106880 101212
rect 106880 101156 106884 101212
rect 106820 101152 106884 101156
rect 106900 101212 106964 101216
rect 106900 101156 106904 101212
rect 106904 101156 106960 101212
rect 106960 101156 106964 101212
rect 106900 101152 106964 101156
rect 4216 100668 4280 100672
rect 4216 100612 4220 100668
rect 4220 100612 4276 100668
rect 4276 100612 4280 100668
rect 4216 100608 4280 100612
rect 4296 100668 4360 100672
rect 4296 100612 4300 100668
rect 4300 100612 4356 100668
rect 4356 100612 4360 100668
rect 4296 100608 4360 100612
rect 4376 100668 4440 100672
rect 4376 100612 4380 100668
rect 4380 100612 4436 100668
rect 4436 100612 4440 100668
rect 4376 100608 4440 100612
rect 4456 100668 4520 100672
rect 4456 100612 4460 100668
rect 4460 100612 4516 100668
rect 4516 100612 4520 100668
rect 4456 100608 4520 100612
rect 105924 100668 105988 100672
rect 105924 100612 105928 100668
rect 105928 100612 105984 100668
rect 105984 100612 105988 100668
rect 105924 100608 105988 100612
rect 106004 100668 106068 100672
rect 106004 100612 106008 100668
rect 106008 100612 106064 100668
rect 106064 100612 106068 100668
rect 106004 100608 106068 100612
rect 106084 100668 106148 100672
rect 106084 100612 106088 100668
rect 106088 100612 106144 100668
rect 106144 100612 106148 100668
rect 106084 100608 106148 100612
rect 106164 100668 106228 100672
rect 106164 100612 106168 100668
rect 106168 100612 106224 100668
rect 106224 100612 106228 100668
rect 106164 100608 106228 100612
rect 4876 100124 4940 100128
rect 4876 100068 4880 100124
rect 4880 100068 4936 100124
rect 4936 100068 4940 100124
rect 4876 100064 4940 100068
rect 4956 100124 5020 100128
rect 4956 100068 4960 100124
rect 4960 100068 5016 100124
rect 5016 100068 5020 100124
rect 4956 100064 5020 100068
rect 5036 100124 5100 100128
rect 5036 100068 5040 100124
rect 5040 100068 5096 100124
rect 5096 100068 5100 100124
rect 5036 100064 5100 100068
rect 5116 100124 5180 100128
rect 5116 100068 5120 100124
rect 5120 100068 5176 100124
rect 5176 100068 5180 100124
rect 5116 100064 5180 100068
rect 106660 100124 106724 100128
rect 106660 100068 106664 100124
rect 106664 100068 106720 100124
rect 106720 100068 106724 100124
rect 106660 100064 106724 100068
rect 106740 100124 106804 100128
rect 106740 100068 106744 100124
rect 106744 100068 106800 100124
rect 106800 100068 106804 100124
rect 106740 100064 106804 100068
rect 106820 100124 106884 100128
rect 106820 100068 106824 100124
rect 106824 100068 106880 100124
rect 106880 100068 106884 100124
rect 106820 100064 106884 100068
rect 106900 100124 106964 100128
rect 106900 100068 106904 100124
rect 106904 100068 106960 100124
rect 106960 100068 106964 100124
rect 106900 100064 106964 100068
rect 4216 99580 4280 99584
rect 4216 99524 4220 99580
rect 4220 99524 4276 99580
rect 4276 99524 4280 99580
rect 4216 99520 4280 99524
rect 4296 99580 4360 99584
rect 4296 99524 4300 99580
rect 4300 99524 4356 99580
rect 4356 99524 4360 99580
rect 4296 99520 4360 99524
rect 4376 99580 4440 99584
rect 4376 99524 4380 99580
rect 4380 99524 4436 99580
rect 4436 99524 4440 99580
rect 4376 99520 4440 99524
rect 4456 99580 4520 99584
rect 4456 99524 4460 99580
rect 4460 99524 4516 99580
rect 4516 99524 4520 99580
rect 4456 99520 4520 99524
rect 105924 99580 105988 99584
rect 105924 99524 105928 99580
rect 105928 99524 105984 99580
rect 105984 99524 105988 99580
rect 105924 99520 105988 99524
rect 106004 99580 106068 99584
rect 106004 99524 106008 99580
rect 106008 99524 106064 99580
rect 106064 99524 106068 99580
rect 106004 99520 106068 99524
rect 106084 99580 106148 99584
rect 106084 99524 106088 99580
rect 106088 99524 106144 99580
rect 106144 99524 106148 99580
rect 106084 99520 106148 99524
rect 106164 99580 106228 99584
rect 106164 99524 106168 99580
rect 106168 99524 106224 99580
rect 106224 99524 106228 99580
rect 106164 99520 106228 99524
rect 4876 99036 4940 99040
rect 4876 98980 4880 99036
rect 4880 98980 4936 99036
rect 4936 98980 4940 99036
rect 4876 98976 4940 98980
rect 4956 99036 5020 99040
rect 4956 98980 4960 99036
rect 4960 98980 5016 99036
rect 5016 98980 5020 99036
rect 4956 98976 5020 98980
rect 5036 99036 5100 99040
rect 5036 98980 5040 99036
rect 5040 98980 5096 99036
rect 5096 98980 5100 99036
rect 5036 98976 5100 98980
rect 5116 99036 5180 99040
rect 5116 98980 5120 99036
rect 5120 98980 5176 99036
rect 5176 98980 5180 99036
rect 5116 98976 5180 98980
rect 106660 99036 106724 99040
rect 106660 98980 106664 99036
rect 106664 98980 106720 99036
rect 106720 98980 106724 99036
rect 106660 98976 106724 98980
rect 106740 99036 106804 99040
rect 106740 98980 106744 99036
rect 106744 98980 106800 99036
rect 106800 98980 106804 99036
rect 106740 98976 106804 98980
rect 106820 99036 106884 99040
rect 106820 98980 106824 99036
rect 106824 98980 106880 99036
rect 106880 98980 106884 99036
rect 106820 98976 106884 98980
rect 106900 99036 106964 99040
rect 106900 98980 106904 99036
rect 106904 98980 106960 99036
rect 106960 98980 106964 99036
rect 106900 98976 106964 98980
rect 4216 98492 4280 98496
rect 4216 98436 4220 98492
rect 4220 98436 4276 98492
rect 4276 98436 4280 98492
rect 4216 98432 4280 98436
rect 4296 98492 4360 98496
rect 4296 98436 4300 98492
rect 4300 98436 4356 98492
rect 4356 98436 4360 98492
rect 4296 98432 4360 98436
rect 4376 98492 4440 98496
rect 4376 98436 4380 98492
rect 4380 98436 4436 98492
rect 4436 98436 4440 98492
rect 4376 98432 4440 98436
rect 4456 98492 4520 98496
rect 4456 98436 4460 98492
rect 4460 98436 4516 98492
rect 4516 98436 4520 98492
rect 4456 98432 4520 98436
rect 105924 98492 105988 98496
rect 105924 98436 105928 98492
rect 105928 98436 105984 98492
rect 105984 98436 105988 98492
rect 105924 98432 105988 98436
rect 106004 98492 106068 98496
rect 106004 98436 106008 98492
rect 106008 98436 106064 98492
rect 106064 98436 106068 98492
rect 106004 98432 106068 98436
rect 106084 98492 106148 98496
rect 106084 98436 106088 98492
rect 106088 98436 106144 98492
rect 106144 98436 106148 98492
rect 106084 98432 106148 98436
rect 106164 98492 106228 98496
rect 106164 98436 106168 98492
rect 106168 98436 106224 98492
rect 106224 98436 106228 98492
rect 106164 98432 106228 98436
rect 4876 97948 4940 97952
rect 4876 97892 4880 97948
rect 4880 97892 4936 97948
rect 4936 97892 4940 97948
rect 4876 97888 4940 97892
rect 4956 97948 5020 97952
rect 4956 97892 4960 97948
rect 4960 97892 5016 97948
rect 5016 97892 5020 97948
rect 4956 97888 5020 97892
rect 5036 97948 5100 97952
rect 5036 97892 5040 97948
rect 5040 97892 5096 97948
rect 5096 97892 5100 97948
rect 5036 97888 5100 97892
rect 5116 97948 5180 97952
rect 5116 97892 5120 97948
rect 5120 97892 5176 97948
rect 5176 97892 5180 97948
rect 5116 97888 5180 97892
rect 106660 97948 106724 97952
rect 106660 97892 106664 97948
rect 106664 97892 106720 97948
rect 106720 97892 106724 97948
rect 106660 97888 106724 97892
rect 106740 97948 106804 97952
rect 106740 97892 106744 97948
rect 106744 97892 106800 97948
rect 106800 97892 106804 97948
rect 106740 97888 106804 97892
rect 106820 97948 106884 97952
rect 106820 97892 106824 97948
rect 106824 97892 106880 97948
rect 106880 97892 106884 97948
rect 106820 97888 106884 97892
rect 106900 97948 106964 97952
rect 106900 97892 106904 97948
rect 106904 97892 106960 97948
rect 106960 97892 106964 97948
rect 106900 97888 106964 97892
rect 4216 97404 4280 97408
rect 4216 97348 4220 97404
rect 4220 97348 4276 97404
rect 4276 97348 4280 97404
rect 4216 97344 4280 97348
rect 4296 97404 4360 97408
rect 4296 97348 4300 97404
rect 4300 97348 4356 97404
rect 4356 97348 4360 97404
rect 4296 97344 4360 97348
rect 4376 97404 4440 97408
rect 4376 97348 4380 97404
rect 4380 97348 4436 97404
rect 4436 97348 4440 97404
rect 4376 97344 4440 97348
rect 4456 97404 4520 97408
rect 4456 97348 4460 97404
rect 4460 97348 4516 97404
rect 4516 97348 4520 97404
rect 4456 97344 4520 97348
rect 105924 97404 105988 97408
rect 105924 97348 105928 97404
rect 105928 97348 105984 97404
rect 105984 97348 105988 97404
rect 105924 97344 105988 97348
rect 106004 97404 106068 97408
rect 106004 97348 106008 97404
rect 106008 97348 106064 97404
rect 106064 97348 106068 97404
rect 106004 97344 106068 97348
rect 106084 97404 106148 97408
rect 106084 97348 106088 97404
rect 106088 97348 106144 97404
rect 106144 97348 106148 97404
rect 106084 97344 106148 97348
rect 106164 97404 106228 97408
rect 106164 97348 106168 97404
rect 106168 97348 106224 97404
rect 106224 97348 106228 97404
rect 106164 97344 106228 97348
rect 4876 96860 4940 96864
rect 4876 96804 4880 96860
rect 4880 96804 4936 96860
rect 4936 96804 4940 96860
rect 4876 96800 4940 96804
rect 4956 96860 5020 96864
rect 4956 96804 4960 96860
rect 4960 96804 5016 96860
rect 5016 96804 5020 96860
rect 4956 96800 5020 96804
rect 5036 96860 5100 96864
rect 5036 96804 5040 96860
rect 5040 96804 5096 96860
rect 5096 96804 5100 96860
rect 5036 96800 5100 96804
rect 5116 96860 5180 96864
rect 5116 96804 5120 96860
rect 5120 96804 5176 96860
rect 5176 96804 5180 96860
rect 5116 96800 5180 96804
rect 106660 96860 106724 96864
rect 106660 96804 106664 96860
rect 106664 96804 106720 96860
rect 106720 96804 106724 96860
rect 106660 96800 106724 96804
rect 106740 96860 106804 96864
rect 106740 96804 106744 96860
rect 106744 96804 106800 96860
rect 106800 96804 106804 96860
rect 106740 96800 106804 96804
rect 106820 96860 106884 96864
rect 106820 96804 106824 96860
rect 106824 96804 106880 96860
rect 106880 96804 106884 96860
rect 106820 96800 106884 96804
rect 106900 96860 106964 96864
rect 106900 96804 106904 96860
rect 106904 96804 106960 96860
rect 106960 96804 106964 96860
rect 106900 96800 106964 96804
rect 4216 96316 4280 96320
rect 4216 96260 4220 96316
rect 4220 96260 4276 96316
rect 4276 96260 4280 96316
rect 4216 96256 4280 96260
rect 4296 96316 4360 96320
rect 4296 96260 4300 96316
rect 4300 96260 4356 96316
rect 4356 96260 4360 96316
rect 4296 96256 4360 96260
rect 4376 96316 4440 96320
rect 4376 96260 4380 96316
rect 4380 96260 4436 96316
rect 4436 96260 4440 96316
rect 4376 96256 4440 96260
rect 4456 96316 4520 96320
rect 4456 96260 4460 96316
rect 4460 96260 4516 96316
rect 4516 96260 4520 96316
rect 4456 96256 4520 96260
rect 105924 96316 105988 96320
rect 105924 96260 105928 96316
rect 105928 96260 105984 96316
rect 105984 96260 105988 96316
rect 105924 96256 105988 96260
rect 106004 96316 106068 96320
rect 106004 96260 106008 96316
rect 106008 96260 106064 96316
rect 106064 96260 106068 96316
rect 106004 96256 106068 96260
rect 106084 96316 106148 96320
rect 106084 96260 106088 96316
rect 106088 96260 106144 96316
rect 106144 96260 106148 96316
rect 106084 96256 106148 96260
rect 106164 96316 106228 96320
rect 106164 96260 106168 96316
rect 106168 96260 106224 96316
rect 106224 96260 106228 96316
rect 106164 96256 106228 96260
rect 4876 95772 4940 95776
rect 4876 95716 4880 95772
rect 4880 95716 4936 95772
rect 4936 95716 4940 95772
rect 4876 95712 4940 95716
rect 4956 95772 5020 95776
rect 4956 95716 4960 95772
rect 4960 95716 5016 95772
rect 5016 95716 5020 95772
rect 4956 95712 5020 95716
rect 5036 95772 5100 95776
rect 5036 95716 5040 95772
rect 5040 95716 5096 95772
rect 5096 95716 5100 95772
rect 5036 95712 5100 95716
rect 5116 95772 5180 95776
rect 5116 95716 5120 95772
rect 5120 95716 5176 95772
rect 5176 95716 5180 95772
rect 5116 95712 5180 95716
rect 106660 95772 106724 95776
rect 106660 95716 106664 95772
rect 106664 95716 106720 95772
rect 106720 95716 106724 95772
rect 106660 95712 106724 95716
rect 106740 95772 106804 95776
rect 106740 95716 106744 95772
rect 106744 95716 106800 95772
rect 106800 95716 106804 95772
rect 106740 95712 106804 95716
rect 106820 95772 106884 95776
rect 106820 95716 106824 95772
rect 106824 95716 106880 95772
rect 106880 95716 106884 95772
rect 106820 95712 106884 95716
rect 106900 95772 106964 95776
rect 106900 95716 106904 95772
rect 106904 95716 106960 95772
rect 106960 95716 106964 95772
rect 106900 95712 106964 95716
rect 4216 95228 4280 95232
rect 4216 95172 4220 95228
rect 4220 95172 4276 95228
rect 4276 95172 4280 95228
rect 4216 95168 4280 95172
rect 4296 95228 4360 95232
rect 4296 95172 4300 95228
rect 4300 95172 4356 95228
rect 4356 95172 4360 95228
rect 4296 95168 4360 95172
rect 4376 95228 4440 95232
rect 4376 95172 4380 95228
rect 4380 95172 4436 95228
rect 4436 95172 4440 95228
rect 4376 95168 4440 95172
rect 4456 95228 4520 95232
rect 4456 95172 4460 95228
rect 4460 95172 4516 95228
rect 4516 95172 4520 95228
rect 4456 95168 4520 95172
rect 105924 95228 105988 95232
rect 105924 95172 105928 95228
rect 105928 95172 105984 95228
rect 105984 95172 105988 95228
rect 105924 95168 105988 95172
rect 106004 95228 106068 95232
rect 106004 95172 106008 95228
rect 106008 95172 106064 95228
rect 106064 95172 106068 95228
rect 106004 95168 106068 95172
rect 106084 95228 106148 95232
rect 106084 95172 106088 95228
rect 106088 95172 106144 95228
rect 106144 95172 106148 95228
rect 106084 95168 106148 95172
rect 106164 95228 106228 95232
rect 106164 95172 106168 95228
rect 106168 95172 106224 95228
rect 106224 95172 106228 95228
rect 106164 95168 106228 95172
rect 4876 94684 4940 94688
rect 4876 94628 4880 94684
rect 4880 94628 4936 94684
rect 4936 94628 4940 94684
rect 4876 94624 4940 94628
rect 4956 94684 5020 94688
rect 4956 94628 4960 94684
rect 4960 94628 5016 94684
rect 5016 94628 5020 94684
rect 4956 94624 5020 94628
rect 5036 94684 5100 94688
rect 5036 94628 5040 94684
rect 5040 94628 5096 94684
rect 5096 94628 5100 94684
rect 5036 94624 5100 94628
rect 5116 94684 5180 94688
rect 5116 94628 5120 94684
rect 5120 94628 5176 94684
rect 5176 94628 5180 94684
rect 5116 94624 5180 94628
rect 106660 94684 106724 94688
rect 106660 94628 106664 94684
rect 106664 94628 106720 94684
rect 106720 94628 106724 94684
rect 106660 94624 106724 94628
rect 106740 94684 106804 94688
rect 106740 94628 106744 94684
rect 106744 94628 106800 94684
rect 106800 94628 106804 94684
rect 106740 94624 106804 94628
rect 106820 94684 106884 94688
rect 106820 94628 106824 94684
rect 106824 94628 106880 94684
rect 106880 94628 106884 94684
rect 106820 94624 106884 94628
rect 106900 94684 106964 94688
rect 106900 94628 106904 94684
rect 106904 94628 106960 94684
rect 106960 94628 106964 94684
rect 106900 94624 106964 94628
rect 4216 94140 4280 94144
rect 4216 94084 4220 94140
rect 4220 94084 4276 94140
rect 4276 94084 4280 94140
rect 4216 94080 4280 94084
rect 4296 94140 4360 94144
rect 4296 94084 4300 94140
rect 4300 94084 4356 94140
rect 4356 94084 4360 94140
rect 4296 94080 4360 94084
rect 4376 94140 4440 94144
rect 4376 94084 4380 94140
rect 4380 94084 4436 94140
rect 4436 94084 4440 94140
rect 4376 94080 4440 94084
rect 4456 94140 4520 94144
rect 4456 94084 4460 94140
rect 4460 94084 4516 94140
rect 4516 94084 4520 94140
rect 4456 94080 4520 94084
rect 105924 94140 105988 94144
rect 105924 94084 105928 94140
rect 105928 94084 105984 94140
rect 105984 94084 105988 94140
rect 105924 94080 105988 94084
rect 106004 94140 106068 94144
rect 106004 94084 106008 94140
rect 106008 94084 106064 94140
rect 106064 94084 106068 94140
rect 106004 94080 106068 94084
rect 106084 94140 106148 94144
rect 106084 94084 106088 94140
rect 106088 94084 106144 94140
rect 106144 94084 106148 94140
rect 106084 94080 106148 94084
rect 106164 94140 106228 94144
rect 106164 94084 106168 94140
rect 106168 94084 106224 94140
rect 106224 94084 106228 94140
rect 106164 94080 106228 94084
rect 4876 93596 4940 93600
rect 4876 93540 4880 93596
rect 4880 93540 4936 93596
rect 4936 93540 4940 93596
rect 4876 93536 4940 93540
rect 4956 93596 5020 93600
rect 4956 93540 4960 93596
rect 4960 93540 5016 93596
rect 5016 93540 5020 93596
rect 4956 93536 5020 93540
rect 5036 93596 5100 93600
rect 5036 93540 5040 93596
rect 5040 93540 5096 93596
rect 5096 93540 5100 93596
rect 5036 93536 5100 93540
rect 5116 93596 5180 93600
rect 5116 93540 5120 93596
rect 5120 93540 5176 93596
rect 5176 93540 5180 93596
rect 5116 93536 5180 93540
rect 106660 93596 106724 93600
rect 106660 93540 106664 93596
rect 106664 93540 106720 93596
rect 106720 93540 106724 93596
rect 106660 93536 106724 93540
rect 106740 93596 106804 93600
rect 106740 93540 106744 93596
rect 106744 93540 106800 93596
rect 106800 93540 106804 93596
rect 106740 93536 106804 93540
rect 106820 93596 106884 93600
rect 106820 93540 106824 93596
rect 106824 93540 106880 93596
rect 106880 93540 106884 93596
rect 106820 93536 106884 93540
rect 106900 93596 106964 93600
rect 106900 93540 106904 93596
rect 106904 93540 106960 93596
rect 106960 93540 106964 93596
rect 106900 93536 106964 93540
rect 4216 93052 4280 93056
rect 4216 92996 4220 93052
rect 4220 92996 4276 93052
rect 4276 92996 4280 93052
rect 4216 92992 4280 92996
rect 4296 93052 4360 93056
rect 4296 92996 4300 93052
rect 4300 92996 4356 93052
rect 4356 92996 4360 93052
rect 4296 92992 4360 92996
rect 4376 93052 4440 93056
rect 4376 92996 4380 93052
rect 4380 92996 4436 93052
rect 4436 92996 4440 93052
rect 4376 92992 4440 92996
rect 4456 93052 4520 93056
rect 4456 92996 4460 93052
rect 4460 92996 4516 93052
rect 4516 92996 4520 93052
rect 4456 92992 4520 92996
rect 105924 93052 105988 93056
rect 105924 92996 105928 93052
rect 105928 92996 105984 93052
rect 105984 92996 105988 93052
rect 105924 92992 105988 92996
rect 106004 93052 106068 93056
rect 106004 92996 106008 93052
rect 106008 92996 106064 93052
rect 106064 92996 106068 93052
rect 106004 92992 106068 92996
rect 106084 93052 106148 93056
rect 106084 92996 106088 93052
rect 106088 92996 106144 93052
rect 106144 92996 106148 93052
rect 106084 92992 106148 92996
rect 106164 93052 106228 93056
rect 106164 92996 106168 93052
rect 106168 92996 106224 93052
rect 106224 92996 106228 93052
rect 106164 92992 106228 92996
rect 4876 92508 4940 92512
rect 4876 92452 4880 92508
rect 4880 92452 4936 92508
rect 4936 92452 4940 92508
rect 4876 92448 4940 92452
rect 4956 92508 5020 92512
rect 4956 92452 4960 92508
rect 4960 92452 5016 92508
rect 5016 92452 5020 92508
rect 4956 92448 5020 92452
rect 5036 92508 5100 92512
rect 5036 92452 5040 92508
rect 5040 92452 5096 92508
rect 5096 92452 5100 92508
rect 5036 92448 5100 92452
rect 5116 92508 5180 92512
rect 5116 92452 5120 92508
rect 5120 92452 5176 92508
rect 5176 92452 5180 92508
rect 5116 92448 5180 92452
rect 106660 92508 106724 92512
rect 106660 92452 106664 92508
rect 106664 92452 106720 92508
rect 106720 92452 106724 92508
rect 106660 92448 106724 92452
rect 106740 92508 106804 92512
rect 106740 92452 106744 92508
rect 106744 92452 106800 92508
rect 106800 92452 106804 92508
rect 106740 92448 106804 92452
rect 106820 92508 106884 92512
rect 106820 92452 106824 92508
rect 106824 92452 106880 92508
rect 106880 92452 106884 92508
rect 106820 92448 106884 92452
rect 106900 92508 106964 92512
rect 106900 92452 106904 92508
rect 106904 92452 106960 92508
rect 106960 92452 106964 92508
rect 106900 92448 106964 92452
rect 4216 91964 4280 91968
rect 4216 91908 4220 91964
rect 4220 91908 4276 91964
rect 4276 91908 4280 91964
rect 4216 91904 4280 91908
rect 4296 91964 4360 91968
rect 4296 91908 4300 91964
rect 4300 91908 4356 91964
rect 4356 91908 4360 91964
rect 4296 91904 4360 91908
rect 4376 91964 4440 91968
rect 4376 91908 4380 91964
rect 4380 91908 4436 91964
rect 4436 91908 4440 91964
rect 4376 91904 4440 91908
rect 4456 91964 4520 91968
rect 4456 91908 4460 91964
rect 4460 91908 4516 91964
rect 4516 91908 4520 91964
rect 4456 91904 4520 91908
rect 105924 91964 105988 91968
rect 105924 91908 105928 91964
rect 105928 91908 105984 91964
rect 105984 91908 105988 91964
rect 105924 91904 105988 91908
rect 106004 91964 106068 91968
rect 106004 91908 106008 91964
rect 106008 91908 106064 91964
rect 106064 91908 106068 91964
rect 106004 91904 106068 91908
rect 106084 91964 106148 91968
rect 106084 91908 106088 91964
rect 106088 91908 106144 91964
rect 106144 91908 106148 91964
rect 106084 91904 106148 91908
rect 106164 91964 106228 91968
rect 106164 91908 106168 91964
rect 106168 91908 106224 91964
rect 106224 91908 106228 91964
rect 106164 91904 106228 91908
rect 4876 91420 4940 91424
rect 4876 91364 4880 91420
rect 4880 91364 4936 91420
rect 4936 91364 4940 91420
rect 4876 91360 4940 91364
rect 4956 91420 5020 91424
rect 4956 91364 4960 91420
rect 4960 91364 5016 91420
rect 5016 91364 5020 91420
rect 4956 91360 5020 91364
rect 5036 91420 5100 91424
rect 5036 91364 5040 91420
rect 5040 91364 5096 91420
rect 5096 91364 5100 91420
rect 5036 91360 5100 91364
rect 5116 91420 5180 91424
rect 5116 91364 5120 91420
rect 5120 91364 5176 91420
rect 5176 91364 5180 91420
rect 5116 91360 5180 91364
rect 106660 91420 106724 91424
rect 106660 91364 106664 91420
rect 106664 91364 106720 91420
rect 106720 91364 106724 91420
rect 106660 91360 106724 91364
rect 106740 91420 106804 91424
rect 106740 91364 106744 91420
rect 106744 91364 106800 91420
rect 106800 91364 106804 91420
rect 106740 91360 106804 91364
rect 106820 91420 106884 91424
rect 106820 91364 106824 91420
rect 106824 91364 106880 91420
rect 106880 91364 106884 91420
rect 106820 91360 106884 91364
rect 106900 91420 106964 91424
rect 106900 91364 106904 91420
rect 106904 91364 106960 91420
rect 106960 91364 106964 91420
rect 106900 91360 106964 91364
rect 4216 90876 4280 90880
rect 4216 90820 4220 90876
rect 4220 90820 4276 90876
rect 4276 90820 4280 90876
rect 4216 90816 4280 90820
rect 4296 90876 4360 90880
rect 4296 90820 4300 90876
rect 4300 90820 4356 90876
rect 4356 90820 4360 90876
rect 4296 90816 4360 90820
rect 4376 90876 4440 90880
rect 4376 90820 4380 90876
rect 4380 90820 4436 90876
rect 4436 90820 4440 90876
rect 4376 90816 4440 90820
rect 4456 90876 4520 90880
rect 4456 90820 4460 90876
rect 4460 90820 4516 90876
rect 4516 90820 4520 90876
rect 4456 90816 4520 90820
rect 105924 90876 105988 90880
rect 105924 90820 105928 90876
rect 105928 90820 105984 90876
rect 105984 90820 105988 90876
rect 105924 90816 105988 90820
rect 106004 90876 106068 90880
rect 106004 90820 106008 90876
rect 106008 90820 106064 90876
rect 106064 90820 106068 90876
rect 106004 90816 106068 90820
rect 106084 90876 106148 90880
rect 106084 90820 106088 90876
rect 106088 90820 106144 90876
rect 106144 90820 106148 90876
rect 106084 90816 106148 90820
rect 106164 90876 106228 90880
rect 106164 90820 106168 90876
rect 106168 90820 106224 90876
rect 106224 90820 106228 90876
rect 106164 90816 106228 90820
rect 4876 90332 4940 90336
rect 4876 90276 4880 90332
rect 4880 90276 4936 90332
rect 4936 90276 4940 90332
rect 4876 90272 4940 90276
rect 4956 90332 5020 90336
rect 4956 90276 4960 90332
rect 4960 90276 5016 90332
rect 5016 90276 5020 90332
rect 4956 90272 5020 90276
rect 5036 90332 5100 90336
rect 5036 90276 5040 90332
rect 5040 90276 5096 90332
rect 5096 90276 5100 90332
rect 5036 90272 5100 90276
rect 5116 90332 5180 90336
rect 5116 90276 5120 90332
rect 5120 90276 5176 90332
rect 5176 90276 5180 90332
rect 5116 90272 5180 90276
rect 106660 90332 106724 90336
rect 106660 90276 106664 90332
rect 106664 90276 106720 90332
rect 106720 90276 106724 90332
rect 106660 90272 106724 90276
rect 106740 90332 106804 90336
rect 106740 90276 106744 90332
rect 106744 90276 106800 90332
rect 106800 90276 106804 90332
rect 106740 90272 106804 90276
rect 106820 90332 106884 90336
rect 106820 90276 106824 90332
rect 106824 90276 106880 90332
rect 106880 90276 106884 90332
rect 106820 90272 106884 90276
rect 106900 90332 106964 90336
rect 106900 90276 106904 90332
rect 106904 90276 106960 90332
rect 106960 90276 106964 90332
rect 106900 90272 106964 90276
rect 4216 89788 4280 89792
rect 4216 89732 4220 89788
rect 4220 89732 4276 89788
rect 4276 89732 4280 89788
rect 4216 89728 4280 89732
rect 4296 89788 4360 89792
rect 4296 89732 4300 89788
rect 4300 89732 4356 89788
rect 4356 89732 4360 89788
rect 4296 89728 4360 89732
rect 4376 89788 4440 89792
rect 4376 89732 4380 89788
rect 4380 89732 4436 89788
rect 4436 89732 4440 89788
rect 4376 89728 4440 89732
rect 4456 89788 4520 89792
rect 4456 89732 4460 89788
rect 4460 89732 4516 89788
rect 4516 89732 4520 89788
rect 4456 89728 4520 89732
rect 105924 89788 105988 89792
rect 105924 89732 105928 89788
rect 105928 89732 105984 89788
rect 105984 89732 105988 89788
rect 105924 89728 105988 89732
rect 106004 89788 106068 89792
rect 106004 89732 106008 89788
rect 106008 89732 106064 89788
rect 106064 89732 106068 89788
rect 106004 89728 106068 89732
rect 106084 89788 106148 89792
rect 106084 89732 106088 89788
rect 106088 89732 106144 89788
rect 106144 89732 106148 89788
rect 106084 89728 106148 89732
rect 106164 89788 106228 89792
rect 106164 89732 106168 89788
rect 106168 89732 106224 89788
rect 106224 89732 106228 89788
rect 106164 89728 106228 89732
rect 4876 89244 4940 89248
rect 4876 89188 4880 89244
rect 4880 89188 4936 89244
rect 4936 89188 4940 89244
rect 4876 89184 4940 89188
rect 4956 89244 5020 89248
rect 4956 89188 4960 89244
rect 4960 89188 5016 89244
rect 5016 89188 5020 89244
rect 4956 89184 5020 89188
rect 5036 89244 5100 89248
rect 5036 89188 5040 89244
rect 5040 89188 5096 89244
rect 5096 89188 5100 89244
rect 5036 89184 5100 89188
rect 5116 89244 5180 89248
rect 5116 89188 5120 89244
rect 5120 89188 5176 89244
rect 5176 89188 5180 89244
rect 5116 89184 5180 89188
rect 106660 89244 106724 89248
rect 106660 89188 106664 89244
rect 106664 89188 106720 89244
rect 106720 89188 106724 89244
rect 106660 89184 106724 89188
rect 106740 89244 106804 89248
rect 106740 89188 106744 89244
rect 106744 89188 106800 89244
rect 106800 89188 106804 89244
rect 106740 89184 106804 89188
rect 106820 89244 106884 89248
rect 106820 89188 106824 89244
rect 106824 89188 106880 89244
rect 106880 89188 106884 89244
rect 106820 89184 106884 89188
rect 106900 89244 106964 89248
rect 106900 89188 106904 89244
rect 106904 89188 106960 89244
rect 106960 89188 106964 89244
rect 106900 89184 106964 89188
rect 4216 88700 4280 88704
rect 4216 88644 4220 88700
rect 4220 88644 4276 88700
rect 4276 88644 4280 88700
rect 4216 88640 4280 88644
rect 4296 88700 4360 88704
rect 4296 88644 4300 88700
rect 4300 88644 4356 88700
rect 4356 88644 4360 88700
rect 4296 88640 4360 88644
rect 4376 88700 4440 88704
rect 4376 88644 4380 88700
rect 4380 88644 4436 88700
rect 4436 88644 4440 88700
rect 4376 88640 4440 88644
rect 4456 88700 4520 88704
rect 4456 88644 4460 88700
rect 4460 88644 4516 88700
rect 4516 88644 4520 88700
rect 4456 88640 4520 88644
rect 105924 88700 105988 88704
rect 105924 88644 105928 88700
rect 105928 88644 105984 88700
rect 105984 88644 105988 88700
rect 105924 88640 105988 88644
rect 106004 88700 106068 88704
rect 106004 88644 106008 88700
rect 106008 88644 106064 88700
rect 106064 88644 106068 88700
rect 106004 88640 106068 88644
rect 106084 88700 106148 88704
rect 106084 88644 106088 88700
rect 106088 88644 106144 88700
rect 106144 88644 106148 88700
rect 106084 88640 106148 88644
rect 106164 88700 106228 88704
rect 106164 88644 106168 88700
rect 106168 88644 106224 88700
rect 106224 88644 106228 88700
rect 106164 88640 106228 88644
rect 4876 88156 4940 88160
rect 4876 88100 4880 88156
rect 4880 88100 4936 88156
rect 4936 88100 4940 88156
rect 4876 88096 4940 88100
rect 4956 88156 5020 88160
rect 4956 88100 4960 88156
rect 4960 88100 5016 88156
rect 5016 88100 5020 88156
rect 4956 88096 5020 88100
rect 5036 88156 5100 88160
rect 5036 88100 5040 88156
rect 5040 88100 5096 88156
rect 5096 88100 5100 88156
rect 5036 88096 5100 88100
rect 5116 88156 5180 88160
rect 5116 88100 5120 88156
rect 5120 88100 5176 88156
rect 5176 88100 5180 88156
rect 5116 88096 5180 88100
rect 106660 88156 106724 88160
rect 106660 88100 106664 88156
rect 106664 88100 106720 88156
rect 106720 88100 106724 88156
rect 106660 88096 106724 88100
rect 106740 88156 106804 88160
rect 106740 88100 106744 88156
rect 106744 88100 106800 88156
rect 106800 88100 106804 88156
rect 106740 88096 106804 88100
rect 106820 88156 106884 88160
rect 106820 88100 106824 88156
rect 106824 88100 106880 88156
rect 106880 88100 106884 88156
rect 106820 88096 106884 88100
rect 106900 88156 106964 88160
rect 106900 88100 106904 88156
rect 106904 88100 106960 88156
rect 106960 88100 106964 88156
rect 106900 88096 106964 88100
rect 4216 87612 4280 87616
rect 4216 87556 4220 87612
rect 4220 87556 4276 87612
rect 4276 87556 4280 87612
rect 4216 87552 4280 87556
rect 4296 87612 4360 87616
rect 4296 87556 4300 87612
rect 4300 87556 4356 87612
rect 4356 87556 4360 87612
rect 4296 87552 4360 87556
rect 4376 87612 4440 87616
rect 4376 87556 4380 87612
rect 4380 87556 4436 87612
rect 4436 87556 4440 87612
rect 4376 87552 4440 87556
rect 4456 87612 4520 87616
rect 4456 87556 4460 87612
rect 4460 87556 4516 87612
rect 4516 87556 4520 87612
rect 4456 87552 4520 87556
rect 105924 87612 105988 87616
rect 105924 87556 105928 87612
rect 105928 87556 105984 87612
rect 105984 87556 105988 87612
rect 105924 87552 105988 87556
rect 106004 87612 106068 87616
rect 106004 87556 106008 87612
rect 106008 87556 106064 87612
rect 106064 87556 106068 87612
rect 106004 87552 106068 87556
rect 106084 87612 106148 87616
rect 106084 87556 106088 87612
rect 106088 87556 106144 87612
rect 106144 87556 106148 87612
rect 106084 87552 106148 87556
rect 106164 87612 106228 87616
rect 106164 87556 106168 87612
rect 106168 87556 106224 87612
rect 106224 87556 106228 87612
rect 106164 87552 106228 87556
rect 4876 87068 4940 87072
rect 4876 87012 4880 87068
rect 4880 87012 4936 87068
rect 4936 87012 4940 87068
rect 4876 87008 4940 87012
rect 4956 87068 5020 87072
rect 4956 87012 4960 87068
rect 4960 87012 5016 87068
rect 5016 87012 5020 87068
rect 4956 87008 5020 87012
rect 5036 87068 5100 87072
rect 5036 87012 5040 87068
rect 5040 87012 5096 87068
rect 5096 87012 5100 87068
rect 5036 87008 5100 87012
rect 5116 87068 5180 87072
rect 5116 87012 5120 87068
rect 5120 87012 5176 87068
rect 5176 87012 5180 87068
rect 5116 87008 5180 87012
rect 106660 87068 106724 87072
rect 106660 87012 106664 87068
rect 106664 87012 106720 87068
rect 106720 87012 106724 87068
rect 106660 87008 106724 87012
rect 106740 87068 106804 87072
rect 106740 87012 106744 87068
rect 106744 87012 106800 87068
rect 106800 87012 106804 87068
rect 106740 87008 106804 87012
rect 106820 87068 106884 87072
rect 106820 87012 106824 87068
rect 106824 87012 106880 87068
rect 106880 87012 106884 87068
rect 106820 87008 106884 87012
rect 106900 87068 106964 87072
rect 106900 87012 106904 87068
rect 106904 87012 106960 87068
rect 106960 87012 106964 87068
rect 106900 87008 106964 87012
rect 4216 86524 4280 86528
rect 4216 86468 4220 86524
rect 4220 86468 4276 86524
rect 4276 86468 4280 86524
rect 4216 86464 4280 86468
rect 4296 86524 4360 86528
rect 4296 86468 4300 86524
rect 4300 86468 4356 86524
rect 4356 86468 4360 86524
rect 4296 86464 4360 86468
rect 4376 86524 4440 86528
rect 4376 86468 4380 86524
rect 4380 86468 4436 86524
rect 4436 86468 4440 86524
rect 4376 86464 4440 86468
rect 4456 86524 4520 86528
rect 4456 86468 4460 86524
rect 4460 86468 4516 86524
rect 4516 86468 4520 86524
rect 4456 86464 4520 86468
rect 105924 86524 105988 86528
rect 105924 86468 105928 86524
rect 105928 86468 105984 86524
rect 105984 86468 105988 86524
rect 105924 86464 105988 86468
rect 106004 86524 106068 86528
rect 106004 86468 106008 86524
rect 106008 86468 106064 86524
rect 106064 86468 106068 86524
rect 106004 86464 106068 86468
rect 106084 86524 106148 86528
rect 106084 86468 106088 86524
rect 106088 86468 106144 86524
rect 106144 86468 106148 86524
rect 106084 86464 106148 86468
rect 106164 86524 106228 86528
rect 106164 86468 106168 86524
rect 106168 86468 106224 86524
rect 106224 86468 106228 86524
rect 106164 86464 106228 86468
rect 4876 85980 4940 85984
rect 4876 85924 4880 85980
rect 4880 85924 4936 85980
rect 4936 85924 4940 85980
rect 4876 85920 4940 85924
rect 4956 85980 5020 85984
rect 4956 85924 4960 85980
rect 4960 85924 5016 85980
rect 5016 85924 5020 85980
rect 4956 85920 5020 85924
rect 5036 85980 5100 85984
rect 5036 85924 5040 85980
rect 5040 85924 5096 85980
rect 5096 85924 5100 85980
rect 5036 85920 5100 85924
rect 5116 85980 5180 85984
rect 5116 85924 5120 85980
rect 5120 85924 5176 85980
rect 5176 85924 5180 85980
rect 5116 85920 5180 85924
rect 106660 85980 106724 85984
rect 106660 85924 106664 85980
rect 106664 85924 106720 85980
rect 106720 85924 106724 85980
rect 106660 85920 106724 85924
rect 106740 85980 106804 85984
rect 106740 85924 106744 85980
rect 106744 85924 106800 85980
rect 106800 85924 106804 85980
rect 106740 85920 106804 85924
rect 106820 85980 106884 85984
rect 106820 85924 106824 85980
rect 106824 85924 106880 85980
rect 106880 85924 106884 85980
rect 106820 85920 106884 85924
rect 106900 85980 106964 85984
rect 106900 85924 106904 85980
rect 106904 85924 106960 85980
rect 106960 85924 106964 85980
rect 106900 85920 106964 85924
rect 4216 85436 4280 85440
rect 4216 85380 4220 85436
rect 4220 85380 4276 85436
rect 4276 85380 4280 85436
rect 4216 85376 4280 85380
rect 4296 85436 4360 85440
rect 4296 85380 4300 85436
rect 4300 85380 4356 85436
rect 4356 85380 4360 85436
rect 4296 85376 4360 85380
rect 4376 85436 4440 85440
rect 4376 85380 4380 85436
rect 4380 85380 4436 85436
rect 4436 85380 4440 85436
rect 4376 85376 4440 85380
rect 4456 85436 4520 85440
rect 4456 85380 4460 85436
rect 4460 85380 4516 85436
rect 4516 85380 4520 85436
rect 4456 85376 4520 85380
rect 105924 85436 105988 85440
rect 105924 85380 105928 85436
rect 105928 85380 105984 85436
rect 105984 85380 105988 85436
rect 105924 85376 105988 85380
rect 106004 85436 106068 85440
rect 106004 85380 106008 85436
rect 106008 85380 106064 85436
rect 106064 85380 106068 85436
rect 106004 85376 106068 85380
rect 106084 85436 106148 85440
rect 106084 85380 106088 85436
rect 106088 85380 106144 85436
rect 106144 85380 106148 85436
rect 106084 85376 106148 85380
rect 106164 85436 106228 85440
rect 106164 85380 106168 85436
rect 106168 85380 106224 85436
rect 106224 85380 106228 85436
rect 106164 85376 106228 85380
rect 4876 84892 4940 84896
rect 4876 84836 4880 84892
rect 4880 84836 4936 84892
rect 4936 84836 4940 84892
rect 4876 84832 4940 84836
rect 4956 84892 5020 84896
rect 4956 84836 4960 84892
rect 4960 84836 5016 84892
rect 5016 84836 5020 84892
rect 4956 84832 5020 84836
rect 5036 84892 5100 84896
rect 5036 84836 5040 84892
rect 5040 84836 5096 84892
rect 5096 84836 5100 84892
rect 5036 84832 5100 84836
rect 5116 84892 5180 84896
rect 5116 84836 5120 84892
rect 5120 84836 5176 84892
rect 5176 84836 5180 84892
rect 5116 84832 5180 84836
rect 106660 84892 106724 84896
rect 106660 84836 106664 84892
rect 106664 84836 106720 84892
rect 106720 84836 106724 84892
rect 106660 84832 106724 84836
rect 106740 84892 106804 84896
rect 106740 84836 106744 84892
rect 106744 84836 106800 84892
rect 106800 84836 106804 84892
rect 106740 84832 106804 84836
rect 106820 84892 106884 84896
rect 106820 84836 106824 84892
rect 106824 84836 106880 84892
rect 106880 84836 106884 84892
rect 106820 84832 106884 84836
rect 106900 84892 106964 84896
rect 106900 84836 106904 84892
rect 106904 84836 106960 84892
rect 106960 84836 106964 84892
rect 106900 84832 106964 84836
rect 4216 84348 4280 84352
rect 4216 84292 4220 84348
rect 4220 84292 4276 84348
rect 4276 84292 4280 84348
rect 4216 84288 4280 84292
rect 4296 84348 4360 84352
rect 4296 84292 4300 84348
rect 4300 84292 4356 84348
rect 4356 84292 4360 84348
rect 4296 84288 4360 84292
rect 4376 84348 4440 84352
rect 4376 84292 4380 84348
rect 4380 84292 4436 84348
rect 4436 84292 4440 84348
rect 4376 84288 4440 84292
rect 4456 84348 4520 84352
rect 4456 84292 4460 84348
rect 4460 84292 4516 84348
rect 4516 84292 4520 84348
rect 4456 84288 4520 84292
rect 105924 84348 105988 84352
rect 105924 84292 105928 84348
rect 105928 84292 105984 84348
rect 105984 84292 105988 84348
rect 105924 84288 105988 84292
rect 106004 84348 106068 84352
rect 106004 84292 106008 84348
rect 106008 84292 106064 84348
rect 106064 84292 106068 84348
rect 106004 84288 106068 84292
rect 106084 84348 106148 84352
rect 106084 84292 106088 84348
rect 106088 84292 106144 84348
rect 106144 84292 106148 84348
rect 106084 84288 106148 84292
rect 106164 84348 106228 84352
rect 106164 84292 106168 84348
rect 106168 84292 106224 84348
rect 106224 84292 106228 84348
rect 106164 84288 106228 84292
rect 4876 83804 4940 83808
rect 4876 83748 4880 83804
rect 4880 83748 4936 83804
rect 4936 83748 4940 83804
rect 4876 83744 4940 83748
rect 4956 83804 5020 83808
rect 4956 83748 4960 83804
rect 4960 83748 5016 83804
rect 5016 83748 5020 83804
rect 4956 83744 5020 83748
rect 5036 83804 5100 83808
rect 5036 83748 5040 83804
rect 5040 83748 5096 83804
rect 5096 83748 5100 83804
rect 5036 83744 5100 83748
rect 5116 83804 5180 83808
rect 5116 83748 5120 83804
rect 5120 83748 5176 83804
rect 5176 83748 5180 83804
rect 5116 83744 5180 83748
rect 106660 83804 106724 83808
rect 106660 83748 106664 83804
rect 106664 83748 106720 83804
rect 106720 83748 106724 83804
rect 106660 83744 106724 83748
rect 106740 83804 106804 83808
rect 106740 83748 106744 83804
rect 106744 83748 106800 83804
rect 106800 83748 106804 83804
rect 106740 83744 106804 83748
rect 106820 83804 106884 83808
rect 106820 83748 106824 83804
rect 106824 83748 106880 83804
rect 106880 83748 106884 83804
rect 106820 83744 106884 83748
rect 106900 83804 106964 83808
rect 106900 83748 106904 83804
rect 106904 83748 106960 83804
rect 106960 83748 106964 83804
rect 106900 83744 106964 83748
rect 4216 83260 4280 83264
rect 4216 83204 4220 83260
rect 4220 83204 4276 83260
rect 4276 83204 4280 83260
rect 4216 83200 4280 83204
rect 4296 83260 4360 83264
rect 4296 83204 4300 83260
rect 4300 83204 4356 83260
rect 4356 83204 4360 83260
rect 4296 83200 4360 83204
rect 4376 83260 4440 83264
rect 4376 83204 4380 83260
rect 4380 83204 4436 83260
rect 4436 83204 4440 83260
rect 4376 83200 4440 83204
rect 4456 83260 4520 83264
rect 4456 83204 4460 83260
rect 4460 83204 4516 83260
rect 4516 83204 4520 83260
rect 4456 83200 4520 83204
rect 105924 83260 105988 83264
rect 105924 83204 105928 83260
rect 105928 83204 105984 83260
rect 105984 83204 105988 83260
rect 105924 83200 105988 83204
rect 106004 83260 106068 83264
rect 106004 83204 106008 83260
rect 106008 83204 106064 83260
rect 106064 83204 106068 83260
rect 106004 83200 106068 83204
rect 106084 83260 106148 83264
rect 106084 83204 106088 83260
rect 106088 83204 106144 83260
rect 106144 83204 106148 83260
rect 106084 83200 106148 83204
rect 106164 83260 106228 83264
rect 106164 83204 106168 83260
rect 106168 83204 106224 83260
rect 106224 83204 106228 83260
rect 106164 83200 106228 83204
rect 4876 82716 4940 82720
rect 4876 82660 4880 82716
rect 4880 82660 4936 82716
rect 4936 82660 4940 82716
rect 4876 82656 4940 82660
rect 4956 82716 5020 82720
rect 4956 82660 4960 82716
rect 4960 82660 5016 82716
rect 5016 82660 5020 82716
rect 4956 82656 5020 82660
rect 5036 82716 5100 82720
rect 5036 82660 5040 82716
rect 5040 82660 5096 82716
rect 5096 82660 5100 82716
rect 5036 82656 5100 82660
rect 5116 82716 5180 82720
rect 5116 82660 5120 82716
rect 5120 82660 5176 82716
rect 5176 82660 5180 82716
rect 5116 82656 5180 82660
rect 106660 82716 106724 82720
rect 106660 82660 106664 82716
rect 106664 82660 106720 82716
rect 106720 82660 106724 82716
rect 106660 82656 106724 82660
rect 106740 82716 106804 82720
rect 106740 82660 106744 82716
rect 106744 82660 106800 82716
rect 106800 82660 106804 82716
rect 106740 82656 106804 82660
rect 106820 82716 106884 82720
rect 106820 82660 106824 82716
rect 106824 82660 106880 82716
rect 106880 82660 106884 82716
rect 106820 82656 106884 82660
rect 106900 82716 106964 82720
rect 106900 82660 106904 82716
rect 106904 82660 106960 82716
rect 106960 82660 106964 82716
rect 106900 82656 106964 82660
rect 4216 82172 4280 82176
rect 4216 82116 4220 82172
rect 4220 82116 4276 82172
rect 4276 82116 4280 82172
rect 4216 82112 4280 82116
rect 4296 82172 4360 82176
rect 4296 82116 4300 82172
rect 4300 82116 4356 82172
rect 4356 82116 4360 82172
rect 4296 82112 4360 82116
rect 4376 82172 4440 82176
rect 4376 82116 4380 82172
rect 4380 82116 4436 82172
rect 4436 82116 4440 82172
rect 4376 82112 4440 82116
rect 4456 82172 4520 82176
rect 4456 82116 4460 82172
rect 4460 82116 4516 82172
rect 4516 82116 4520 82172
rect 4456 82112 4520 82116
rect 105924 82172 105988 82176
rect 105924 82116 105928 82172
rect 105928 82116 105984 82172
rect 105984 82116 105988 82172
rect 105924 82112 105988 82116
rect 106004 82172 106068 82176
rect 106004 82116 106008 82172
rect 106008 82116 106064 82172
rect 106064 82116 106068 82172
rect 106004 82112 106068 82116
rect 106084 82172 106148 82176
rect 106084 82116 106088 82172
rect 106088 82116 106144 82172
rect 106144 82116 106148 82172
rect 106084 82112 106148 82116
rect 106164 82172 106228 82176
rect 106164 82116 106168 82172
rect 106168 82116 106224 82172
rect 106224 82116 106228 82172
rect 106164 82112 106228 82116
rect 4876 81628 4940 81632
rect 4876 81572 4880 81628
rect 4880 81572 4936 81628
rect 4936 81572 4940 81628
rect 4876 81568 4940 81572
rect 4956 81628 5020 81632
rect 4956 81572 4960 81628
rect 4960 81572 5016 81628
rect 5016 81572 5020 81628
rect 4956 81568 5020 81572
rect 5036 81628 5100 81632
rect 5036 81572 5040 81628
rect 5040 81572 5096 81628
rect 5096 81572 5100 81628
rect 5036 81568 5100 81572
rect 5116 81628 5180 81632
rect 5116 81572 5120 81628
rect 5120 81572 5176 81628
rect 5176 81572 5180 81628
rect 5116 81568 5180 81572
rect 106660 81628 106724 81632
rect 106660 81572 106664 81628
rect 106664 81572 106720 81628
rect 106720 81572 106724 81628
rect 106660 81568 106724 81572
rect 106740 81628 106804 81632
rect 106740 81572 106744 81628
rect 106744 81572 106800 81628
rect 106800 81572 106804 81628
rect 106740 81568 106804 81572
rect 106820 81628 106884 81632
rect 106820 81572 106824 81628
rect 106824 81572 106880 81628
rect 106880 81572 106884 81628
rect 106820 81568 106884 81572
rect 106900 81628 106964 81632
rect 106900 81572 106904 81628
rect 106904 81572 106960 81628
rect 106960 81572 106964 81628
rect 106900 81568 106964 81572
rect 4216 81084 4280 81088
rect 4216 81028 4220 81084
rect 4220 81028 4276 81084
rect 4276 81028 4280 81084
rect 4216 81024 4280 81028
rect 4296 81084 4360 81088
rect 4296 81028 4300 81084
rect 4300 81028 4356 81084
rect 4356 81028 4360 81084
rect 4296 81024 4360 81028
rect 4376 81084 4440 81088
rect 4376 81028 4380 81084
rect 4380 81028 4436 81084
rect 4436 81028 4440 81084
rect 4376 81024 4440 81028
rect 4456 81084 4520 81088
rect 4456 81028 4460 81084
rect 4460 81028 4516 81084
rect 4516 81028 4520 81084
rect 4456 81024 4520 81028
rect 105924 81084 105988 81088
rect 105924 81028 105928 81084
rect 105928 81028 105984 81084
rect 105984 81028 105988 81084
rect 105924 81024 105988 81028
rect 106004 81084 106068 81088
rect 106004 81028 106008 81084
rect 106008 81028 106064 81084
rect 106064 81028 106068 81084
rect 106004 81024 106068 81028
rect 106084 81084 106148 81088
rect 106084 81028 106088 81084
rect 106088 81028 106144 81084
rect 106144 81028 106148 81084
rect 106084 81024 106148 81028
rect 106164 81084 106228 81088
rect 106164 81028 106168 81084
rect 106168 81028 106224 81084
rect 106224 81028 106228 81084
rect 106164 81024 106228 81028
rect 4876 80540 4940 80544
rect 4876 80484 4880 80540
rect 4880 80484 4936 80540
rect 4936 80484 4940 80540
rect 4876 80480 4940 80484
rect 4956 80540 5020 80544
rect 4956 80484 4960 80540
rect 4960 80484 5016 80540
rect 5016 80484 5020 80540
rect 4956 80480 5020 80484
rect 5036 80540 5100 80544
rect 5036 80484 5040 80540
rect 5040 80484 5096 80540
rect 5096 80484 5100 80540
rect 5036 80480 5100 80484
rect 5116 80540 5180 80544
rect 5116 80484 5120 80540
rect 5120 80484 5176 80540
rect 5176 80484 5180 80540
rect 5116 80480 5180 80484
rect 106660 80540 106724 80544
rect 106660 80484 106664 80540
rect 106664 80484 106720 80540
rect 106720 80484 106724 80540
rect 106660 80480 106724 80484
rect 106740 80540 106804 80544
rect 106740 80484 106744 80540
rect 106744 80484 106800 80540
rect 106800 80484 106804 80540
rect 106740 80480 106804 80484
rect 106820 80540 106884 80544
rect 106820 80484 106824 80540
rect 106824 80484 106880 80540
rect 106880 80484 106884 80540
rect 106820 80480 106884 80484
rect 106900 80540 106964 80544
rect 106900 80484 106904 80540
rect 106904 80484 106960 80540
rect 106960 80484 106964 80540
rect 106900 80480 106964 80484
rect 4216 79996 4280 80000
rect 4216 79940 4220 79996
rect 4220 79940 4276 79996
rect 4276 79940 4280 79996
rect 4216 79936 4280 79940
rect 4296 79996 4360 80000
rect 4296 79940 4300 79996
rect 4300 79940 4356 79996
rect 4356 79940 4360 79996
rect 4296 79936 4360 79940
rect 4376 79996 4440 80000
rect 4376 79940 4380 79996
rect 4380 79940 4436 79996
rect 4436 79940 4440 79996
rect 4376 79936 4440 79940
rect 4456 79996 4520 80000
rect 4456 79940 4460 79996
rect 4460 79940 4516 79996
rect 4516 79940 4520 79996
rect 4456 79936 4520 79940
rect 105924 79996 105988 80000
rect 105924 79940 105928 79996
rect 105928 79940 105984 79996
rect 105984 79940 105988 79996
rect 105924 79936 105988 79940
rect 106004 79996 106068 80000
rect 106004 79940 106008 79996
rect 106008 79940 106064 79996
rect 106064 79940 106068 79996
rect 106004 79936 106068 79940
rect 106084 79996 106148 80000
rect 106084 79940 106088 79996
rect 106088 79940 106144 79996
rect 106144 79940 106148 79996
rect 106084 79936 106148 79940
rect 106164 79996 106228 80000
rect 106164 79940 106168 79996
rect 106168 79940 106224 79996
rect 106224 79940 106228 79996
rect 106164 79936 106228 79940
rect 4876 79452 4940 79456
rect 4876 79396 4880 79452
rect 4880 79396 4936 79452
rect 4936 79396 4940 79452
rect 4876 79392 4940 79396
rect 4956 79452 5020 79456
rect 4956 79396 4960 79452
rect 4960 79396 5016 79452
rect 5016 79396 5020 79452
rect 4956 79392 5020 79396
rect 5036 79452 5100 79456
rect 5036 79396 5040 79452
rect 5040 79396 5096 79452
rect 5096 79396 5100 79452
rect 5036 79392 5100 79396
rect 5116 79452 5180 79456
rect 5116 79396 5120 79452
rect 5120 79396 5176 79452
rect 5176 79396 5180 79452
rect 5116 79392 5180 79396
rect 106660 79452 106724 79456
rect 106660 79396 106664 79452
rect 106664 79396 106720 79452
rect 106720 79396 106724 79452
rect 106660 79392 106724 79396
rect 106740 79452 106804 79456
rect 106740 79396 106744 79452
rect 106744 79396 106800 79452
rect 106800 79396 106804 79452
rect 106740 79392 106804 79396
rect 106820 79452 106884 79456
rect 106820 79396 106824 79452
rect 106824 79396 106880 79452
rect 106880 79396 106884 79452
rect 106820 79392 106884 79396
rect 106900 79452 106964 79456
rect 106900 79396 106904 79452
rect 106904 79396 106960 79452
rect 106960 79396 106964 79452
rect 106900 79392 106964 79396
rect 4216 78908 4280 78912
rect 4216 78852 4220 78908
rect 4220 78852 4276 78908
rect 4276 78852 4280 78908
rect 4216 78848 4280 78852
rect 4296 78908 4360 78912
rect 4296 78852 4300 78908
rect 4300 78852 4356 78908
rect 4356 78852 4360 78908
rect 4296 78848 4360 78852
rect 4376 78908 4440 78912
rect 4376 78852 4380 78908
rect 4380 78852 4436 78908
rect 4436 78852 4440 78908
rect 4376 78848 4440 78852
rect 4456 78908 4520 78912
rect 4456 78852 4460 78908
rect 4460 78852 4516 78908
rect 4516 78852 4520 78908
rect 4456 78848 4520 78852
rect 105924 78908 105988 78912
rect 105924 78852 105928 78908
rect 105928 78852 105984 78908
rect 105984 78852 105988 78908
rect 105924 78848 105988 78852
rect 106004 78908 106068 78912
rect 106004 78852 106008 78908
rect 106008 78852 106064 78908
rect 106064 78852 106068 78908
rect 106004 78848 106068 78852
rect 106084 78908 106148 78912
rect 106084 78852 106088 78908
rect 106088 78852 106144 78908
rect 106144 78852 106148 78908
rect 106084 78848 106148 78852
rect 106164 78908 106228 78912
rect 106164 78852 106168 78908
rect 106168 78852 106224 78908
rect 106224 78852 106228 78908
rect 106164 78848 106228 78852
rect 4876 78364 4940 78368
rect 4876 78308 4880 78364
rect 4880 78308 4936 78364
rect 4936 78308 4940 78364
rect 4876 78304 4940 78308
rect 4956 78364 5020 78368
rect 4956 78308 4960 78364
rect 4960 78308 5016 78364
rect 5016 78308 5020 78364
rect 4956 78304 5020 78308
rect 5036 78364 5100 78368
rect 5036 78308 5040 78364
rect 5040 78308 5096 78364
rect 5096 78308 5100 78364
rect 5036 78304 5100 78308
rect 5116 78364 5180 78368
rect 5116 78308 5120 78364
rect 5120 78308 5176 78364
rect 5176 78308 5180 78364
rect 5116 78304 5180 78308
rect 106660 78364 106724 78368
rect 106660 78308 106664 78364
rect 106664 78308 106720 78364
rect 106720 78308 106724 78364
rect 106660 78304 106724 78308
rect 106740 78364 106804 78368
rect 106740 78308 106744 78364
rect 106744 78308 106800 78364
rect 106800 78308 106804 78364
rect 106740 78304 106804 78308
rect 106820 78364 106884 78368
rect 106820 78308 106824 78364
rect 106824 78308 106880 78364
rect 106880 78308 106884 78364
rect 106820 78304 106884 78308
rect 106900 78364 106964 78368
rect 106900 78308 106904 78364
rect 106904 78308 106960 78364
rect 106960 78308 106964 78364
rect 106900 78304 106964 78308
rect 4216 77820 4280 77824
rect 4216 77764 4220 77820
rect 4220 77764 4276 77820
rect 4276 77764 4280 77820
rect 4216 77760 4280 77764
rect 4296 77820 4360 77824
rect 4296 77764 4300 77820
rect 4300 77764 4356 77820
rect 4356 77764 4360 77820
rect 4296 77760 4360 77764
rect 4376 77820 4440 77824
rect 4376 77764 4380 77820
rect 4380 77764 4436 77820
rect 4436 77764 4440 77820
rect 4376 77760 4440 77764
rect 4456 77820 4520 77824
rect 4456 77764 4460 77820
rect 4460 77764 4516 77820
rect 4516 77764 4520 77820
rect 4456 77760 4520 77764
rect 105924 77820 105988 77824
rect 105924 77764 105928 77820
rect 105928 77764 105984 77820
rect 105984 77764 105988 77820
rect 105924 77760 105988 77764
rect 106004 77820 106068 77824
rect 106004 77764 106008 77820
rect 106008 77764 106064 77820
rect 106064 77764 106068 77820
rect 106004 77760 106068 77764
rect 106084 77820 106148 77824
rect 106084 77764 106088 77820
rect 106088 77764 106144 77820
rect 106144 77764 106148 77820
rect 106084 77760 106148 77764
rect 106164 77820 106228 77824
rect 106164 77764 106168 77820
rect 106168 77764 106224 77820
rect 106224 77764 106228 77820
rect 106164 77760 106228 77764
rect 4876 77276 4940 77280
rect 4876 77220 4880 77276
rect 4880 77220 4936 77276
rect 4936 77220 4940 77276
rect 4876 77216 4940 77220
rect 4956 77276 5020 77280
rect 4956 77220 4960 77276
rect 4960 77220 5016 77276
rect 5016 77220 5020 77276
rect 4956 77216 5020 77220
rect 5036 77276 5100 77280
rect 5036 77220 5040 77276
rect 5040 77220 5096 77276
rect 5096 77220 5100 77276
rect 5036 77216 5100 77220
rect 5116 77276 5180 77280
rect 5116 77220 5120 77276
rect 5120 77220 5176 77276
rect 5176 77220 5180 77276
rect 5116 77216 5180 77220
rect 106660 77276 106724 77280
rect 106660 77220 106664 77276
rect 106664 77220 106720 77276
rect 106720 77220 106724 77276
rect 106660 77216 106724 77220
rect 106740 77276 106804 77280
rect 106740 77220 106744 77276
rect 106744 77220 106800 77276
rect 106800 77220 106804 77276
rect 106740 77216 106804 77220
rect 106820 77276 106884 77280
rect 106820 77220 106824 77276
rect 106824 77220 106880 77276
rect 106880 77220 106884 77276
rect 106820 77216 106884 77220
rect 106900 77276 106964 77280
rect 106900 77220 106904 77276
rect 106904 77220 106960 77276
rect 106960 77220 106964 77276
rect 106900 77216 106964 77220
rect 4216 76732 4280 76736
rect 4216 76676 4220 76732
rect 4220 76676 4276 76732
rect 4276 76676 4280 76732
rect 4216 76672 4280 76676
rect 4296 76732 4360 76736
rect 4296 76676 4300 76732
rect 4300 76676 4356 76732
rect 4356 76676 4360 76732
rect 4296 76672 4360 76676
rect 4376 76732 4440 76736
rect 4376 76676 4380 76732
rect 4380 76676 4436 76732
rect 4436 76676 4440 76732
rect 4376 76672 4440 76676
rect 4456 76732 4520 76736
rect 4456 76676 4460 76732
rect 4460 76676 4516 76732
rect 4516 76676 4520 76732
rect 4456 76672 4520 76676
rect 105924 76732 105988 76736
rect 105924 76676 105928 76732
rect 105928 76676 105984 76732
rect 105984 76676 105988 76732
rect 105924 76672 105988 76676
rect 106004 76732 106068 76736
rect 106004 76676 106008 76732
rect 106008 76676 106064 76732
rect 106064 76676 106068 76732
rect 106004 76672 106068 76676
rect 106084 76732 106148 76736
rect 106084 76676 106088 76732
rect 106088 76676 106144 76732
rect 106144 76676 106148 76732
rect 106084 76672 106148 76676
rect 106164 76732 106228 76736
rect 106164 76676 106168 76732
rect 106168 76676 106224 76732
rect 106224 76676 106228 76732
rect 106164 76672 106228 76676
rect 4876 76188 4940 76192
rect 4876 76132 4880 76188
rect 4880 76132 4936 76188
rect 4936 76132 4940 76188
rect 4876 76128 4940 76132
rect 4956 76188 5020 76192
rect 4956 76132 4960 76188
rect 4960 76132 5016 76188
rect 5016 76132 5020 76188
rect 4956 76128 5020 76132
rect 5036 76188 5100 76192
rect 5036 76132 5040 76188
rect 5040 76132 5096 76188
rect 5096 76132 5100 76188
rect 5036 76128 5100 76132
rect 5116 76188 5180 76192
rect 5116 76132 5120 76188
rect 5120 76132 5176 76188
rect 5176 76132 5180 76188
rect 5116 76128 5180 76132
rect 106660 76188 106724 76192
rect 106660 76132 106664 76188
rect 106664 76132 106720 76188
rect 106720 76132 106724 76188
rect 106660 76128 106724 76132
rect 106740 76188 106804 76192
rect 106740 76132 106744 76188
rect 106744 76132 106800 76188
rect 106800 76132 106804 76188
rect 106740 76128 106804 76132
rect 106820 76188 106884 76192
rect 106820 76132 106824 76188
rect 106824 76132 106880 76188
rect 106880 76132 106884 76188
rect 106820 76128 106884 76132
rect 106900 76188 106964 76192
rect 106900 76132 106904 76188
rect 106904 76132 106960 76188
rect 106960 76132 106964 76188
rect 106900 76128 106964 76132
rect 4216 75644 4280 75648
rect 4216 75588 4220 75644
rect 4220 75588 4276 75644
rect 4276 75588 4280 75644
rect 4216 75584 4280 75588
rect 4296 75644 4360 75648
rect 4296 75588 4300 75644
rect 4300 75588 4356 75644
rect 4356 75588 4360 75644
rect 4296 75584 4360 75588
rect 4376 75644 4440 75648
rect 4376 75588 4380 75644
rect 4380 75588 4436 75644
rect 4436 75588 4440 75644
rect 4376 75584 4440 75588
rect 4456 75644 4520 75648
rect 4456 75588 4460 75644
rect 4460 75588 4516 75644
rect 4516 75588 4520 75644
rect 4456 75584 4520 75588
rect 105924 75644 105988 75648
rect 105924 75588 105928 75644
rect 105928 75588 105984 75644
rect 105984 75588 105988 75644
rect 105924 75584 105988 75588
rect 106004 75644 106068 75648
rect 106004 75588 106008 75644
rect 106008 75588 106064 75644
rect 106064 75588 106068 75644
rect 106004 75584 106068 75588
rect 106084 75644 106148 75648
rect 106084 75588 106088 75644
rect 106088 75588 106144 75644
rect 106144 75588 106148 75644
rect 106084 75584 106148 75588
rect 106164 75644 106228 75648
rect 106164 75588 106168 75644
rect 106168 75588 106224 75644
rect 106224 75588 106228 75644
rect 106164 75584 106228 75588
rect 4876 75100 4940 75104
rect 4876 75044 4880 75100
rect 4880 75044 4936 75100
rect 4936 75044 4940 75100
rect 4876 75040 4940 75044
rect 4956 75100 5020 75104
rect 4956 75044 4960 75100
rect 4960 75044 5016 75100
rect 5016 75044 5020 75100
rect 4956 75040 5020 75044
rect 5036 75100 5100 75104
rect 5036 75044 5040 75100
rect 5040 75044 5096 75100
rect 5096 75044 5100 75100
rect 5036 75040 5100 75044
rect 5116 75100 5180 75104
rect 5116 75044 5120 75100
rect 5120 75044 5176 75100
rect 5176 75044 5180 75100
rect 5116 75040 5180 75044
rect 106660 75100 106724 75104
rect 106660 75044 106664 75100
rect 106664 75044 106720 75100
rect 106720 75044 106724 75100
rect 106660 75040 106724 75044
rect 106740 75100 106804 75104
rect 106740 75044 106744 75100
rect 106744 75044 106800 75100
rect 106800 75044 106804 75100
rect 106740 75040 106804 75044
rect 106820 75100 106884 75104
rect 106820 75044 106824 75100
rect 106824 75044 106880 75100
rect 106880 75044 106884 75100
rect 106820 75040 106884 75044
rect 106900 75100 106964 75104
rect 106900 75044 106904 75100
rect 106904 75044 106960 75100
rect 106960 75044 106964 75100
rect 106900 75040 106964 75044
rect 4216 74556 4280 74560
rect 4216 74500 4220 74556
rect 4220 74500 4276 74556
rect 4276 74500 4280 74556
rect 4216 74496 4280 74500
rect 4296 74556 4360 74560
rect 4296 74500 4300 74556
rect 4300 74500 4356 74556
rect 4356 74500 4360 74556
rect 4296 74496 4360 74500
rect 4376 74556 4440 74560
rect 4376 74500 4380 74556
rect 4380 74500 4436 74556
rect 4436 74500 4440 74556
rect 4376 74496 4440 74500
rect 4456 74556 4520 74560
rect 4456 74500 4460 74556
rect 4460 74500 4516 74556
rect 4516 74500 4520 74556
rect 4456 74496 4520 74500
rect 105924 74556 105988 74560
rect 105924 74500 105928 74556
rect 105928 74500 105984 74556
rect 105984 74500 105988 74556
rect 105924 74496 105988 74500
rect 106004 74556 106068 74560
rect 106004 74500 106008 74556
rect 106008 74500 106064 74556
rect 106064 74500 106068 74556
rect 106004 74496 106068 74500
rect 106084 74556 106148 74560
rect 106084 74500 106088 74556
rect 106088 74500 106144 74556
rect 106144 74500 106148 74556
rect 106084 74496 106148 74500
rect 106164 74556 106228 74560
rect 106164 74500 106168 74556
rect 106168 74500 106224 74556
rect 106224 74500 106228 74556
rect 106164 74496 106228 74500
rect 4876 74012 4940 74016
rect 4876 73956 4880 74012
rect 4880 73956 4936 74012
rect 4936 73956 4940 74012
rect 4876 73952 4940 73956
rect 4956 74012 5020 74016
rect 4956 73956 4960 74012
rect 4960 73956 5016 74012
rect 5016 73956 5020 74012
rect 4956 73952 5020 73956
rect 5036 74012 5100 74016
rect 5036 73956 5040 74012
rect 5040 73956 5096 74012
rect 5096 73956 5100 74012
rect 5036 73952 5100 73956
rect 5116 74012 5180 74016
rect 5116 73956 5120 74012
rect 5120 73956 5176 74012
rect 5176 73956 5180 74012
rect 5116 73952 5180 73956
rect 106660 74012 106724 74016
rect 106660 73956 106664 74012
rect 106664 73956 106720 74012
rect 106720 73956 106724 74012
rect 106660 73952 106724 73956
rect 106740 74012 106804 74016
rect 106740 73956 106744 74012
rect 106744 73956 106800 74012
rect 106800 73956 106804 74012
rect 106740 73952 106804 73956
rect 106820 74012 106884 74016
rect 106820 73956 106824 74012
rect 106824 73956 106880 74012
rect 106880 73956 106884 74012
rect 106820 73952 106884 73956
rect 106900 74012 106964 74016
rect 106900 73956 106904 74012
rect 106904 73956 106960 74012
rect 106960 73956 106964 74012
rect 106900 73952 106964 73956
rect 4216 73468 4280 73472
rect 4216 73412 4220 73468
rect 4220 73412 4276 73468
rect 4276 73412 4280 73468
rect 4216 73408 4280 73412
rect 4296 73468 4360 73472
rect 4296 73412 4300 73468
rect 4300 73412 4356 73468
rect 4356 73412 4360 73468
rect 4296 73408 4360 73412
rect 4376 73468 4440 73472
rect 4376 73412 4380 73468
rect 4380 73412 4436 73468
rect 4436 73412 4440 73468
rect 4376 73408 4440 73412
rect 4456 73468 4520 73472
rect 4456 73412 4460 73468
rect 4460 73412 4516 73468
rect 4516 73412 4520 73468
rect 4456 73408 4520 73412
rect 105924 73468 105988 73472
rect 105924 73412 105928 73468
rect 105928 73412 105984 73468
rect 105984 73412 105988 73468
rect 105924 73408 105988 73412
rect 106004 73468 106068 73472
rect 106004 73412 106008 73468
rect 106008 73412 106064 73468
rect 106064 73412 106068 73468
rect 106004 73408 106068 73412
rect 106084 73468 106148 73472
rect 106084 73412 106088 73468
rect 106088 73412 106144 73468
rect 106144 73412 106148 73468
rect 106084 73408 106148 73412
rect 106164 73468 106228 73472
rect 106164 73412 106168 73468
rect 106168 73412 106224 73468
rect 106224 73412 106228 73468
rect 106164 73408 106228 73412
rect 4876 72924 4940 72928
rect 4876 72868 4880 72924
rect 4880 72868 4936 72924
rect 4936 72868 4940 72924
rect 4876 72864 4940 72868
rect 4956 72924 5020 72928
rect 4956 72868 4960 72924
rect 4960 72868 5016 72924
rect 5016 72868 5020 72924
rect 4956 72864 5020 72868
rect 5036 72924 5100 72928
rect 5036 72868 5040 72924
rect 5040 72868 5096 72924
rect 5096 72868 5100 72924
rect 5036 72864 5100 72868
rect 5116 72924 5180 72928
rect 5116 72868 5120 72924
rect 5120 72868 5176 72924
rect 5176 72868 5180 72924
rect 5116 72864 5180 72868
rect 106660 72924 106724 72928
rect 106660 72868 106664 72924
rect 106664 72868 106720 72924
rect 106720 72868 106724 72924
rect 106660 72864 106724 72868
rect 106740 72924 106804 72928
rect 106740 72868 106744 72924
rect 106744 72868 106800 72924
rect 106800 72868 106804 72924
rect 106740 72864 106804 72868
rect 106820 72924 106884 72928
rect 106820 72868 106824 72924
rect 106824 72868 106880 72924
rect 106880 72868 106884 72924
rect 106820 72864 106884 72868
rect 106900 72924 106964 72928
rect 106900 72868 106904 72924
rect 106904 72868 106960 72924
rect 106960 72868 106964 72924
rect 106900 72864 106964 72868
rect 4216 72380 4280 72384
rect 4216 72324 4220 72380
rect 4220 72324 4276 72380
rect 4276 72324 4280 72380
rect 4216 72320 4280 72324
rect 4296 72380 4360 72384
rect 4296 72324 4300 72380
rect 4300 72324 4356 72380
rect 4356 72324 4360 72380
rect 4296 72320 4360 72324
rect 4376 72380 4440 72384
rect 4376 72324 4380 72380
rect 4380 72324 4436 72380
rect 4436 72324 4440 72380
rect 4376 72320 4440 72324
rect 4456 72380 4520 72384
rect 4456 72324 4460 72380
rect 4460 72324 4516 72380
rect 4516 72324 4520 72380
rect 4456 72320 4520 72324
rect 105924 72380 105988 72384
rect 105924 72324 105928 72380
rect 105928 72324 105984 72380
rect 105984 72324 105988 72380
rect 105924 72320 105988 72324
rect 106004 72380 106068 72384
rect 106004 72324 106008 72380
rect 106008 72324 106064 72380
rect 106064 72324 106068 72380
rect 106004 72320 106068 72324
rect 106084 72380 106148 72384
rect 106084 72324 106088 72380
rect 106088 72324 106144 72380
rect 106144 72324 106148 72380
rect 106084 72320 106148 72324
rect 106164 72380 106228 72384
rect 106164 72324 106168 72380
rect 106168 72324 106224 72380
rect 106224 72324 106228 72380
rect 106164 72320 106228 72324
rect 4876 71836 4940 71840
rect 4876 71780 4880 71836
rect 4880 71780 4936 71836
rect 4936 71780 4940 71836
rect 4876 71776 4940 71780
rect 4956 71836 5020 71840
rect 4956 71780 4960 71836
rect 4960 71780 5016 71836
rect 5016 71780 5020 71836
rect 4956 71776 5020 71780
rect 5036 71836 5100 71840
rect 5036 71780 5040 71836
rect 5040 71780 5096 71836
rect 5096 71780 5100 71836
rect 5036 71776 5100 71780
rect 5116 71836 5180 71840
rect 5116 71780 5120 71836
rect 5120 71780 5176 71836
rect 5176 71780 5180 71836
rect 5116 71776 5180 71780
rect 106660 71836 106724 71840
rect 106660 71780 106664 71836
rect 106664 71780 106720 71836
rect 106720 71780 106724 71836
rect 106660 71776 106724 71780
rect 106740 71836 106804 71840
rect 106740 71780 106744 71836
rect 106744 71780 106800 71836
rect 106800 71780 106804 71836
rect 106740 71776 106804 71780
rect 106820 71836 106884 71840
rect 106820 71780 106824 71836
rect 106824 71780 106880 71836
rect 106880 71780 106884 71836
rect 106820 71776 106884 71780
rect 106900 71836 106964 71840
rect 106900 71780 106904 71836
rect 106904 71780 106960 71836
rect 106960 71780 106964 71836
rect 106900 71776 106964 71780
rect 4216 71292 4280 71296
rect 4216 71236 4220 71292
rect 4220 71236 4276 71292
rect 4276 71236 4280 71292
rect 4216 71232 4280 71236
rect 4296 71292 4360 71296
rect 4296 71236 4300 71292
rect 4300 71236 4356 71292
rect 4356 71236 4360 71292
rect 4296 71232 4360 71236
rect 4376 71292 4440 71296
rect 4376 71236 4380 71292
rect 4380 71236 4436 71292
rect 4436 71236 4440 71292
rect 4376 71232 4440 71236
rect 4456 71292 4520 71296
rect 4456 71236 4460 71292
rect 4460 71236 4516 71292
rect 4516 71236 4520 71292
rect 4456 71232 4520 71236
rect 105924 71292 105988 71296
rect 105924 71236 105928 71292
rect 105928 71236 105984 71292
rect 105984 71236 105988 71292
rect 105924 71232 105988 71236
rect 106004 71292 106068 71296
rect 106004 71236 106008 71292
rect 106008 71236 106064 71292
rect 106064 71236 106068 71292
rect 106004 71232 106068 71236
rect 106084 71292 106148 71296
rect 106084 71236 106088 71292
rect 106088 71236 106144 71292
rect 106144 71236 106148 71292
rect 106084 71232 106148 71236
rect 106164 71292 106228 71296
rect 106164 71236 106168 71292
rect 106168 71236 106224 71292
rect 106224 71236 106228 71292
rect 106164 71232 106228 71236
rect 4876 70748 4940 70752
rect 4876 70692 4880 70748
rect 4880 70692 4936 70748
rect 4936 70692 4940 70748
rect 4876 70688 4940 70692
rect 4956 70748 5020 70752
rect 4956 70692 4960 70748
rect 4960 70692 5016 70748
rect 5016 70692 5020 70748
rect 4956 70688 5020 70692
rect 5036 70748 5100 70752
rect 5036 70692 5040 70748
rect 5040 70692 5096 70748
rect 5096 70692 5100 70748
rect 5036 70688 5100 70692
rect 5116 70748 5180 70752
rect 5116 70692 5120 70748
rect 5120 70692 5176 70748
rect 5176 70692 5180 70748
rect 5116 70688 5180 70692
rect 106660 70748 106724 70752
rect 106660 70692 106664 70748
rect 106664 70692 106720 70748
rect 106720 70692 106724 70748
rect 106660 70688 106724 70692
rect 106740 70748 106804 70752
rect 106740 70692 106744 70748
rect 106744 70692 106800 70748
rect 106800 70692 106804 70748
rect 106740 70688 106804 70692
rect 106820 70748 106884 70752
rect 106820 70692 106824 70748
rect 106824 70692 106880 70748
rect 106880 70692 106884 70748
rect 106820 70688 106884 70692
rect 106900 70748 106964 70752
rect 106900 70692 106904 70748
rect 106904 70692 106960 70748
rect 106960 70692 106964 70748
rect 106900 70688 106964 70692
rect 4216 70204 4280 70208
rect 4216 70148 4220 70204
rect 4220 70148 4276 70204
rect 4276 70148 4280 70204
rect 4216 70144 4280 70148
rect 4296 70204 4360 70208
rect 4296 70148 4300 70204
rect 4300 70148 4356 70204
rect 4356 70148 4360 70204
rect 4296 70144 4360 70148
rect 4376 70204 4440 70208
rect 4376 70148 4380 70204
rect 4380 70148 4436 70204
rect 4436 70148 4440 70204
rect 4376 70144 4440 70148
rect 4456 70204 4520 70208
rect 4456 70148 4460 70204
rect 4460 70148 4516 70204
rect 4516 70148 4520 70204
rect 4456 70144 4520 70148
rect 105924 70204 105988 70208
rect 105924 70148 105928 70204
rect 105928 70148 105984 70204
rect 105984 70148 105988 70204
rect 105924 70144 105988 70148
rect 106004 70204 106068 70208
rect 106004 70148 106008 70204
rect 106008 70148 106064 70204
rect 106064 70148 106068 70204
rect 106004 70144 106068 70148
rect 106084 70204 106148 70208
rect 106084 70148 106088 70204
rect 106088 70148 106144 70204
rect 106144 70148 106148 70204
rect 106084 70144 106148 70148
rect 106164 70204 106228 70208
rect 106164 70148 106168 70204
rect 106168 70148 106224 70204
rect 106224 70148 106228 70204
rect 106164 70144 106228 70148
rect 33950 69804 34014 69868
rect 37454 69864 37518 69868
rect 37454 69808 37462 69864
rect 37462 69808 37518 69864
rect 37454 69804 37518 69808
rect 38622 69864 38686 69868
rect 38622 69808 38658 69864
rect 38658 69808 38686 69864
rect 38622 69804 38686 69808
rect 39790 69864 39854 69868
rect 39790 69808 39818 69864
rect 39818 69808 39854 69864
rect 39790 69804 39854 69808
rect 40958 69864 41022 69868
rect 40958 69808 41014 69864
rect 41014 69808 41022 69864
rect 40958 69804 41022 69808
rect 43294 69864 43358 69868
rect 43294 69808 43314 69864
rect 43314 69808 43358 69864
rect 43294 69804 43358 69808
rect 90680 69804 90744 69868
rect 4876 69660 4940 69664
rect 4876 69604 4880 69660
rect 4880 69604 4936 69660
rect 4936 69604 4940 69660
rect 4876 69600 4940 69604
rect 4956 69660 5020 69664
rect 4956 69604 4960 69660
rect 4960 69604 5016 69660
rect 5016 69604 5020 69660
rect 4956 69600 5020 69604
rect 5036 69660 5100 69664
rect 5036 69604 5040 69660
rect 5040 69604 5096 69660
rect 5096 69604 5100 69660
rect 5036 69600 5100 69604
rect 5116 69660 5180 69664
rect 5116 69604 5120 69660
rect 5120 69604 5176 69660
rect 5176 69604 5180 69660
rect 5116 69600 5180 69604
rect 23438 69592 23502 69596
rect 23438 69536 23478 69592
rect 23478 69536 23502 69592
rect 23438 69532 23502 69536
rect 24624 69592 24688 69596
rect 24624 69536 24674 69592
rect 24674 69536 24688 69592
rect 24624 69532 24688 69536
rect 25774 69592 25838 69596
rect 25774 69536 25778 69592
rect 25778 69536 25834 69592
rect 25834 69536 25838 69592
rect 25774 69532 25838 69536
rect 26942 69592 27006 69596
rect 26942 69536 26974 69592
rect 26974 69536 27006 69592
rect 26942 69532 27006 69536
rect 28110 69592 28174 69596
rect 28110 69536 28134 69592
rect 28134 69536 28174 69592
rect 28110 69532 28174 69536
rect 30446 69592 30510 69596
rect 30446 69536 30470 69592
rect 30470 69536 30510 69592
rect 30446 69532 30510 69536
rect 106660 69660 106724 69664
rect 106660 69604 106664 69660
rect 106664 69604 106720 69660
rect 106720 69604 106724 69660
rect 106660 69600 106724 69604
rect 106740 69660 106804 69664
rect 106740 69604 106744 69660
rect 106744 69604 106800 69660
rect 106800 69604 106804 69660
rect 106740 69600 106804 69604
rect 106820 69660 106884 69664
rect 106820 69604 106824 69660
rect 106824 69604 106880 69660
rect 106880 69604 106884 69660
rect 106820 69600 106884 69604
rect 106900 69660 106964 69664
rect 106900 69604 106904 69660
rect 106904 69604 106960 69660
rect 106960 69604 106964 69660
rect 106900 69600 106964 69604
rect 31614 69532 31678 69596
rect 32812 69592 32876 69596
rect 32812 69536 32862 69592
rect 32862 69536 32876 69592
rect 32812 69532 32876 69536
rect 33950 69592 34014 69596
rect 33950 69536 33966 69592
rect 33966 69536 34014 69592
rect 33950 69532 34014 69536
rect 35118 69592 35182 69596
rect 35118 69536 35162 69592
rect 35162 69536 35182 69592
rect 35118 69532 35182 69536
rect 36308 69592 36372 69596
rect 36308 69536 36358 69592
rect 36358 69536 36372 69592
rect 36308 69532 36372 69536
rect 42126 69592 42190 69596
rect 42126 69536 42154 69592
rect 42154 69536 42190 69592
rect 42126 69532 42190 69536
rect 90527 69532 90591 69596
rect 29316 69260 29380 69324
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 105924 69116 105988 69120
rect 105924 69060 105928 69116
rect 105928 69060 105984 69116
rect 105984 69060 105988 69116
rect 105924 69056 105988 69060
rect 106004 69116 106068 69120
rect 106004 69060 106008 69116
rect 106008 69060 106064 69116
rect 106064 69060 106068 69116
rect 106004 69056 106068 69060
rect 106084 69116 106148 69120
rect 106084 69060 106088 69116
rect 106088 69060 106144 69116
rect 106144 69060 106148 69116
rect 106084 69056 106148 69060
rect 106164 69116 106228 69120
rect 106164 69060 106168 69116
rect 106168 69060 106224 69116
rect 106224 69060 106228 69116
rect 106164 69056 106228 69060
rect 90772 68776 90836 68780
rect 90772 68720 90822 68776
rect 90822 68720 90836 68776
rect 90772 68716 90836 68720
rect 4876 68572 4940 68576
rect 4876 68516 4880 68572
rect 4880 68516 4936 68572
rect 4936 68516 4940 68572
rect 4876 68512 4940 68516
rect 4956 68572 5020 68576
rect 4956 68516 4960 68572
rect 4960 68516 5016 68572
rect 5016 68516 5020 68572
rect 4956 68512 5020 68516
rect 5036 68572 5100 68576
rect 5036 68516 5040 68572
rect 5040 68516 5096 68572
rect 5096 68516 5100 68572
rect 5036 68512 5100 68516
rect 5116 68572 5180 68576
rect 5116 68516 5120 68572
rect 5120 68516 5176 68572
rect 5176 68516 5180 68572
rect 5116 68512 5180 68516
rect 106660 68572 106724 68576
rect 106660 68516 106664 68572
rect 106664 68516 106720 68572
rect 106720 68516 106724 68572
rect 106660 68512 106724 68516
rect 106740 68572 106804 68576
rect 106740 68516 106744 68572
rect 106744 68516 106800 68572
rect 106800 68516 106804 68572
rect 106740 68512 106804 68516
rect 106820 68572 106884 68576
rect 106820 68516 106824 68572
rect 106824 68516 106880 68572
rect 106880 68516 106884 68572
rect 106820 68512 106884 68516
rect 106900 68572 106964 68576
rect 106900 68516 106904 68572
rect 106904 68516 106960 68572
rect 106960 68516 106964 68572
rect 106900 68512 106964 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 65656 68028 65720 68032
rect 65656 67972 65660 68028
rect 65660 67972 65716 68028
rect 65716 67972 65720 68028
rect 65656 67968 65720 67972
rect 65736 68028 65800 68032
rect 65736 67972 65740 68028
rect 65740 67972 65796 68028
rect 65796 67972 65800 68028
rect 65736 67968 65800 67972
rect 65816 68028 65880 68032
rect 65816 67972 65820 68028
rect 65820 67972 65876 68028
rect 65876 67972 65880 68028
rect 65816 67968 65880 67972
rect 65896 68028 65960 68032
rect 65896 67972 65900 68028
rect 65900 67972 65956 68028
rect 65956 67972 65960 68028
rect 65896 67968 65960 67972
rect 96376 68028 96440 68032
rect 96376 67972 96380 68028
rect 96380 67972 96436 68028
rect 96436 67972 96440 68028
rect 96376 67968 96440 67972
rect 96456 68028 96520 68032
rect 96456 67972 96460 68028
rect 96460 67972 96516 68028
rect 96516 67972 96520 68028
rect 96456 67968 96520 67972
rect 96536 68028 96600 68032
rect 96536 67972 96540 68028
rect 96540 67972 96596 68028
rect 96596 67972 96600 68028
rect 96536 67968 96600 67972
rect 96616 68028 96680 68032
rect 96616 67972 96620 68028
rect 96620 67972 96676 68028
rect 96676 67972 96680 68028
rect 96616 67968 96680 67972
rect 105924 68028 105988 68032
rect 105924 67972 105928 68028
rect 105928 67972 105984 68028
rect 105984 67972 105988 68028
rect 105924 67968 105988 67972
rect 106004 68028 106068 68032
rect 106004 67972 106008 68028
rect 106008 67972 106064 68028
rect 106064 67972 106068 68028
rect 106004 67968 106068 67972
rect 106084 68028 106148 68032
rect 106084 67972 106088 68028
rect 106088 67972 106144 68028
rect 106144 67972 106148 68028
rect 106084 67968 106148 67972
rect 106164 68028 106228 68032
rect 106164 67972 106168 68028
rect 106168 67972 106224 68028
rect 106224 67972 106228 68028
rect 106164 67968 106228 67972
rect 16068 67628 16132 67692
rect 86172 67628 86236 67692
rect 4876 67484 4940 67488
rect 4876 67428 4880 67484
rect 4880 67428 4936 67484
rect 4936 67428 4940 67484
rect 4876 67424 4940 67428
rect 4956 67484 5020 67488
rect 4956 67428 4960 67484
rect 4960 67428 5016 67484
rect 5016 67428 5020 67484
rect 4956 67424 5020 67428
rect 5036 67484 5100 67488
rect 5036 67428 5040 67484
rect 5040 67428 5096 67484
rect 5096 67428 5100 67484
rect 5036 67424 5100 67428
rect 5116 67484 5180 67488
rect 5116 67428 5120 67484
rect 5120 67428 5176 67484
rect 5176 67428 5180 67484
rect 5116 67424 5180 67428
rect 35596 67484 35660 67488
rect 35596 67428 35600 67484
rect 35600 67428 35656 67484
rect 35656 67428 35660 67484
rect 35596 67424 35660 67428
rect 35676 67484 35740 67488
rect 35676 67428 35680 67484
rect 35680 67428 35736 67484
rect 35736 67428 35740 67484
rect 35676 67424 35740 67428
rect 35756 67484 35820 67488
rect 35756 67428 35760 67484
rect 35760 67428 35816 67484
rect 35816 67428 35820 67484
rect 35756 67424 35820 67428
rect 35836 67484 35900 67488
rect 35836 67428 35840 67484
rect 35840 67428 35896 67484
rect 35896 67428 35900 67484
rect 35836 67424 35900 67428
rect 66316 67484 66380 67488
rect 66316 67428 66320 67484
rect 66320 67428 66376 67484
rect 66376 67428 66380 67484
rect 66316 67424 66380 67428
rect 66396 67484 66460 67488
rect 66396 67428 66400 67484
rect 66400 67428 66456 67484
rect 66456 67428 66460 67484
rect 66396 67424 66460 67428
rect 66476 67484 66540 67488
rect 66476 67428 66480 67484
rect 66480 67428 66536 67484
rect 66536 67428 66540 67484
rect 66476 67424 66540 67428
rect 66556 67484 66620 67488
rect 66556 67428 66560 67484
rect 66560 67428 66616 67484
rect 66616 67428 66620 67484
rect 66556 67424 66620 67428
rect 97036 67484 97100 67488
rect 97036 67428 97040 67484
rect 97040 67428 97096 67484
rect 97096 67428 97100 67484
rect 97036 67424 97100 67428
rect 97116 67484 97180 67488
rect 97116 67428 97120 67484
rect 97120 67428 97176 67484
rect 97176 67428 97180 67484
rect 97116 67424 97180 67428
rect 97196 67484 97260 67488
rect 97196 67428 97200 67484
rect 97200 67428 97256 67484
rect 97256 67428 97260 67484
rect 97196 67424 97260 67428
rect 97276 67484 97340 67488
rect 97276 67428 97280 67484
rect 97280 67428 97336 67484
rect 97336 67428 97340 67484
rect 97276 67424 97340 67428
rect 106660 67484 106724 67488
rect 106660 67428 106664 67484
rect 106664 67428 106720 67484
rect 106720 67428 106724 67484
rect 106660 67424 106724 67428
rect 106740 67484 106804 67488
rect 106740 67428 106744 67484
rect 106744 67428 106800 67484
rect 106800 67428 106804 67484
rect 106740 67424 106804 67428
rect 106820 67484 106884 67488
rect 106820 67428 106824 67484
rect 106824 67428 106880 67484
rect 106880 67428 106884 67484
rect 106820 67424 106884 67428
rect 106900 67484 106964 67488
rect 106900 67428 106904 67484
rect 106904 67428 106960 67484
rect 106960 67428 106964 67484
rect 106900 67424 106964 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 96376 66940 96440 66944
rect 96376 66884 96380 66940
rect 96380 66884 96436 66940
rect 96436 66884 96440 66940
rect 96376 66880 96440 66884
rect 96456 66940 96520 66944
rect 96456 66884 96460 66940
rect 96460 66884 96516 66940
rect 96516 66884 96520 66940
rect 96456 66880 96520 66884
rect 96536 66940 96600 66944
rect 96536 66884 96540 66940
rect 96540 66884 96596 66940
rect 96596 66884 96600 66940
rect 96536 66880 96600 66884
rect 96616 66940 96680 66944
rect 96616 66884 96620 66940
rect 96620 66884 96676 66940
rect 96676 66884 96680 66940
rect 96616 66880 96680 66884
rect 63540 66676 63604 66740
rect 36124 66540 36188 66604
rect 51028 66540 51092 66604
rect 66116 66540 66180 66604
rect 4876 66396 4940 66400
rect 4876 66340 4880 66396
rect 4880 66340 4936 66396
rect 4936 66340 4940 66396
rect 4876 66336 4940 66340
rect 4956 66396 5020 66400
rect 4956 66340 4960 66396
rect 4960 66340 5016 66396
rect 5016 66340 5020 66396
rect 4956 66336 5020 66340
rect 5036 66396 5100 66400
rect 5036 66340 5040 66396
rect 5040 66340 5096 66396
rect 5096 66340 5100 66396
rect 5036 66336 5100 66340
rect 5116 66396 5180 66400
rect 5116 66340 5120 66396
rect 5120 66340 5176 66396
rect 5176 66340 5180 66396
rect 5116 66336 5180 66340
rect 35596 66396 35660 66400
rect 35596 66340 35600 66396
rect 35600 66340 35656 66396
rect 35656 66340 35660 66396
rect 35596 66336 35660 66340
rect 35676 66396 35740 66400
rect 35676 66340 35680 66396
rect 35680 66340 35736 66396
rect 35736 66340 35740 66396
rect 35676 66336 35740 66340
rect 35756 66396 35820 66400
rect 35756 66340 35760 66396
rect 35760 66340 35816 66396
rect 35816 66340 35820 66396
rect 35756 66336 35820 66340
rect 35836 66396 35900 66400
rect 35836 66340 35840 66396
rect 35840 66340 35896 66396
rect 35896 66340 35900 66396
rect 35836 66336 35900 66340
rect 66316 66396 66380 66400
rect 66316 66340 66320 66396
rect 66320 66340 66376 66396
rect 66376 66340 66380 66396
rect 66316 66336 66380 66340
rect 66396 66396 66460 66400
rect 66396 66340 66400 66396
rect 66400 66340 66456 66396
rect 66456 66340 66460 66396
rect 66396 66336 66460 66340
rect 66476 66396 66540 66400
rect 66476 66340 66480 66396
rect 66480 66340 66536 66396
rect 66536 66340 66540 66396
rect 66476 66336 66540 66340
rect 66556 66396 66620 66400
rect 66556 66340 66560 66396
rect 66560 66340 66616 66396
rect 66616 66340 66620 66396
rect 66556 66336 66620 66340
rect 97036 66396 97100 66400
rect 97036 66340 97040 66396
rect 97040 66340 97096 66396
rect 97096 66340 97100 66396
rect 97036 66336 97100 66340
rect 97116 66396 97180 66400
rect 97116 66340 97120 66396
rect 97120 66340 97176 66396
rect 97176 66340 97180 66396
rect 97116 66336 97180 66340
rect 97196 66396 97260 66400
rect 97196 66340 97200 66396
rect 97200 66340 97256 66396
rect 97256 66340 97260 66396
rect 97196 66336 97260 66340
rect 97276 66396 97340 66400
rect 97276 66340 97280 66396
rect 97280 66340 97336 66396
rect 97336 66340 97340 66396
rect 97276 66336 97340 66340
rect 106660 66396 106724 66400
rect 106660 66340 106664 66396
rect 106664 66340 106720 66396
rect 106720 66340 106724 66396
rect 106660 66336 106724 66340
rect 106740 66396 106804 66400
rect 106740 66340 106744 66396
rect 106744 66340 106800 66396
rect 106800 66340 106804 66396
rect 106740 66336 106804 66340
rect 106820 66396 106884 66400
rect 106820 66340 106824 66396
rect 106824 66340 106880 66396
rect 106880 66340 106884 66396
rect 106820 66336 106884 66340
rect 106900 66396 106964 66400
rect 106900 66340 106904 66396
rect 106904 66340 106960 66396
rect 106960 66340 106964 66396
rect 106900 66336 106964 66340
rect 41092 66268 41156 66332
rect 71084 66268 71148 66332
rect 87276 66268 87340 66332
rect 46060 66132 46124 66196
rect 53604 65920 53668 65924
rect 53604 65864 53654 65920
rect 53654 65864 53668 65920
rect 53604 65860 53668 65864
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 96376 65852 96440 65856
rect 96376 65796 96380 65852
rect 96380 65796 96436 65852
rect 96436 65796 96440 65852
rect 96376 65792 96440 65796
rect 96456 65852 96520 65856
rect 96456 65796 96460 65852
rect 96460 65796 96516 65852
rect 96516 65796 96520 65852
rect 96456 65792 96520 65796
rect 96536 65852 96600 65856
rect 96536 65796 96540 65852
rect 96540 65796 96596 65852
rect 96596 65796 96600 65852
rect 96536 65792 96600 65796
rect 96616 65852 96680 65856
rect 96616 65796 96620 65852
rect 96620 65796 96676 65852
rect 96676 65796 96680 65852
rect 96616 65792 96680 65796
rect 105924 65852 105988 65856
rect 105924 65796 105928 65852
rect 105928 65796 105984 65852
rect 105984 65796 105988 65852
rect 105924 65792 105988 65796
rect 106004 65852 106068 65856
rect 106004 65796 106008 65852
rect 106008 65796 106064 65852
rect 106064 65796 106068 65852
rect 106004 65792 106068 65796
rect 106084 65852 106148 65856
rect 106084 65796 106088 65852
rect 106088 65796 106144 65852
rect 106144 65796 106148 65852
rect 106084 65792 106148 65796
rect 106164 65852 106228 65856
rect 106164 65796 106168 65852
rect 106168 65796 106224 65852
rect 106224 65796 106228 65852
rect 106164 65792 106228 65796
rect 43484 65452 43548 65516
rect 73476 65452 73540 65516
rect 4876 65308 4940 65312
rect 4876 65252 4880 65308
rect 4880 65252 4936 65308
rect 4936 65252 4940 65308
rect 4876 65248 4940 65252
rect 4956 65308 5020 65312
rect 4956 65252 4960 65308
rect 4960 65252 5016 65308
rect 5016 65252 5020 65308
rect 4956 65248 5020 65252
rect 5036 65308 5100 65312
rect 5036 65252 5040 65308
rect 5040 65252 5096 65308
rect 5096 65252 5100 65308
rect 5036 65248 5100 65252
rect 5116 65308 5180 65312
rect 5116 65252 5120 65308
rect 5120 65252 5176 65308
rect 5176 65252 5180 65308
rect 5116 65248 5180 65252
rect 106660 65308 106724 65312
rect 106660 65252 106664 65308
rect 106664 65252 106720 65308
rect 106720 65252 106724 65308
rect 106660 65248 106724 65252
rect 106740 65308 106804 65312
rect 106740 65252 106744 65308
rect 106744 65252 106800 65308
rect 106800 65252 106804 65308
rect 106740 65248 106804 65252
rect 106820 65308 106884 65312
rect 106820 65252 106824 65308
rect 106824 65252 106880 65308
rect 106880 65252 106884 65308
rect 106820 65248 106884 65252
rect 106900 65308 106964 65312
rect 106900 65252 106904 65308
rect 106904 65252 106960 65308
rect 106960 65252 106964 65308
rect 106900 65248 106964 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 105924 64764 105988 64768
rect 105924 64708 105928 64764
rect 105928 64708 105984 64764
rect 105984 64708 105988 64764
rect 105924 64704 105988 64708
rect 106004 64764 106068 64768
rect 106004 64708 106008 64764
rect 106008 64708 106064 64764
rect 106064 64708 106068 64764
rect 106004 64704 106068 64708
rect 106084 64764 106148 64768
rect 106084 64708 106088 64764
rect 106088 64708 106144 64764
rect 106144 64708 106148 64764
rect 106084 64704 106148 64708
rect 106164 64764 106228 64768
rect 106164 64708 106168 64764
rect 106168 64708 106224 64764
rect 106224 64708 106228 64764
rect 106164 64704 106228 64708
rect 4876 64220 4940 64224
rect 4876 64164 4880 64220
rect 4880 64164 4936 64220
rect 4936 64164 4940 64220
rect 4876 64160 4940 64164
rect 4956 64220 5020 64224
rect 4956 64164 4960 64220
rect 4960 64164 5016 64220
rect 5016 64164 5020 64220
rect 4956 64160 5020 64164
rect 5036 64220 5100 64224
rect 5036 64164 5040 64220
rect 5040 64164 5096 64220
rect 5096 64164 5100 64220
rect 5036 64160 5100 64164
rect 5116 64220 5180 64224
rect 5116 64164 5120 64220
rect 5120 64164 5176 64220
rect 5176 64164 5180 64220
rect 5116 64160 5180 64164
rect 106660 64220 106724 64224
rect 106660 64164 106664 64220
rect 106664 64164 106720 64220
rect 106720 64164 106724 64220
rect 106660 64160 106724 64164
rect 106740 64220 106804 64224
rect 106740 64164 106744 64220
rect 106744 64164 106800 64220
rect 106800 64164 106804 64220
rect 106740 64160 106804 64164
rect 106820 64220 106884 64224
rect 106820 64164 106824 64220
rect 106824 64164 106880 64220
rect 106880 64164 106884 64220
rect 106820 64160 106884 64164
rect 106900 64220 106964 64224
rect 106900 64164 106904 64220
rect 106904 64164 106960 64220
rect 106960 64164 106964 64220
rect 106900 64160 106964 64164
rect 38571 64092 38635 64156
rect 48544 64092 48608 64156
rect 56043 64092 56107 64156
rect 68523 64092 68587 64156
rect 58539 63956 58603 64020
rect 61056 63820 61120 63884
rect 95858 63820 95922 63884
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 105924 63676 105988 63680
rect 105924 63620 105928 63676
rect 105928 63620 105984 63676
rect 105984 63620 105988 63676
rect 105924 63616 105988 63620
rect 106004 63676 106068 63680
rect 106004 63620 106008 63676
rect 106008 63620 106064 63676
rect 106064 63620 106068 63676
rect 106004 63616 106068 63620
rect 106084 63676 106148 63680
rect 106084 63620 106088 63676
rect 106088 63620 106144 63676
rect 106144 63620 106148 63676
rect 106084 63616 106148 63620
rect 106164 63676 106228 63680
rect 106164 63620 106168 63676
rect 106168 63620 106224 63676
rect 106224 63620 106228 63676
rect 106164 63616 106228 63620
rect 4876 63132 4940 63136
rect 4876 63076 4880 63132
rect 4880 63076 4936 63132
rect 4936 63076 4940 63132
rect 4876 63072 4940 63076
rect 4956 63132 5020 63136
rect 4956 63076 4960 63132
rect 4960 63076 5016 63132
rect 5016 63076 5020 63132
rect 4956 63072 5020 63076
rect 5036 63132 5100 63136
rect 5036 63076 5040 63132
rect 5040 63076 5096 63132
rect 5096 63076 5100 63132
rect 5036 63072 5100 63076
rect 5116 63132 5180 63136
rect 5116 63076 5120 63132
rect 5120 63076 5176 63132
rect 5176 63076 5180 63132
rect 5116 63072 5180 63076
rect 106660 63132 106724 63136
rect 106660 63076 106664 63132
rect 106664 63076 106720 63132
rect 106720 63076 106724 63132
rect 106660 63072 106724 63076
rect 106740 63132 106804 63136
rect 106740 63076 106744 63132
rect 106744 63076 106800 63132
rect 106800 63076 106804 63132
rect 106740 63072 106804 63076
rect 106820 63132 106884 63136
rect 106820 63076 106824 63132
rect 106824 63076 106880 63132
rect 106880 63076 106884 63132
rect 106820 63072 106884 63076
rect 106900 63132 106964 63136
rect 106900 63076 106904 63132
rect 106904 63076 106960 63132
rect 106960 63076 106964 63132
rect 106900 63072 106964 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 105924 62588 105988 62592
rect 105924 62532 105928 62588
rect 105928 62532 105984 62588
rect 105984 62532 105988 62588
rect 105924 62528 105988 62532
rect 106004 62588 106068 62592
rect 106004 62532 106008 62588
rect 106008 62532 106064 62588
rect 106064 62532 106068 62588
rect 106004 62528 106068 62532
rect 106084 62588 106148 62592
rect 106084 62532 106088 62588
rect 106088 62532 106144 62588
rect 106144 62532 106148 62588
rect 106084 62528 106148 62532
rect 106164 62588 106228 62592
rect 106164 62532 106168 62588
rect 106168 62532 106224 62588
rect 106224 62532 106228 62588
rect 106164 62528 106228 62532
rect 4876 62044 4940 62048
rect 4876 61988 4880 62044
rect 4880 61988 4936 62044
rect 4936 61988 4940 62044
rect 4876 61984 4940 61988
rect 4956 62044 5020 62048
rect 4956 61988 4960 62044
rect 4960 61988 5016 62044
rect 5016 61988 5020 62044
rect 4956 61984 5020 61988
rect 5036 62044 5100 62048
rect 5036 61988 5040 62044
rect 5040 61988 5096 62044
rect 5096 61988 5100 62044
rect 5036 61984 5100 61988
rect 5116 62044 5180 62048
rect 5116 61988 5120 62044
rect 5120 61988 5176 62044
rect 5176 61988 5180 62044
rect 5116 61984 5180 61988
rect 106660 62044 106724 62048
rect 106660 61988 106664 62044
rect 106664 61988 106720 62044
rect 106720 61988 106724 62044
rect 106660 61984 106724 61988
rect 106740 62044 106804 62048
rect 106740 61988 106744 62044
rect 106744 61988 106800 62044
rect 106800 61988 106804 62044
rect 106740 61984 106804 61988
rect 106820 62044 106884 62048
rect 106820 61988 106824 62044
rect 106824 61988 106880 62044
rect 106880 61988 106884 62044
rect 106820 61984 106884 61988
rect 106900 62044 106964 62048
rect 106900 61988 106904 62044
rect 106904 61988 106960 62044
rect 106960 61988 106964 62044
rect 106900 61984 106964 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 105924 61500 105988 61504
rect 105924 61444 105928 61500
rect 105928 61444 105984 61500
rect 105984 61444 105988 61500
rect 105924 61440 105988 61444
rect 106004 61500 106068 61504
rect 106004 61444 106008 61500
rect 106008 61444 106064 61500
rect 106064 61444 106068 61500
rect 106004 61440 106068 61444
rect 106084 61500 106148 61504
rect 106084 61444 106088 61500
rect 106088 61444 106144 61500
rect 106144 61444 106148 61500
rect 106084 61440 106148 61444
rect 106164 61500 106228 61504
rect 106164 61444 106168 61500
rect 106168 61444 106224 61500
rect 106224 61444 106228 61500
rect 106164 61440 106228 61444
rect 4876 60956 4940 60960
rect 4876 60900 4880 60956
rect 4880 60900 4936 60956
rect 4936 60900 4940 60956
rect 4876 60896 4940 60900
rect 4956 60956 5020 60960
rect 4956 60900 4960 60956
rect 4960 60900 5016 60956
rect 5016 60900 5020 60956
rect 4956 60896 5020 60900
rect 5036 60956 5100 60960
rect 5036 60900 5040 60956
rect 5040 60900 5096 60956
rect 5096 60900 5100 60956
rect 5036 60896 5100 60900
rect 5116 60956 5180 60960
rect 5116 60900 5120 60956
rect 5120 60900 5176 60956
rect 5176 60900 5180 60956
rect 5116 60896 5180 60900
rect 106660 60956 106724 60960
rect 106660 60900 106664 60956
rect 106664 60900 106720 60956
rect 106720 60900 106724 60956
rect 106660 60896 106724 60900
rect 106740 60956 106804 60960
rect 106740 60900 106744 60956
rect 106744 60900 106800 60956
rect 106800 60900 106804 60956
rect 106740 60896 106804 60900
rect 106820 60956 106884 60960
rect 106820 60900 106824 60956
rect 106824 60900 106880 60956
rect 106880 60900 106884 60956
rect 106820 60896 106884 60900
rect 106900 60956 106964 60960
rect 106900 60900 106904 60956
rect 106904 60900 106960 60956
rect 106960 60900 106964 60956
rect 106900 60896 106964 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 105924 60412 105988 60416
rect 105924 60356 105928 60412
rect 105928 60356 105984 60412
rect 105984 60356 105988 60412
rect 105924 60352 105988 60356
rect 106004 60412 106068 60416
rect 106004 60356 106008 60412
rect 106008 60356 106064 60412
rect 106064 60356 106068 60412
rect 106004 60352 106068 60356
rect 106084 60412 106148 60416
rect 106084 60356 106088 60412
rect 106088 60356 106144 60412
rect 106144 60356 106148 60412
rect 106084 60352 106148 60356
rect 106164 60412 106228 60416
rect 106164 60356 106168 60412
rect 106168 60356 106224 60412
rect 106224 60356 106228 60412
rect 106164 60352 106228 60356
rect 4876 59868 4940 59872
rect 4876 59812 4880 59868
rect 4880 59812 4936 59868
rect 4936 59812 4940 59868
rect 4876 59808 4940 59812
rect 4956 59868 5020 59872
rect 4956 59812 4960 59868
rect 4960 59812 5016 59868
rect 5016 59812 5020 59868
rect 4956 59808 5020 59812
rect 5036 59868 5100 59872
rect 5036 59812 5040 59868
rect 5040 59812 5096 59868
rect 5096 59812 5100 59868
rect 5036 59808 5100 59812
rect 5116 59868 5180 59872
rect 5116 59812 5120 59868
rect 5120 59812 5176 59868
rect 5176 59812 5180 59868
rect 5116 59808 5180 59812
rect 106660 59868 106724 59872
rect 106660 59812 106664 59868
rect 106664 59812 106720 59868
rect 106720 59812 106724 59868
rect 106660 59808 106724 59812
rect 106740 59868 106804 59872
rect 106740 59812 106744 59868
rect 106744 59812 106800 59868
rect 106800 59812 106804 59868
rect 106740 59808 106804 59812
rect 106820 59868 106884 59872
rect 106820 59812 106824 59868
rect 106824 59812 106880 59868
rect 106880 59812 106884 59868
rect 106820 59808 106884 59812
rect 106900 59868 106964 59872
rect 106900 59812 106904 59868
rect 106904 59812 106960 59868
rect 106960 59812 106964 59868
rect 106900 59808 106964 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 105924 59324 105988 59328
rect 105924 59268 105928 59324
rect 105928 59268 105984 59324
rect 105984 59268 105988 59324
rect 105924 59264 105988 59268
rect 106004 59324 106068 59328
rect 106004 59268 106008 59324
rect 106008 59268 106064 59324
rect 106064 59268 106068 59324
rect 106004 59264 106068 59268
rect 106084 59324 106148 59328
rect 106084 59268 106088 59324
rect 106088 59268 106144 59324
rect 106144 59268 106148 59324
rect 106084 59264 106148 59268
rect 106164 59324 106228 59328
rect 106164 59268 106168 59324
rect 106168 59268 106224 59324
rect 106224 59268 106228 59324
rect 106164 59264 106228 59268
rect 4876 58780 4940 58784
rect 4876 58724 4880 58780
rect 4880 58724 4936 58780
rect 4936 58724 4940 58780
rect 4876 58720 4940 58724
rect 4956 58780 5020 58784
rect 4956 58724 4960 58780
rect 4960 58724 5016 58780
rect 5016 58724 5020 58780
rect 4956 58720 5020 58724
rect 5036 58780 5100 58784
rect 5036 58724 5040 58780
rect 5040 58724 5096 58780
rect 5096 58724 5100 58780
rect 5036 58720 5100 58724
rect 5116 58780 5180 58784
rect 5116 58724 5120 58780
rect 5120 58724 5176 58780
rect 5176 58724 5180 58780
rect 5116 58720 5180 58724
rect 106660 58780 106724 58784
rect 106660 58724 106664 58780
rect 106664 58724 106720 58780
rect 106720 58724 106724 58780
rect 106660 58720 106724 58724
rect 106740 58780 106804 58784
rect 106740 58724 106744 58780
rect 106744 58724 106800 58780
rect 106800 58724 106804 58780
rect 106740 58720 106804 58724
rect 106820 58780 106884 58784
rect 106820 58724 106824 58780
rect 106824 58724 106880 58780
rect 106880 58724 106884 58780
rect 106820 58720 106884 58724
rect 106900 58780 106964 58784
rect 106900 58724 106904 58780
rect 106904 58724 106960 58780
rect 106960 58724 106964 58780
rect 106900 58720 106964 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 105924 58236 105988 58240
rect 105924 58180 105928 58236
rect 105928 58180 105984 58236
rect 105984 58180 105988 58236
rect 105924 58176 105988 58180
rect 106004 58236 106068 58240
rect 106004 58180 106008 58236
rect 106008 58180 106064 58236
rect 106064 58180 106068 58236
rect 106004 58176 106068 58180
rect 106084 58236 106148 58240
rect 106084 58180 106088 58236
rect 106088 58180 106144 58236
rect 106144 58180 106148 58236
rect 106084 58176 106148 58180
rect 106164 58236 106228 58240
rect 106164 58180 106168 58236
rect 106168 58180 106224 58236
rect 106224 58180 106228 58236
rect 106164 58176 106228 58180
rect 4876 57692 4940 57696
rect 4876 57636 4880 57692
rect 4880 57636 4936 57692
rect 4936 57636 4940 57692
rect 4876 57632 4940 57636
rect 4956 57692 5020 57696
rect 4956 57636 4960 57692
rect 4960 57636 5016 57692
rect 5016 57636 5020 57692
rect 4956 57632 5020 57636
rect 5036 57692 5100 57696
rect 5036 57636 5040 57692
rect 5040 57636 5096 57692
rect 5096 57636 5100 57692
rect 5036 57632 5100 57636
rect 5116 57692 5180 57696
rect 5116 57636 5120 57692
rect 5120 57636 5176 57692
rect 5176 57636 5180 57692
rect 5116 57632 5180 57636
rect 106660 57692 106724 57696
rect 106660 57636 106664 57692
rect 106664 57636 106720 57692
rect 106720 57636 106724 57692
rect 106660 57632 106724 57636
rect 106740 57692 106804 57696
rect 106740 57636 106744 57692
rect 106744 57636 106800 57692
rect 106800 57636 106804 57692
rect 106740 57632 106804 57636
rect 106820 57692 106884 57696
rect 106820 57636 106824 57692
rect 106824 57636 106880 57692
rect 106880 57636 106884 57692
rect 106820 57632 106884 57636
rect 106900 57692 106964 57696
rect 106900 57636 106904 57692
rect 106904 57636 106960 57692
rect 106960 57636 106964 57692
rect 106900 57632 106964 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 105924 57148 105988 57152
rect 105924 57092 105928 57148
rect 105928 57092 105984 57148
rect 105984 57092 105988 57148
rect 105924 57088 105988 57092
rect 106004 57148 106068 57152
rect 106004 57092 106008 57148
rect 106008 57092 106064 57148
rect 106064 57092 106068 57148
rect 106004 57088 106068 57092
rect 106084 57148 106148 57152
rect 106084 57092 106088 57148
rect 106088 57092 106144 57148
rect 106144 57092 106148 57148
rect 106084 57088 106148 57092
rect 106164 57148 106228 57152
rect 106164 57092 106168 57148
rect 106168 57092 106224 57148
rect 106224 57092 106228 57148
rect 106164 57088 106228 57092
rect 4876 56604 4940 56608
rect 4876 56548 4880 56604
rect 4880 56548 4936 56604
rect 4936 56548 4940 56604
rect 4876 56544 4940 56548
rect 4956 56604 5020 56608
rect 4956 56548 4960 56604
rect 4960 56548 5016 56604
rect 5016 56548 5020 56604
rect 4956 56544 5020 56548
rect 5036 56604 5100 56608
rect 5036 56548 5040 56604
rect 5040 56548 5096 56604
rect 5096 56548 5100 56604
rect 5036 56544 5100 56548
rect 5116 56604 5180 56608
rect 5116 56548 5120 56604
rect 5120 56548 5176 56604
rect 5176 56548 5180 56604
rect 5116 56544 5180 56548
rect 106660 56604 106724 56608
rect 106660 56548 106664 56604
rect 106664 56548 106720 56604
rect 106720 56548 106724 56604
rect 106660 56544 106724 56548
rect 106740 56604 106804 56608
rect 106740 56548 106744 56604
rect 106744 56548 106800 56604
rect 106800 56548 106804 56604
rect 106740 56544 106804 56548
rect 106820 56604 106884 56608
rect 106820 56548 106824 56604
rect 106824 56548 106880 56604
rect 106880 56548 106884 56604
rect 106820 56544 106884 56548
rect 106900 56604 106964 56608
rect 106900 56548 106904 56604
rect 106904 56548 106960 56604
rect 106960 56548 106964 56604
rect 106900 56544 106964 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 105924 56060 105988 56064
rect 105924 56004 105928 56060
rect 105928 56004 105984 56060
rect 105984 56004 105988 56060
rect 105924 56000 105988 56004
rect 106004 56060 106068 56064
rect 106004 56004 106008 56060
rect 106008 56004 106064 56060
rect 106064 56004 106068 56060
rect 106004 56000 106068 56004
rect 106084 56060 106148 56064
rect 106084 56004 106088 56060
rect 106088 56004 106144 56060
rect 106144 56004 106148 56060
rect 106084 56000 106148 56004
rect 106164 56060 106228 56064
rect 106164 56004 106168 56060
rect 106168 56004 106224 56060
rect 106224 56004 106228 56060
rect 106164 56000 106228 56004
rect 4876 55516 4940 55520
rect 4876 55460 4880 55516
rect 4880 55460 4936 55516
rect 4936 55460 4940 55516
rect 4876 55456 4940 55460
rect 4956 55516 5020 55520
rect 4956 55460 4960 55516
rect 4960 55460 5016 55516
rect 5016 55460 5020 55516
rect 4956 55456 5020 55460
rect 5036 55516 5100 55520
rect 5036 55460 5040 55516
rect 5040 55460 5096 55516
rect 5096 55460 5100 55516
rect 5036 55456 5100 55460
rect 5116 55516 5180 55520
rect 5116 55460 5120 55516
rect 5120 55460 5176 55516
rect 5176 55460 5180 55516
rect 5116 55456 5180 55460
rect 106660 55516 106724 55520
rect 106660 55460 106664 55516
rect 106664 55460 106720 55516
rect 106720 55460 106724 55516
rect 106660 55456 106724 55460
rect 106740 55516 106804 55520
rect 106740 55460 106744 55516
rect 106744 55460 106800 55516
rect 106800 55460 106804 55516
rect 106740 55456 106804 55460
rect 106820 55516 106884 55520
rect 106820 55460 106824 55516
rect 106824 55460 106880 55516
rect 106880 55460 106884 55516
rect 106820 55456 106884 55460
rect 106900 55516 106964 55520
rect 106900 55460 106904 55516
rect 106904 55460 106960 55516
rect 106960 55460 106964 55516
rect 106900 55456 106964 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 105924 54972 105988 54976
rect 105924 54916 105928 54972
rect 105928 54916 105984 54972
rect 105984 54916 105988 54972
rect 105924 54912 105988 54916
rect 106004 54972 106068 54976
rect 106004 54916 106008 54972
rect 106008 54916 106064 54972
rect 106064 54916 106068 54972
rect 106004 54912 106068 54916
rect 106084 54972 106148 54976
rect 106084 54916 106088 54972
rect 106088 54916 106144 54972
rect 106144 54916 106148 54972
rect 106084 54912 106148 54916
rect 106164 54972 106228 54976
rect 106164 54916 106168 54972
rect 106168 54916 106224 54972
rect 106224 54916 106228 54972
rect 106164 54912 106228 54916
rect 4876 54428 4940 54432
rect 4876 54372 4880 54428
rect 4880 54372 4936 54428
rect 4936 54372 4940 54428
rect 4876 54368 4940 54372
rect 4956 54428 5020 54432
rect 4956 54372 4960 54428
rect 4960 54372 5016 54428
rect 5016 54372 5020 54428
rect 4956 54368 5020 54372
rect 5036 54428 5100 54432
rect 5036 54372 5040 54428
rect 5040 54372 5096 54428
rect 5096 54372 5100 54428
rect 5036 54368 5100 54372
rect 5116 54428 5180 54432
rect 5116 54372 5120 54428
rect 5120 54372 5176 54428
rect 5176 54372 5180 54428
rect 5116 54368 5180 54372
rect 106660 54428 106724 54432
rect 106660 54372 106664 54428
rect 106664 54372 106720 54428
rect 106720 54372 106724 54428
rect 106660 54368 106724 54372
rect 106740 54428 106804 54432
rect 106740 54372 106744 54428
rect 106744 54372 106800 54428
rect 106800 54372 106804 54428
rect 106740 54368 106804 54372
rect 106820 54428 106884 54432
rect 106820 54372 106824 54428
rect 106824 54372 106880 54428
rect 106880 54372 106884 54428
rect 106820 54368 106884 54372
rect 106900 54428 106964 54432
rect 106900 54372 106904 54428
rect 106904 54372 106960 54428
rect 106960 54372 106964 54428
rect 106900 54368 106964 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 105924 53884 105988 53888
rect 105924 53828 105928 53884
rect 105928 53828 105984 53884
rect 105984 53828 105988 53884
rect 105924 53824 105988 53828
rect 106004 53884 106068 53888
rect 106004 53828 106008 53884
rect 106008 53828 106064 53884
rect 106064 53828 106068 53884
rect 106004 53824 106068 53828
rect 106084 53884 106148 53888
rect 106084 53828 106088 53884
rect 106088 53828 106144 53884
rect 106144 53828 106148 53884
rect 106084 53824 106148 53828
rect 106164 53884 106228 53888
rect 106164 53828 106168 53884
rect 106168 53828 106224 53884
rect 106224 53828 106228 53884
rect 106164 53824 106228 53828
rect 4876 53340 4940 53344
rect 4876 53284 4880 53340
rect 4880 53284 4936 53340
rect 4936 53284 4940 53340
rect 4876 53280 4940 53284
rect 4956 53340 5020 53344
rect 4956 53284 4960 53340
rect 4960 53284 5016 53340
rect 5016 53284 5020 53340
rect 4956 53280 5020 53284
rect 5036 53340 5100 53344
rect 5036 53284 5040 53340
rect 5040 53284 5096 53340
rect 5096 53284 5100 53340
rect 5036 53280 5100 53284
rect 5116 53340 5180 53344
rect 5116 53284 5120 53340
rect 5120 53284 5176 53340
rect 5176 53284 5180 53340
rect 5116 53280 5180 53284
rect 106660 53340 106724 53344
rect 106660 53284 106664 53340
rect 106664 53284 106720 53340
rect 106720 53284 106724 53340
rect 106660 53280 106724 53284
rect 106740 53340 106804 53344
rect 106740 53284 106744 53340
rect 106744 53284 106800 53340
rect 106800 53284 106804 53340
rect 106740 53280 106804 53284
rect 106820 53340 106884 53344
rect 106820 53284 106824 53340
rect 106824 53284 106880 53340
rect 106880 53284 106884 53340
rect 106820 53280 106884 53284
rect 106900 53340 106964 53344
rect 106900 53284 106904 53340
rect 106904 53284 106960 53340
rect 106960 53284 106964 53340
rect 106900 53280 106964 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 105924 52796 105988 52800
rect 105924 52740 105928 52796
rect 105928 52740 105984 52796
rect 105984 52740 105988 52796
rect 105924 52736 105988 52740
rect 106004 52796 106068 52800
rect 106004 52740 106008 52796
rect 106008 52740 106064 52796
rect 106064 52740 106068 52796
rect 106004 52736 106068 52740
rect 106084 52796 106148 52800
rect 106084 52740 106088 52796
rect 106088 52740 106144 52796
rect 106144 52740 106148 52796
rect 106084 52736 106148 52740
rect 106164 52796 106228 52800
rect 106164 52740 106168 52796
rect 106168 52740 106224 52796
rect 106224 52740 106228 52796
rect 106164 52736 106228 52740
rect 4876 52252 4940 52256
rect 4876 52196 4880 52252
rect 4880 52196 4936 52252
rect 4936 52196 4940 52252
rect 4876 52192 4940 52196
rect 4956 52252 5020 52256
rect 4956 52196 4960 52252
rect 4960 52196 5016 52252
rect 5016 52196 5020 52252
rect 4956 52192 5020 52196
rect 5036 52252 5100 52256
rect 5036 52196 5040 52252
rect 5040 52196 5096 52252
rect 5096 52196 5100 52252
rect 5036 52192 5100 52196
rect 5116 52252 5180 52256
rect 5116 52196 5120 52252
rect 5120 52196 5176 52252
rect 5176 52196 5180 52252
rect 5116 52192 5180 52196
rect 106660 52252 106724 52256
rect 106660 52196 106664 52252
rect 106664 52196 106720 52252
rect 106720 52196 106724 52252
rect 106660 52192 106724 52196
rect 106740 52252 106804 52256
rect 106740 52196 106744 52252
rect 106744 52196 106800 52252
rect 106800 52196 106804 52252
rect 106740 52192 106804 52196
rect 106820 52252 106884 52256
rect 106820 52196 106824 52252
rect 106824 52196 106880 52252
rect 106880 52196 106884 52252
rect 106820 52192 106884 52196
rect 106900 52252 106964 52256
rect 106900 52196 106904 52252
rect 106904 52196 106960 52252
rect 106960 52196 106964 52252
rect 106900 52192 106964 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 105924 51708 105988 51712
rect 105924 51652 105928 51708
rect 105928 51652 105984 51708
rect 105984 51652 105988 51708
rect 105924 51648 105988 51652
rect 106004 51708 106068 51712
rect 106004 51652 106008 51708
rect 106008 51652 106064 51708
rect 106064 51652 106068 51708
rect 106004 51648 106068 51652
rect 106084 51708 106148 51712
rect 106084 51652 106088 51708
rect 106088 51652 106144 51708
rect 106144 51652 106148 51708
rect 106084 51648 106148 51652
rect 106164 51708 106228 51712
rect 106164 51652 106168 51708
rect 106168 51652 106224 51708
rect 106224 51652 106228 51708
rect 106164 51648 106228 51652
rect 4876 51164 4940 51168
rect 4876 51108 4880 51164
rect 4880 51108 4936 51164
rect 4936 51108 4940 51164
rect 4876 51104 4940 51108
rect 4956 51164 5020 51168
rect 4956 51108 4960 51164
rect 4960 51108 5016 51164
rect 5016 51108 5020 51164
rect 4956 51104 5020 51108
rect 5036 51164 5100 51168
rect 5036 51108 5040 51164
rect 5040 51108 5096 51164
rect 5096 51108 5100 51164
rect 5036 51104 5100 51108
rect 5116 51164 5180 51168
rect 5116 51108 5120 51164
rect 5120 51108 5176 51164
rect 5176 51108 5180 51164
rect 5116 51104 5180 51108
rect 106660 51164 106724 51168
rect 106660 51108 106664 51164
rect 106664 51108 106720 51164
rect 106720 51108 106724 51164
rect 106660 51104 106724 51108
rect 106740 51164 106804 51168
rect 106740 51108 106744 51164
rect 106744 51108 106800 51164
rect 106800 51108 106804 51164
rect 106740 51104 106804 51108
rect 106820 51164 106884 51168
rect 106820 51108 106824 51164
rect 106824 51108 106880 51164
rect 106880 51108 106884 51164
rect 106820 51104 106884 51108
rect 106900 51164 106964 51168
rect 106900 51108 106904 51164
rect 106904 51108 106960 51164
rect 106960 51108 106964 51164
rect 106900 51104 106964 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 105924 50620 105988 50624
rect 105924 50564 105928 50620
rect 105928 50564 105984 50620
rect 105984 50564 105988 50620
rect 105924 50560 105988 50564
rect 106004 50620 106068 50624
rect 106004 50564 106008 50620
rect 106008 50564 106064 50620
rect 106064 50564 106068 50620
rect 106004 50560 106068 50564
rect 106084 50620 106148 50624
rect 106084 50564 106088 50620
rect 106088 50564 106144 50620
rect 106144 50564 106148 50620
rect 106084 50560 106148 50564
rect 106164 50620 106228 50624
rect 106164 50564 106168 50620
rect 106168 50564 106224 50620
rect 106224 50564 106228 50620
rect 106164 50560 106228 50564
rect 4876 50076 4940 50080
rect 4876 50020 4880 50076
rect 4880 50020 4936 50076
rect 4936 50020 4940 50076
rect 4876 50016 4940 50020
rect 4956 50076 5020 50080
rect 4956 50020 4960 50076
rect 4960 50020 5016 50076
rect 5016 50020 5020 50076
rect 4956 50016 5020 50020
rect 5036 50076 5100 50080
rect 5036 50020 5040 50076
rect 5040 50020 5096 50076
rect 5096 50020 5100 50076
rect 5036 50016 5100 50020
rect 5116 50076 5180 50080
rect 5116 50020 5120 50076
rect 5120 50020 5176 50076
rect 5176 50020 5180 50076
rect 5116 50016 5180 50020
rect 106660 50076 106724 50080
rect 106660 50020 106664 50076
rect 106664 50020 106720 50076
rect 106720 50020 106724 50076
rect 106660 50016 106724 50020
rect 106740 50076 106804 50080
rect 106740 50020 106744 50076
rect 106744 50020 106800 50076
rect 106800 50020 106804 50076
rect 106740 50016 106804 50020
rect 106820 50076 106884 50080
rect 106820 50020 106824 50076
rect 106824 50020 106880 50076
rect 106880 50020 106884 50076
rect 106820 50016 106884 50020
rect 106900 50076 106964 50080
rect 106900 50020 106904 50076
rect 106904 50020 106960 50076
rect 106960 50020 106964 50076
rect 106900 50016 106964 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 105924 49532 105988 49536
rect 105924 49476 105928 49532
rect 105928 49476 105984 49532
rect 105984 49476 105988 49532
rect 105924 49472 105988 49476
rect 106004 49532 106068 49536
rect 106004 49476 106008 49532
rect 106008 49476 106064 49532
rect 106064 49476 106068 49532
rect 106004 49472 106068 49476
rect 106084 49532 106148 49536
rect 106084 49476 106088 49532
rect 106088 49476 106144 49532
rect 106144 49476 106148 49532
rect 106084 49472 106148 49476
rect 106164 49532 106228 49536
rect 106164 49476 106168 49532
rect 106168 49476 106224 49532
rect 106224 49476 106228 49532
rect 106164 49472 106228 49476
rect 4876 48988 4940 48992
rect 4876 48932 4880 48988
rect 4880 48932 4936 48988
rect 4936 48932 4940 48988
rect 4876 48928 4940 48932
rect 4956 48988 5020 48992
rect 4956 48932 4960 48988
rect 4960 48932 5016 48988
rect 5016 48932 5020 48988
rect 4956 48928 5020 48932
rect 5036 48988 5100 48992
rect 5036 48932 5040 48988
rect 5040 48932 5096 48988
rect 5096 48932 5100 48988
rect 5036 48928 5100 48932
rect 5116 48988 5180 48992
rect 5116 48932 5120 48988
rect 5120 48932 5176 48988
rect 5176 48932 5180 48988
rect 5116 48928 5180 48932
rect 106660 48988 106724 48992
rect 106660 48932 106664 48988
rect 106664 48932 106720 48988
rect 106720 48932 106724 48988
rect 106660 48928 106724 48932
rect 106740 48988 106804 48992
rect 106740 48932 106744 48988
rect 106744 48932 106800 48988
rect 106800 48932 106804 48988
rect 106740 48928 106804 48932
rect 106820 48988 106884 48992
rect 106820 48932 106824 48988
rect 106824 48932 106880 48988
rect 106880 48932 106884 48988
rect 106820 48928 106884 48932
rect 106900 48988 106964 48992
rect 106900 48932 106904 48988
rect 106904 48932 106960 48988
rect 106960 48932 106964 48988
rect 106900 48928 106964 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 105924 48444 105988 48448
rect 105924 48388 105928 48444
rect 105928 48388 105984 48444
rect 105984 48388 105988 48444
rect 105924 48384 105988 48388
rect 106004 48444 106068 48448
rect 106004 48388 106008 48444
rect 106008 48388 106064 48444
rect 106064 48388 106068 48444
rect 106004 48384 106068 48388
rect 106084 48444 106148 48448
rect 106084 48388 106088 48444
rect 106088 48388 106144 48444
rect 106144 48388 106148 48444
rect 106084 48384 106148 48388
rect 106164 48444 106228 48448
rect 106164 48388 106168 48444
rect 106168 48388 106224 48444
rect 106224 48388 106228 48444
rect 106164 48384 106228 48388
rect 4876 47900 4940 47904
rect 4876 47844 4880 47900
rect 4880 47844 4936 47900
rect 4936 47844 4940 47900
rect 4876 47840 4940 47844
rect 4956 47900 5020 47904
rect 4956 47844 4960 47900
rect 4960 47844 5016 47900
rect 5016 47844 5020 47900
rect 4956 47840 5020 47844
rect 5036 47900 5100 47904
rect 5036 47844 5040 47900
rect 5040 47844 5096 47900
rect 5096 47844 5100 47900
rect 5036 47840 5100 47844
rect 5116 47900 5180 47904
rect 5116 47844 5120 47900
rect 5120 47844 5176 47900
rect 5176 47844 5180 47900
rect 5116 47840 5180 47844
rect 106660 47900 106724 47904
rect 106660 47844 106664 47900
rect 106664 47844 106720 47900
rect 106720 47844 106724 47900
rect 106660 47840 106724 47844
rect 106740 47900 106804 47904
rect 106740 47844 106744 47900
rect 106744 47844 106800 47900
rect 106800 47844 106804 47900
rect 106740 47840 106804 47844
rect 106820 47900 106884 47904
rect 106820 47844 106824 47900
rect 106824 47844 106880 47900
rect 106880 47844 106884 47900
rect 106820 47840 106884 47844
rect 106900 47900 106964 47904
rect 106900 47844 106904 47900
rect 106904 47844 106960 47900
rect 106960 47844 106964 47900
rect 106900 47840 106964 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 105924 47356 105988 47360
rect 105924 47300 105928 47356
rect 105928 47300 105984 47356
rect 105984 47300 105988 47356
rect 105924 47296 105988 47300
rect 106004 47356 106068 47360
rect 106004 47300 106008 47356
rect 106008 47300 106064 47356
rect 106064 47300 106068 47356
rect 106004 47296 106068 47300
rect 106084 47356 106148 47360
rect 106084 47300 106088 47356
rect 106088 47300 106144 47356
rect 106144 47300 106148 47356
rect 106084 47296 106148 47300
rect 106164 47356 106228 47360
rect 106164 47300 106168 47356
rect 106168 47300 106224 47356
rect 106224 47300 106228 47356
rect 106164 47296 106228 47300
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 106660 46812 106724 46816
rect 106660 46756 106664 46812
rect 106664 46756 106720 46812
rect 106720 46756 106724 46812
rect 106660 46752 106724 46756
rect 106740 46812 106804 46816
rect 106740 46756 106744 46812
rect 106744 46756 106800 46812
rect 106800 46756 106804 46812
rect 106740 46752 106804 46756
rect 106820 46812 106884 46816
rect 106820 46756 106824 46812
rect 106824 46756 106880 46812
rect 106880 46756 106884 46812
rect 106820 46752 106884 46756
rect 106900 46812 106964 46816
rect 106900 46756 106904 46812
rect 106904 46756 106960 46812
rect 106960 46756 106964 46812
rect 106900 46752 106964 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 105924 46268 105988 46272
rect 105924 46212 105928 46268
rect 105928 46212 105984 46268
rect 105984 46212 105988 46268
rect 105924 46208 105988 46212
rect 106004 46268 106068 46272
rect 106004 46212 106008 46268
rect 106008 46212 106064 46268
rect 106064 46212 106068 46268
rect 106004 46208 106068 46212
rect 106084 46268 106148 46272
rect 106084 46212 106088 46268
rect 106088 46212 106144 46268
rect 106144 46212 106148 46268
rect 106084 46208 106148 46212
rect 106164 46268 106228 46272
rect 106164 46212 106168 46268
rect 106168 46212 106224 46268
rect 106224 46212 106228 46268
rect 106164 46208 106228 46212
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 106660 45724 106724 45728
rect 106660 45668 106664 45724
rect 106664 45668 106720 45724
rect 106720 45668 106724 45724
rect 106660 45664 106724 45668
rect 106740 45724 106804 45728
rect 106740 45668 106744 45724
rect 106744 45668 106800 45724
rect 106800 45668 106804 45724
rect 106740 45664 106804 45668
rect 106820 45724 106884 45728
rect 106820 45668 106824 45724
rect 106824 45668 106880 45724
rect 106880 45668 106884 45724
rect 106820 45664 106884 45668
rect 106900 45724 106964 45728
rect 106900 45668 106904 45724
rect 106904 45668 106960 45724
rect 106960 45668 106964 45724
rect 106900 45664 106964 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 105924 45180 105988 45184
rect 105924 45124 105928 45180
rect 105928 45124 105984 45180
rect 105984 45124 105988 45180
rect 105924 45120 105988 45124
rect 106004 45180 106068 45184
rect 106004 45124 106008 45180
rect 106008 45124 106064 45180
rect 106064 45124 106068 45180
rect 106004 45120 106068 45124
rect 106084 45180 106148 45184
rect 106084 45124 106088 45180
rect 106088 45124 106144 45180
rect 106144 45124 106148 45180
rect 106084 45120 106148 45124
rect 106164 45180 106228 45184
rect 106164 45124 106168 45180
rect 106168 45124 106224 45180
rect 106224 45124 106228 45180
rect 106164 45120 106228 45124
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 106660 44636 106724 44640
rect 106660 44580 106664 44636
rect 106664 44580 106720 44636
rect 106720 44580 106724 44636
rect 106660 44576 106724 44580
rect 106740 44636 106804 44640
rect 106740 44580 106744 44636
rect 106744 44580 106800 44636
rect 106800 44580 106804 44636
rect 106740 44576 106804 44580
rect 106820 44636 106884 44640
rect 106820 44580 106824 44636
rect 106824 44580 106880 44636
rect 106880 44580 106884 44636
rect 106820 44576 106884 44580
rect 106900 44636 106964 44640
rect 106900 44580 106904 44636
rect 106904 44580 106960 44636
rect 106960 44580 106964 44636
rect 106900 44576 106964 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 105924 44092 105988 44096
rect 105924 44036 105928 44092
rect 105928 44036 105984 44092
rect 105984 44036 105988 44092
rect 105924 44032 105988 44036
rect 106004 44092 106068 44096
rect 106004 44036 106008 44092
rect 106008 44036 106064 44092
rect 106064 44036 106068 44092
rect 106004 44032 106068 44036
rect 106084 44092 106148 44096
rect 106084 44036 106088 44092
rect 106088 44036 106144 44092
rect 106144 44036 106148 44092
rect 106084 44032 106148 44036
rect 106164 44092 106228 44096
rect 106164 44036 106168 44092
rect 106168 44036 106224 44092
rect 106224 44036 106228 44092
rect 106164 44032 106228 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 106660 43548 106724 43552
rect 106660 43492 106664 43548
rect 106664 43492 106720 43548
rect 106720 43492 106724 43548
rect 106660 43488 106724 43492
rect 106740 43548 106804 43552
rect 106740 43492 106744 43548
rect 106744 43492 106800 43548
rect 106800 43492 106804 43548
rect 106740 43488 106804 43492
rect 106820 43548 106884 43552
rect 106820 43492 106824 43548
rect 106824 43492 106880 43548
rect 106880 43492 106884 43548
rect 106820 43488 106884 43492
rect 106900 43548 106964 43552
rect 106900 43492 106904 43548
rect 106904 43492 106960 43548
rect 106960 43492 106964 43548
rect 106900 43488 106964 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 105924 43004 105988 43008
rect 105924 42948 105928 43004
rect 105928 42948 105984 43004
rect 105984 42948 105988 43004
rect 105924 42944 105988 42948
rect 106004 43004 106068 43008
rect 106004 42948 106008 43004
rect 106008 42948 106064 43004
rect 106064 42948 106068 43004
rect 106004 42944 106068 42948
rect 106084 43004 106148 43008
rect 106084 42948 106088 43004
rect 106088 42948 106144 43004
rect 106144 42948 106148 43004
rect 106084 42944 106148 42948
rect 106164 43004 106228 43008
rect 106164 42948 106168 43004
rect 106168 42948 106224 43004
rect 106224 42948 106228 43004
rect 106164 42944 106228 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 106660 42460 106724 42464
rect 106660 42404 106664 42460
rect 106664 42404 106720 42460
rect 106720 42404 106724 42460
rect 106660 42400 106724 42404
rect 106740 42460 106804 42464
rect 106740 42404 106744 42460
rect 106744 42404 106800 42460
rect 106800 42404 106804 42460
rect 106740 42400 106804 42404
rect 106820 42460 106884 42464
rect 106820 42404 106824 42460
rect 106824 42404 106880 42460
rect 106880 42404 106884 42460
rect 106820 42400 106884 42404
rect 106900 42460 106964 42464
rect 106900 42404 106904 42460
rect 106904 42404 106960 42460
rect 106960 42404 106964 42460
rect 106900 42400 106964 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 105924 41916 105988 41920
rect 105924 41860 105928 41916
rect 105928 41860 105984 41916
rect 105984 41860 105988 41916
rect 105924 41856 105988 41860
rect 106004 41916 106068 41920
rect 106004 41860 106008 41916
rect 106008 41860 106064 41916
rect 106064 41860 106068 41916
rect 106004 41856 106068 41860
rect 106084 41916 106148 41920
rect 106084 41860 106088 41916
rect 106088 41860 106144 41916
rect 106144 41860 106148 41916
rect 106084 41856 106148 41860
rect 106164 41916 106228 41920
rect 106164 41860 106168 41916
rect 106168 41860 106224 41916
rect 106224 41860 106228 41916
rect 106164 41856 106228 41860
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 106660 41372 106724 41376
rect 106660 41316 106664 41372
rect 106664 41316 106720 41372
rect 106720 41316 106724 41372
rect 106660 41312 106724 41316
rect 106740 41372 106804 41376
rect 106740 41316 106744 41372
rect 106744 41316 106800 41372
rect 106800 41316 106804 41372
rect 106740 41312 106804 41316
rect 106820 41372 106884 41376
rect 106820 41316 106824 41372
rect 106824 41316 106880 41372
rect 106880 41316 106884 41372
rect 106820 41312 106884 41316
rect 106900 41372 106964 41376
rect 106900 41316 106904 41372
rect 106904 41316 106960 41372
rect 106960 41316 106964 41372
rect 106900 41312 106964 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 105924 40828 105988 40832
rect 105924 40772 105928 40828
rect 105928 40772 105984 40828
rect 105984 40772 105988 40828
rect 105924 40768 105988 40772
rect 106004 40828 106068 40832
rect 106004 40772 106008 40828
rect 106008 40772 106064 40828
rect 106064 40772 106068 40828
rect 106004 40768 106068 40772
rect 106084 40828 106148 40832
rect 106084 40772 106088 40828
rect 106088 40772 106144 40828
rect 106144 40772 106148 40828
rect 106084 40768 106148 40772
rect 106164 40828 106228 40832
rect 106164 40772 106168 40828
rect 106168 40772 106224 40828
rect 106224 40772 106228 40828
rect 106164 40768 106228 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 106660 40284 106724 40288
rect 106660 40228 106664 40284
rect 106664 40228 106720 40284
rect 106720 40228 106724 40284
rect 106660 40224 106724 40228
rect 106740 40284 106804 40288
rect 106740 40228 106744 40284
rect 106744 40228 106800 40284
rect 106800 40228 106804 40284
rect 106740 40224 106804 40228
rect 106820 40284 106884 40288
rect 106820 40228 106824 40284
rect 106824 40228 106880 40284
rect 106880 40228 106884 40284
rect 106820 40224 106884 40228
rect 106900 40284 106964 40288
rect 106900 40228 106904 40284
rect 106904 40228 106960 40284
rect 106960 40228 106964 40284
rect 106900 40224 106964 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 105924 39740 105988 39744
rect 105924 39684 105928 39740
rect 105928 39684 105984 39740
rect 105984 39684 105988 39740
rect 105924 39680 105988 39684
rect 106004 39740 106068 39744
rect 106004 39684 106008 39740
rect 106008 39684 106064 39740
rect 106064 39684 106068 39740
rect 106004 39680 106068 39684
rect 106084 39740 106148 39744
rect 106084 39684 106088 39740
rect 106088 39684 106144 39740
rect 106144 39684 106148 39740
rect 106084 39680 106148 39684
rect 106164 39740 106228 39744
rect 106164 39684 106168 39740
rect 106168 39684 106224 39740
rect 106224 39684 106228 39740
rect 106164 39680 106228 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 106660 39196 106724 39200
rect 106660 39140 106664 39196
rect 106664 39140 106720 39196
rect 106720 39140 106724 39196
rect 106660 39136 106724 39140
rect 106740 39196 106804 39200
rect 106740 39140 106744 39196
rect 106744 39140 106800 39196
rect 106800 39140 106804 39196
rect 106740 39136 106804 39140
rect 106820 39196 106884 39200
rect 106820 39140 106824 39196
rect 106824 39140 106880 39196
rect 106880 39140 106884 39196
rect 106820 39136 106884 39140
rect 106900 39196 106964 39200
rect 106900 39140 106904 39196
rect 106904 39140 106960 39196
rect 106960 39140 106964 39196
rect 106900 39136 106964 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 105924 38652 105988 38656
rect 105924 38596 105928 38652
rect 105928 38596 105984 38652
rect 105984 38596 105988 38652
rect 105924 38592 105988 38596
rect 106004 38652 106068 38656
rect 106004 38596 106008 38652
rect 106008 38596 106064 38652
rect 106064 38596 106068 38652
rect 106004 38592 106068 38596
rect 106084 38652 106148 38656
rect 106084 38596 106088 38652
rect 106088 38596 106144 38652
rect 106144 38596 106148 38652
rect 106084 38592 106148 38596
rect 106164 38652 106228 38656
rect 106164 38596 106168 38652
rect 106168 38596 106224 38652
rect 106224 38596 106228 38652
rect 106164 38592 106228 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 106660 38108 106724 38112
rect 106660 38052 106664 38108
rect 106664 38052 106720 38108
rect 106720 38052 106724 38108
rect 106660 38048 106724 38052
rect 106740 38108 106804 38112
rect 106740 38052 106744 38108
rect 106744 38052 106800 38108
rect 106800 38052 106804 38108
rect 106740 38048 106804 38052
rect 106820 38108 106884 38112
rect 106820 38052 106824 38108
rect 106824 38052 106880 38108
rect 106880 38052 106884 38108
rect 106820 38048 106884 38052
rect 106900 38108 106964 38112
rect 106900 38052 106904 38108
rect 106904 38052 106960 38108
rect 106960 38052 106964 38108
rect 106900 38048 106964 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 105924 37564 105988 37568
rect 105924 37508 105928 37564
rect 105928 37508 105984 37564
rect 105984 37508 105988 37564
rect 105924 37504 105988 37508
rect 106004 37564 106068 37568
rect 106004 37508 106008 37564
rect 106008 37508 106064 37564
rect 106064 37508 106068 37564
rect 106004 37504 106068 37508
rect 106084 37564 106148 37568
rect 106084 37508 106088 37564
rect 106088 37508 106144 37564
rect 106144 37508 106148 37564
rect 106084 37504 106148 37508
rect 106164 37564 106228 37568
rect 106164 37508 106168 37564
rect 106168 37508 106224 37564
rect 106224 37508 106228 37564
rect 106164 37504 106228 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 106660 37020 106724 37024
rect 106660 36964 106664 37020
rect 106664 36964 106720 37020
rect 106720 36964 106724 37020
rect 106660 36960 106724 36964
rect 106740 37020 106804 37024
rect 106740 36964 106744 37020
rect 106744 36964 106800 37020
rect 106800 36964 106804 37020
rect 106740 36960 106804 36964
rect 106820 37020 106884 37024
rect 106820 36964 106824 37020
rect 106824 36964 106880 37020
rect 106880 36964 106884 37020
rect 106820 36960 106884 36964
rect 106900 37020 106964 37024
rect 106900 36964 106904 37020
rect 106904 36964 106960 37020
rect 106960 36964 106964 37020
rect 106900 36960 106964 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 105924 36476 105988 36480
rect 105924 36420 105928 36476
rect 105928 36420 105984 36476
rect 105984 36420 105988 36476
rect 105924 36416 105988 36420
rect 106004 36476 106068 36480
rect 106004 36420 106008 36476
rect 106008 36420 106064 36476
rect 106064 36420 106068 36476
rect 106004 36416 106068 36420
rect 106084 36476 106148 36480
rect 106084 36420 106088 36476
rect 106088 36420 106144 36476
rect 106144 36420 106148 36476
rect 106084 36416 106148 36420
rect 106164 36476 106228 36480
rect 106164 36420 106168 36476
rect 106168 36420 106224 36476
rect 106224 36420 106228 36476
rect 106164 36416 106228 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 106660 35932 106724 35936
rect 106660 35876 106664 35932
rect 106664 35876 106720 35932
rect 106720 35876 106724 35932
rect 106660 35872 106724 35876
rect 106740 35932 106804 35936
rect 106740 35876 106744 35932
rect 106744 35876 106800 35932
rect 106800 35876 106804 35932
rect 106740 35872 106804 35876
rect 106820 35932 106884 35936
rect 106820 35876 106824 35932
rect 106824 35876 106880 35932
rect 106880 35876 106884 35932
rect 106820 35872 106884 35876
rect 106900 35932 106964 35936
rect 106900 35876 106904 35932
rect 106904 35876 106960 35932
rect 106960 35876 106964 35932
rect 106900 35872 106964 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 105924 35388 105988 35392
rect 105924 35332 105928 35388
rect 105928 35332 105984 35388
rect 105984 35332 105988 35388
rect 105924 35328 105988 35332
rect 106004 35388 106068 35392
rect 106004 35332 106008 35388
rect 106008 35332 106064 35388
rect 106064 35332 106068 35388
rect 106004 35328 106068 35332
rect 106084 35388 106148 35392
rect 106084 35332 106088 35388
rect 106088 35332 106144 35388
rect 106144 35332 106148 35388
rect 106084 35328 106148 35332
rect 106164 35388 106228 35392
rect 106164 35332 106168 35388
rect 106168 35332 106224 35388
rect 106224 35332 106228 35388
rect 106164 35328 106228 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 106660 34844 106724 34848
rect 106660 34788 106664 34844
rect 106664 34788 106720 34844
rect 106720 34788 106724 34844
rect 106660 34784 106724 34788
rect 106740 34844 106804 34848
rect 106740 34788 106744 34844
rect 106744 34788 106800 34844
rect 106800 34788 106804 34844
rect 106740 34784 106804 34788
rect 106820 34844 106884 34848
rect 106820 34788 106824 34844
rect 106824 34788 106880 34844
rect 106880 34788 106884 34844
rect 106820 34784 106884 34788
rect 106900 34844 106964 34848
rect 106900 34788 106904 34844
rect 106904 34788 106960 34844
rect 106960 34788 106964 34844
rect 106900 34784 106964 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 105924 34300 105988 34304
rect 105924 34244 105928 34300
rect 105928 34244 105984 34300
rect 105984 34244 105988 34300
rect 105924 34240 105988 34244
rect 106004 34300 106068 34304
rect 106004 34244 106008 34300
rect 106008 34244 106064 34300
rect 106064 34244 106068 34300
rect 106004 34240 106068 34244
rect 106084 34300 106148 34304
rect 106084 34244 106088 34300
rect 106088 34244 106144 34300
rect 106144 34244 106148 34300
rect 106084 34240 106148 34244
rect 106164 34300 106228 34304
rect 106164 34244 106168 34300
rect 106168 34244 106224 34300
rect 106224 34244 106228 34300
rect 106164 34240 106228 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 106660 33756 106724 33760
rect 106660 33700 106664 33756
rect 106664 33700 106720 33756
rect 106720 33700 106724 33756
rect 106660 33696 106724 33700
rect 106740 33756 106804 33760
rect 106740 33700 106744 33756
rect 106744 33700 106800 33756
rect 106800 33700 106804 33756
rect 106740 33696 106804 33700
rect 106820 33756 106884 33760
rect 106820 33700 106824 33756
rect 106824 33700 106880 33756
rect 106880 33700 106884 33756
rect 106820 33696 106884 33700
rect 106900 33756 106964 33760
rect 106900 33700 106904 33756
rect 106904 33700 106960 33756
rect 106960 33700 106964 33756
rect 106900 33696 106964 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 105924 33212 105988 33216
rect 105924 33156 105928 33212
rect 105928 33156 105984 33212
rect 105984 33156 105988 33212
rect 105924 33152 105988 33156
rect 106004 33212 106068 33216
rect 106004 33156 106008 33212
rect 106008 33156 106064 33212
rect 106064 33156 106068 33212
rect 106004 33152 106068 33156
rect 106084 33212 106148 33216
rect 106084 33156 106088 33212
rect 106088 33156 106144 33212
rect 106144 33156 106148 33212
rect 106084 33152 106148 33156
rect 106164 33212 106228 33216
rect 106164 33156 106168 33212
rect 106168 33156 106224 33212
rect 106224 33156 106228 33212
rect 106164 33152 106228 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 106660 32668 106724 32672
rect 106660 32612 106664 32668
rect 106664 32612 106720 32668
rect 106720 32612 106724 32668
rect 106660 32608 106724 32612
rect 106740 32668 106804 32672
rect 106740 32612 106744 32668
rect 106744 32612 106800 32668
rect 106800 32612 106804 32668
rect 106740 32608 106804 32612
rect 106820 32668 106884 32672
rect 106820 32612 106824 32668
rect 106824 32612 106880 32668
rect 106880 32612 106884 32668
rect 106820 32608 106884 32612
rect 106900 32668 106964 32672
rect 106900 32612 106904 32668
rect 106904 32612 106960 32668
rect 106960 32612 106964 32668
rect 106900 32608 106964 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 105924 32124 105988 32128
rect 105924 32068 105928 32124
rect 105928 32068 105984 32124
rect 105984 32068 105988 32124
rect 105924 32064 105988 32068
rect 106004 32124 106068 32128
rect 106004 32068 106008 32124
rect 106008 32068 106064 32124
rect 106064 32068 106068 32124
rect 106004 32064 106068 32068
rect 106084 32124 106148 32128
rect 106084 32068 106088 32124
rect 106088 32068 106144 32124
rect 106144 32068 106148 32124
rect 106084 32064 106148 32068
rect 106164 32124 106228 32128
rect 106164 32068 106168 32124
rect 106168 32068 106224 32124
rect 106224 32068 106228 32124
rect 106164 32064 106228 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 106660 31580 106724 31584
rect 106660 31524 106664 31580
rect 106664 31524 106720 31580
rect 106720 31524 106724 31580
rect 106660 31520 106724 31524
rect 106740 31580 106804 31584
rect 106740 31524 106744 31580
rect 106744 31524 106800 31580
rect 106800 31524 106804 31580
rect 106740 31520 106804 31524
rect 106820 31580 106884 31584
rect 106820 31524 106824 31580
rect 106824 31524 106880 31580
rect 106880 31524 106884 31580
rect 106820 31520 106884 31524
rect 106900 31580 106964 31584
rect 106900 31524 106904 31580
rect 106904 31524 106960 31580
rect 106960 31524 106964 31580
rect 106900 31520 106964 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 105924 31036 105988 31040
rect 105924 30980 105928 31036
rect 105928 30980 105984 31036
rect 105984 30980 105988 31036
rect 105924 30976 105988 30980
rect 106004 31036 106068 31040
rect 106004 30980 106008 31036
rect 106008 30980 106064 31036
rect 106064 30980 106068 31036
rect 106004 30976 106068 30980
rect 106084 31036 106148 31040
rect 106084 30980 106088 31036
rect 106088 30980 106144 31036
rect 106144 30980 106148 31036
rect 106084 30976 106148 30980
rect 106164 31036 106228 31040
rect 106164 30980 106168 31036
rect 106168 30980 106224 31036
rect 106224 30980 106228 31036
rect 106164 30976 106228 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 106660 30492 106724 30496
rect 106660 30436 106664 30492
rect 106664 30436 106720 30492
rect 106720 30436 106724 30492
rect 106660 30432 106724 30436
rect 106740 30492 106804 30496
rect 106740 30436 106744 30492
rect 106744 30436 106800 30492
rect 106800 30436 106804 30492
rect 106740 30432 106804 30436
rect 106820 30492 106884 30496
rect 106820 30436 106824 30492
rect 106824 30436 106880 30492
rect 106880 30436 106884 30492
rect 106820 30432 106884 30436
rect 106900 30492 106964 30496
rect 106900 30436 106904 30492
rect 106904 30436 106960 30492
rect 106960 30436 106964 30492
rect 106900 30432 106964 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 105924 29948 105988 29952
rect 105924 29892 105928 29948
rect 105928 29892 105984 29948
rect 105984 29892 105988 29948
rect 105924 29888 105988 29892
rect 106004 29948 106068 29952
rect 106004 29892 106008 29948
rect 106008 29892 106064 29948
rect 106064 29892 106068 29948
rect 106004 29888 106068 29892
rect 106084 29948 106148 29952
rect 106084 29892 106088 29948
rect 106088 29892 106144 29948
rect 106144 29892 106148 29948
rect 106084 29888 106148 29892
rect 106164 29948 106228 29952
rect 106164 29892 106168 29948
rect 106168 29892 106224 29948
rect 106224 29892 106228 29948
rect 106164 29888 106228 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 106660 29404 106724 29408
rect 106660 29348 106664 29404
rect 106664 29348 106720 29404
rect 106720 29348 106724 29404
rect 106660 29344 106724 29348
rect 106740 29404 106804 29408
rect 106740 29348 106744 29404
rect 106744 29348 106800 29404
rect 106800 29348 106804 29404
rect 106740 29344 106804 29348
rect 106820 29404 106884 29408
rect 106820 29348 106824 29404
rect 106824 29348 106880 29404
rect 106880 29348 106884 29404
rect 106820 29344 106884 29348
rect 106900 29404 106964 29408
rect 106900 29348 106904 29404
rect 106904 29348 106960 29404
rect 106960 29348 106964 29404
rect 106900 29344 106964 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 105924 28860 105988 28864
rect 105924 28804 105928 28860
rect 105928 28804 105984 28860
rect 105984 28804 105988 28860
rect 105924 28800 105988 28804
rect 106004 28860 106068 28864
rect 106004 28804 106008 28860
rect 106008 28804 106064 28860
rect 106064 28804 106068 28860
rect 106004 28800 106068 28804
rect 106084 28860 106148 28864
rect 106084 28804 106088 28860
rect 106088 28804 106144 28860
rect 106144 28804 106148 28860
rect 106084 28800 106148 28804
rect 106164 28860 106228 28864
rect 106164 28804 106168 28860
rect 106168 28804 106224 28860
rect 106224 28804 106228 28860
rect 106164 28800 106228 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 106660 28316 106724 28320
rect 106660 28260 106664 28316
rect 106664 28260 106720 28316
rect 106720 28260 106724 28316
rect 106660 28256 106724 28260
rect 106740 28316 106804 28320
rect 106740 28260 106744 28316
rect 106744 28260 106800 28316
rect 106800 28260 106804 28316
rect 106740 28256 106804 28260
rect 106820 28316 106884 28320
rect 106820 28260 106824 28316
rect 106824 28260 106880 28316
rect 106880 28260 106884 28316
rect 106820 28256 106884 28260
rect 106900 28316 106964 28320
rect 106900 28260 106904 28316
rect 106904 28260 106960 28316
rect 106960 28260 106964 28316
rect 106900 28256 106964 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 105924 27772 105988 27776
rect 105924 27716 105928 27772
rect 105928 27716 105984 27772
rect 105984 27716 105988 27772
rect 105924 27712 105988 27716
rect 106004 27772 106068 27776
rect 106004 27716 106008 27772
rect 106008 27716 106064 27772
rect 106064 27716 106068 27772
rect 106004 27712 106068 27716
rect 106084 27772 106148 27776
rect 106084 27716 106088 27772
rect 106088 27716 106144 27772
rect 106144 27716 106148 27772
rect 106084 27712 106148 27716
rect 106164 27772 106228 27776
rect 106164 27716 106168 27772
rect 106168 27716 106224 27772
rect 106224 27716 106228 27772
rect 106164 27712 106228 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 106660 27228 106724 27232
rect 106660 27172 106664 27228
rect 106664 27172 106720 27228
rect 106720 27172 106724 27228
rect 106660 27168 106724 27172
rect 106740 27228 106804 27232
rect 106740 27172 106744 27228
rect 106744 27172 106800 27228
rect 106800 27172 106804 27228
rect 106740 27168 106804 27172
rect 106820 27228 106884 27232
rect 106820 27172 106824 27228
rect 106824 27172 106880 27228
rect 106880 27172 106884 27228
rect 106820 27168 106884 27172
rect 106900 27228 106964 27232
rect 106900 27172 106904 27228
rect 106904 27172 106960 27228
rect 106960 27172 106964 27228
rect 106900 27168 106964 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 105924 26684 105988 26688
rect 105924 26628 105928 26684
rect 105928 26628 105984 26684
rect 105984 26628 105988 26684
rect 105924 26624 105988 26628
rect 106004 26684 106068 26688
rect 106004 26628 106008 26684
rect 106008 26628 106064 26684
rect 106064 26628 106068 26684
rect 106004 26624 106068 26628
rect 106084 26684 106148 26688
rect 106084 26628 106088 26684
rect 106088 26628 106144 26684
rect 106144 26628 106148 26684
rect 106084 26624 106148 26628
rect 106164 26684 106228 26688
rect 106164 26628 106168 26684
rect 106168 26628 106224 26684
rect 106224 26628 106228 26684
rect 106164 26624 106228 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 106660 26140 106724 26144
rect 106660 26084 106664 26140
rect 106664 26084 106720 26140
rect 106720 26084 106724 26140
rect 106660 26080 106724 26084
rect 106740 26140 106804 26144
rect 106740 26084 106744 26140
rect 106744 26084 106800 26140
rect 106800 26084 106804 26140
rect 106740 26080 106804 26084
rect 106820 26140 106884 26144
rect 106820 26084 106824 26140
rect 106824 26084 106880 26140
rect 106880 26084 106884 26140
rect 106820 26080 106884 26084
rect 106900 26140 106964 26144
rect 106900 26084 106904 26140
rect 106904 26084 106960 26140
rect 106960 26084 106964 26140
rect 106900 26080 106964 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 105924 25596 105988 25600
rect 105924 25540 105928 25596
rect 105928 25540 105984 25596
rect 105984 25540 105988 25596
rect 105924 25536 105988 25540
rect 106004 25596 106068 25600
rect 106004 25540 106008 25596
rect 106008 25540 106064 25596
rect 106064 25540 106068 25596
rect 106004 25536 106068 25540
rect 106084 25596 106148 25600
rect 106084 25540 106088 25596
rect 106088 25540 106144 25596
rect 106144 25540 106148 25596
rect 106084 25536 106148 25540
rect 106164 25596 106228 25600
rect 106164 25540 106168 25596
rect 106168 25540 106224 25596
rect 106224 25540 106228 25596
rect 106164 25536 106228 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 106660 25052 106724 25056
rect 106660 24996 106664 25052
rect 106664 24996 106720 25052
rect 106720 24996 106724 25052
rect 106660 24992 106724 24996
rect 106740 25052 106804 25056
rect 106740 24996 106744 25052
rect 106744 24996 106800 25052
rect 106800 24996 106804 25052
rect 106740 24992 106804 24996
rect 106820 25052 106884 25056
rect 106820 24996 106824 25052
rect 106824 24996 106880 25052
rect 106880 24996 106884 25052
rect 106820 24992 106884 24996
rect 106900 25052 106964 25056
rect 106900 24996 106904 25052
rect 106904 24996 106960 25052
rect 106960 24996 106964 25052
rect 106900 24992 106964 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 105924 24508 105988 24512
rect 105924 24452 105928 24508
rect 105928 24452 105984 24508
rect 105984 24452 105988 24508
rect 105924 24448 105988 24452
rect 106004 24508 106068 24512
rect 106004 24452 106008 24508
rect 106008 24452 106064 24508
rect 106064 24452 106068 24508
rect 106004 24448 106068 24452
rect 106084 24508 106148 24512
rect 106084 24452 106088 24508
rect 106088 24452 106144 24508
rect 106144 24452 106148 24508
rect 106084 24448 106148 24452
rect 106164 24508 106228 24512
rect 106164 24452 106168 24508
rect 106168 24452 106224 24508
rect 106224 24452 106228 24508
rect 106164 24448 106228 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 106660 23964 106724 23968
rect 106660 23908 106664 23964
rect 106664 23908 106720 23964
rect 106720 23908 106724 23964
rect 106660 23904 106724 23908
rect 106740 23964 106804 23968
rect 106740 23908 106744 23964
rect 106744 23908 106800 23964
rect 106800 23908 106804 23964
rect 106740 23904 106804 23908
rect 106820 23964 106884 23968
rect 106820 23908 106824 23964
rect 106824 23908 106880 23964
rect 106880 23908 106884 23964
rect 106820 23904 106884 23908
rect 106900 23964 106964 23968
rect 106900 23908 106904 23964
rect 106904 23908 106960 23964
rect 106960 23908 106964 23964
rect 106900 23904 106964 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 105924 23420 105988 23424
rect 105924 23364 105928 23420
rect 105928 23364 105984 23420
rect 105984 23364 105988 23420
rect 105924 23360 105988 23364
rect 106004 23420 106068 23424
rect 106004 23364 106008 23420
rect 106008 23364 106064 23420
rect 106064 23364 106068 23420
rect 106004 23360 106068 23364
rect 106084 23420 106148 23424
rect 106084 23364 106088 23420
rect 106088 23364 106144 23420
rect 106144 23364 106148 23420
rect 106084 23360 106148 23364
rect 106164 23420 106228 23424
rect 106164 23364 106168 23420
rect 106168 23364 106224 23420
rect 106224 23364 106228 23420
rect 106164 23360 106228 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 106660 22876 106724 22880
rect 106660 22820 106664 22876
rect 106664 22820 106720 22876
rect 106720 22820 106724 22876
rect 106660 22816 106724 22820
rect 106740 22876 106804 22880
rect 106740 22820 106744 22876
rect 106744 22820 106800 22876
rect 106800 22820 106804 22876
rect 106740 22816 106804 22820
rect 106820 22876 106884 22880
rect 106820 22820 106824 22876
rect 106824 22820 106880 22876
rect 106880 22820 106884 22876
rect 106820 22816 106884 22820
rect 106900 22876 106964 22880
rect 106900 22820 106904 22876
rect 106904 22820 106960 22876
rect 106960 22820 106964 22876
rect 106900 22816 106964 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 105924 22332 105988 22336
rect 105924 22276 105928 22332
rect 105928 22276 105984 22332
rect 105984 22276 105988 22332
rect 105924 22272 105988 22276
rect 106004 22332 106068 22336
rect 106004 22276 106008 22332
rect 106008 22276 106064 22332
rect 106064 22276 106068 22332
rect 106004 22272 106068 22276
rect 106084 22332 106148 22336
rect 106084 22276 106088 22332
rect 106088 22276 106144 22332
rect 106144 22276 106148 22332
rect 106084 22272 106148 22276
rect 106164 22332 106228 22336
rect 106164 22276 106168 22332
rect 106168 22276 106224 22332
rect 106224 22276 106228 22332
rect 106164 22272 106228 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 106660 21788 106724 21792
rect 106660 21732 106664 21788
rect 106664 21732 106720 21788
rect 106720 21732 106724 21788
rect 106660 21728 106724 21732
rect 106740 21788 106804 21792
rect 106740 21732 106744 21788
rect 106744 21732 106800 21788
rect 106800 21732 106804 21788
rect 106740 21728 106804 21732
rect 106820 21788 106884 21792
rect 106820 21732 106824 21788
rect 106824 21732 106880 21788
rect 106880 21732 106884 21788
rect 106820 21728 106884 21732
rect 106900 21788 106964 21792
rect 106900 21732 106904 21788
rect 106904 21732 106960 21788
rect 106960 21732 106964 21788
rect 106900 21728 106964 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 105924 21244 105988 21248
rect 105924 21188 105928 21244
rect 105928 21188 105984 21244
rect 105984 21188 105988 21244
rect 105924 21184 105988 21188
rect 106004 21244 106068 21248
rect 106004 21188 106008 21244
rect 106008 21188 106064 21244
rect 106064 21188 106068 21244
rect 106004 21184 106068 21188
rect 106084 21244 106148 21248
rect 106084 21188 106088 21244
rect 106088 21188 106144 21244
rect 106144 21188 106148 21244
rect 106084 21184 106148 21188
rect 106164 21244 106228 21248
rect 106164 21188 106168 21244
rect 106168 21188 106224 21244
rect 106224 21188 106228 21244
rect 106164 21184 106228 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 106660 20700 106724 20704
rect 106660 20644 106664 20700
rect 106664 20644 106720 20700
rect 106720 20644 106724 20700
rect 106660 20640 106724 20644
rect 106740 20700 106804 20704
rect 106740 20644 106744 20700
rect 106744 20644 106800 20700
rect 106800 20644 106804 20700
rect 106740 20640 106804 20644
rect 106820 20700 106884 20704
rect 106820 20644 106824 20700
rect 106824 20644 106880 20700
rect 106880 20644 106884 20700
rect 106820 20640 106884 20644
rect 106900 20700 106964 20704
rect 106900 20644 106904 20700
rect 106904 20644 106960 20700
rect 106960 20644 106964 20700
rect 106900 20640 106964 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 105924 20156 105988 20160
rect 105924 20100 105928 20156
rect 105928 20100 105984 20156
rect 105984 20100 105988 20156
rect 105924 20096 105988 20100
rect 106004 20156 106068 20160
rect 106004 20100 106008 20156
rect 106008 20100 106064 20156
rect 106064 20100 106068 20156
rect 106004 20096 106068 20100
rect 106084 20156 106148 20160
rect 106084 20100 106088 20156
rect 106088 20100 106144 20156
rect 106144 20100 106148 20156
rect 106084 20096 106148 20100
rect 106164 20156 106228 20160
rect 106164 20100 106168 20156
rect 106168 20100 106224 20156
rect 106224 20100 106228 20156
rect 106164 20096 106228 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 106660 19612 106724 19616
rect 106660 19556 106664 19612
rect 106664 19556 106720 19612
rect 106720 19556 106724 19612
rect 106660 19552 106724 19556
rect 106740 19612 106804 19616
rect 106740 19556 106744 19612
rect 106744 19556 106800 19612
rect 106800 19556 106804 19612
rect 106740 19552 106804 19556
rect 106820 19612 106884 19616
rect 106820 19556 106824 19612
rect 106824 19556 106880 19612
rect 106880 19556 106884 19612
rect 106820 19552 106884 19556
rect 106900 19612 106964 19616
rect 106900 19556 106904 19612
rect 106904 19556 106960 19612
rect 106960 19556 106964 19612
rect 106900 19552 106964 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 105924 19068 105988 19072
rect 105924 19012 105928 19068
rect 105928 19012 105984 19068
rect 105984 19012 105988 19068
rect 105924 19008 105988 19012
rect 106004 19068 106068 19072
rect 106004 19012 106008 19068
rect 106008 19012 106064 19068
rect 106064 19012 106068 19068
rect 106004 19008 106068 19012
rect 106084 19068 106148 19072
rect 106084 19012 106088 19068
rect 106088 19012 106144 19068
rect 106144 19012 106148 19068
rect 106084 19008 106148 19012
rect 106164 19068 106228 19072
rect 106164 19012 106168 19068
rect 106168 19012 106224 19068
rect 106224 19012 106228 19068
rect 106164 19008 106228 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 106660 18524 106724 18528
rect 106660 18468 106664 18524
rect 106664 18468 106720 18524
rect 106720 18468 106724 18524
rect 106660 18464 106724 18468
rect 106740 18524 106804 18528
rect 106740 18468 106744 18524
rect 106744 18468 106800 18524
rect 106800 18468 106804 18524
rect 106740 18464 106804 18468
rect 106820 18524 106884 18528
rect 106820 18468 106824 18524
rect 106824 18468 106880 18524
rect 106880 18468 106884 18524
rect 106820 18464 106884 18468
rect 106900 18524 106964 18528
rect 106900 18468 106904 18524
rect 106904 18468 106960 18524
rect 106960 18468 106964 18524
rect 106900 18464 106964 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 105924 17980 105988 17984
rect 105924 17924 105928 17980
rect 105928 17924 105984 17980
rect 105984 17924 105988 17980
rect 105924 17920 105988 17924
rect 106004 17980 106068 17984
rect 106004 17924 106008 17980
rect 106008 17924 106064 17980
rect 106064 17924 106068 17980
rect 106004 17920 106068 17924
rect 106084 17980 106148 17984
rect 106084 17924 106088 17980
rect 106088 17924 106144 17980
rect 106144 17924 106148 17980
rect 106084 17920 106148 17924
rect 106164 17980 106228 17984
rect 106164 17924 106168 17980
rect 106168 17924 106224 17980
rect 106224 17924 106228 17980
rect 106164 17920 106228 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 106660 17436 106724 17440
rect 106660 17380 106664 17436
rect 106664 17380 106720 17436
rect 106720 17380 106724 17436
rect 106660 17376 106724 17380
rect 106740 17436 106804 17440
rect 106740 17380 106744 17436
rect 106744 17380 106800 17436
rect 106800 17380 106804 17436
rect 106740 17376 106804 17380
rect 106820 17436 106884 17440
rect 106820 17380 106824 17436
rect 106824 17380 106880 17436
rect 106880 17380 106884 17436
rect 106820 17376 106884 17380
rect 106900 17436 106964 17440
rect 106900 17380 106904 17436
rect 106904 17380 106960 17436
rect 106960 17380 106964 17436
rect 106900 17376 106964 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 105924 16892 105988 16896
rect 105924 16836 105928 16892
rect 105928 16836 105984 16892
rect 105984 16836 105988 16892
rect 105924 16832 105988 16836
rect 106004 16892 106068 16896
rect 106004 16836 106008 16892
rect 106008 16836 106064 16892
rect 106064 16836 106068 16892
rect 106004 16832 106068 16836
rect 106084 16892 106148 16896
rect 106084 16836 106088 16892
rect 106088 16836 106144 16892
rect 106144 16836 106148 16892
rect 106084 16832 106148 16836
rect 106164 16892 106228 16896
rect 106164 16836 106168 16892
rect 106168 16836 106224 16892
rect 106224 16836 106228 16892
rect 106164 16832 106228 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 106660 16348 106724 16352
rect 106660 16292 106664 16348
rect 106664 16292 106720 16348
rect 106720 16292 106724 16348
rect 106660 16288 106724 16292
rect 106740 16348 106804 16352
rect 106740 16292 106744 16348
rect 106744 16292 106800 16348
rect 106800 16292 106804 16348
rect 106740 16288 106804 16292
rect 106820 16348 106884 16352
rect 106820 16292 106824 16348
rect 106824 16292 106880 16348
rect 106880 16292 106884 16348
rect 106820 16288 106884 16292
rect 106900 16348 106964 16352
rect 106900 16292 106904 16348
rect 106904 16292 106960 16348
rect 106960 16292 106964 16348
rect 106900 16288 106964 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 105924 15804 105988 15808
rect 105924 15748 105928 15804
rect 105928 15748 105984 15804
rect 105984 15748 105988 15804
rect 105924 15744 105988 15748
rect 106004 15804 106068 15808
rect 106004 15748 106008 15804
rect 106008 15748 106064 15804
rect 106064 15748 106068 15804
rect 106004 15744 106068 15748
rect 106084 15804 106148 15808
rect 106084 15748 106088 15804
rect 106088 15748 106144 15804
rect 106144 15748 106148 15804
rect 106084 15744 106148 15748
rect 106164 15804 106228 15808
rect 106164 15748 106168 15804
rect 106168 15748 106224 15804
rect 106224 15748 106228 15804
rect 106164 15744 106228 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 106660 15260 106724 15264
rect 106660 15204 106664 15260
rect 106664 15204 106720 15260
rect 106720 15204 106724 15260
rect 106660 15200 106724 15204
rect 106740 15260 106804 15264
rect 106740 15204 106744 15260
rect 106744 15204 106800 15260
rect 106800 15204 106804 15260
rect 106740 15200 106804 15204
rect 106820 15260 106884 15264
rect 106820 15204 106824 15260
rect 106824 15204 106880 15260
rect 106880 15204 106884 15260
rect 106820 15200 106884 15204
rect 106900 15260 106964 15264
rect 106900 15204 106904 15260
rect 106904 15204 106960 15260
rect 106960 15204 106964 15260
rect 106900 15200 106964 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 105924 14716 105988 14720
rect 105924 14660 105928 14716
rect 105928 14660 105984 14716
rect 105984 14660 105988 14716
rect 105924 14656 105988 14660
rect 106004 14716 106068 14720
rect 106004 14660 106008 14716
rect 106008 14660 106064 14716
rect 106064 14660 106068 14716
rect 106004 14656 106068 14660
rect 106084 14716 106148 14720
rect 106084 14660 106088 14716
rect 106088 14660 106144 14716
rect 106144 14660 106148 14716
rect 106084 14656 106148 14660
rect 106164 14716 106228 14720
rect 106164 14660 106168 14716
rect 106168 14660 106224 14716
rect 106224 14660 106228 14716
rect 106164 14656 106228 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 106660 14172 106724 14176
rect 106660 14116 106664 14172
rect 106664 14116 106720 14172
rect 106720 14116 106724 14172
rect 106660 14112 106724 14116
rect 106740 14172 106804 14176
rect 106740 14116 106744 14172
rect 106744 14116 106800 14172
rect 106800 14116 106804 14172
rect 106740 14112 106804 14116
rect 106820 14172 106884 14176
rect 106820 14116 106824 14172
rect 106824 14116 106880 14172
rect 106880 14116 106884 14172
rect 106820 14112 106884 14116
rect 106900 14172 106964 14176
rect 106900 14116 106904 14172
rect 106904 14116 106960 14172
rect 106960 14116 106964 14172
rect 106900 14112 106964 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 105924 13628 105988 13632
rect 105924 13572 105928 13628
rect 105928 13572 105984 13628
rect 105984 13572 105988 13628
rect 105924 13568 105988 13572
rect 106004 13628 106068 13632
rect 106004 13572 106008 13628
rect 106008 13572 106064 13628
rect 106064 13572 106068 13628
rect 106004 13568 106068 13572
rect 106084 13628 106148 13632
rect 106084 13572 106088 13628
rect 106088 13572 106144 13628
rect 106144 13572 106148 13628
rect 106084 13568 106148 13572
rect 106164 13628 106228 13632
rect 106164 13572 106168 13628
rect 106168 13572 106224 13628
rect 106224 13572 106228 13628
rect 106164 13568 106228 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 106660 13084 106724 13088
rect 106660 13028 106664 13084
rect 106664 13028 106720 13084
rect 106720 13028 106724 13084
rect 106660 13024 106724 13028
rect 106740 13084 106804 13088
rect 106740 13028 106744 13084
rect 106744 13028 106800 13084
rect 106800 13028 106804 13084
rect 106740 13024 106804 13028
rect 106820 13084 106884 13088
rect 106820 13028 106824 13084
rect 106824 13028 106880 13084
rect 106880 13028 106884 13084
rect 106820 13024 106884 13028
rect 106900 13084 106964 13088
rect 106900 13028 106904 13084
rect 106904 13028 106960 13084
rect 106960 13028 106964 13084
rect 106900 13024 106964 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 105924 12540 105988 12544
rect 105924 12484 105928 12540
rect 105928 12484 105984 12540
rect 105984 12484 105988 12540
rect 105924 12480 105988 12484
rect 106004 12540 106068 12544
rect 106004 12484 106008 12540
rect 106008 12484 106064 12540
rect 106064 12484 106068 12540
rect 106004 12480 106068 12484
rect 106084 12540 106148 12544
rect 106084 12484 106088 12540
rect 106088 12484 106144 12540
rect 106144 12484 106148 12540
rect 106084 12480 106148 12484
rect 106164 12540 106228 12544
rect 106164 12484 106168 12540
rect 106168 12484 106224 12540
rect 106224 12484 106228 12540
rect 106164 12480 106228 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 106660 11996 106724 12000
rect 106660 11940 106664 11996
rect 106664 11940 106720 11996
rect 106720 11940 106724 11996
rect 106660 11936 106724 11940
rect 106740 11996 106804 12000
rect 106740 11940 106744 11996
rect 106744 11940 106800 11996
rect 106800 11940 106804 11996
rect 106740 11936 106804 11940
rect 106820 11996 106884 12000
rect 106820 11940 106824 11996
rect 106824 11940 106880 11996
rect 106880 11940 106884 11996
rect 106820 11936 106884 11940
rect 106900 11996 106964 12000
rect 106900 11940 106904 11996
rect 106904 11940 106960 11996
rect 106960 11940 106964 11996
rect 106900 11936 106964 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 105924 11452 105988 11456
rect 105924 11396 105928 11452
rect 105928 11396 105984 11452
rect 105984 11396 105988 11452
rect 105924 11392 105988 11396
rect 106004 11452 106068 11456
rect 106004 11396 106008 11452
rect 106008 11396 106064 11452
rect 106064 11396 106068 11452
rect 106004 11392 106068 11396
rect 106084 11452 106148 11456
rect 106084 11396 106088 11452
rect 106088 11396 106144 11452
rect 106144 11396 106148 11452
rect 106084 11392 106148 11396
rect 106164 11452 106228 11456
rect 106164 11396 106168 11452
rect 106168 11396 106224 11452
rect 106224 11396 106228 11452
rect 106164 11392 106228 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 106660 10908 106724 10912
rect 106660 10852 106664 10908
rect 106664 10852 106720 10908
rect 106720 10852 106724 10908
rect 106660 10848 106724 10852
rect 106740 10908 106804 10912
rect 106740 10852 106744 10908
rect 106744 10852 106800 10908
rect 106800 10852 106804 10908
rect 106740 10848 106804 10852
rect 106820 10908 106884 10912
rect 106820 10852 106824 10908
rect 106824 10852 106880 10908
rect 106880 10852 106884 10908
rect 106820 10848 106884 10852
rect 106900 10908 106964 10912
rect 106900 10852 106904 10908
rect 106904 10852 106960 10908
rect 106960 10852 106964 10908
rect 106900 10848 106964 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 105924 10364 105988 10368
rect 105924 10308 105928 10364
rect 105928 10308 105984 10364
rect 105984 10308 105988 10364
rect 105924 10304 105988 10308
rect 106004 10364 106068 10368
rect 106004 10308 106008 10364
rect 106008 10308 106064 10364
rect 106064 10308 106068 10364
rect 106004 10304 106068 10308
rect 106084 10364 106148 10368
rect 106084 10308 106088 10364
rect 106088 10308 106144 10364
rect 106144 10308 106148 10364
rect 106084 10304 106148 10308
rect 106164 10364 106228 10368
rect 106164 10308 106168 10364
rect 106168 10308 106224 10364
rect 106224 10308 106228 10364
rect 106164 10304 106228 10308
rect 16058 9888 16122 9892
rect 16058 9832 16118 9888
rect 16118 9832 16122 9888
rect 16058 9828 16122 9832
rect 90527 9828 90591 9892
rect 90956 9828 91020 9892
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 106660 9820 106724 9824
rect 106660 9764 106664 9820
rect 106664 9764 106720 9820
rect 106720 9764 106724 9820
rect 106660 9760 106724 9764
rect 106740 9820 106804 9824
rect 106740 9764 106744 9820
rect 106744 9764 106800 9820
rect 106800 9764 106804 9820
rect 106740 9760 106804 9764
rect 106820 9820 106884 9824
rect 106820 9764 106824 9820
rect 106824 9764 106880 9820
rect 106880 9764 106884 9820
rect 106820 9760 106884 9764
rect 106900 9820 106964 9824
rect 106900 9764 106904 9820
rect 106904 9764 106960 9820
rect 106960 9764 106964 9820
rect 106900 9760 106964 9764
rect 90680 9752 90744 9756
rect 90680 9696 90730 9752
rect 90730 9696 90744 9752
rect 90680 9692 90744 9696
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 105924 9276 105988 9280
rect 105924 9220 105928 9276
rect 105928 9220 105984 9276
rect 105984 9220 105988 9276
rect 105924 9216 105988 9220
rect 106004 9276 106068 9280
rect 106004 9220 106008 9276
rect 106008 9220 106064 9276
rect 106064 9220 106068 9276
rect 106004 9216 106068 9220
rect 106084 9276 106148 9280
rect 106084 9220 106088 9276
rect 106088 9220 106144 9276
rect 106144 9220 106148 9276
rect 106084 9216 106148 9220
rect 106164 9276 106228 9280
rect 106164 9220 106168 9276
rect 106168 9220 106224 9276
rect 106224 9220 106228 9276
rect 106164 9216 106228 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 106660 8732 106724 8736
rect 106660 8676 106664 8732
rect 106664 8676 106720 8732
rect 106720 8676 106724 8732
rect 106660 8672 106724 8676
rect 106740 8732 106804 8736
rect 106740 8676 106744 8732
rect 106744 8676 106800 8732
rect 106800 8676 106804 8732
rect 106740 8672 106804 8676
rect 106820 8732 106884 8736
rect 106820 8676 106824 8732
rect 106824 8676 106880 8732
rect 106880 8676 106884 8732
rect 106820 8672 106884 8676
rect 106900 8732 106964 8736
rect 106900 8676 106904 8732
rect 106904 8676 106960 8732
rect 106960 8676 106964 8732
rect 106900 8672 106964 8676
rect 23428 8256 23492 8260
rect 23428 8200 23478 8256
rect 23478 8200 23492 8256
rect 23428 8196 23492 8200
rect 24716 8256 24780 8260
rect 24716 8200 24766 8256
rect 24766 8200 24780 8256
rect 24716 8196 24780 8200
rect 25820 8256 25884 8260
rect 25820 8200 25870 8256
rect 25870 8200 25884 8256
rect 25820 8196 25884 8200
rect 26924 8196 26988 8260
rect 28212 8196 28276 8260
rect 29316 8256 29380 8260
rect 29316 8200 29330 8256
rect 29330 8200 29380 8256
rect 29316 8196 29380 8200
rect 30420 8196 30484 8260
rect 31708 8256 31772 8260
rect 31708 8200 31722 8256
rect 31722 8200 31772 8256
rect 31708 8196 31772 8200
rect 32812 8196 32876 8260
rect 33916 8196 33980 8260
rect 35204 8196 35268 8260
rect 36308 8256 36372 8260
rect 36308 8200 36358 8256
rect 36358 8200 36372 8256
rect 36308 8196 36372 8200
rect 37412 8256 37476 8260
rect 37412 8200 37462 8256
rect 37462 8200 37476 8256
rect 37412 8196 37476 8200
rect 38700 8256 38764 8260
rect 38700 8200 38750 8256
rect 38750 8200 38764 8256
rect 38700 8196 38764 8200
rect 40908 8196 40972 8260
rect 42196 8256 42260 8260
rect 42196 8200 42210 8256
rect 42210 8200 42260 8256
rect 42196 8196 42260 8200
rect 43300 8196 43364 8260
rect 90588 8256 90652 8260
rect 90588 8200 90638 8256
rect 90638 8200 90652 8256
rect 90588 8196 90652 8200
rect 90956 8256 91020 8260
rect 90956 8200 91006 8256
rect 91006 8200 91020 8256
rect 90956 8196 91020 8200
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 105924 8188 105988 8192
rect 105924 8132 105928 8188
rect 105928 8132 105984 8188
rect 105984 8132 105988 8188
rect 105924 8128 105988 8132
rect 106004 8188 106068 8192
rect 106004 8132 106008 8188
rect 106008 8132 106064 8188
rect 106064 8132 106068 8188
rect 106004 8128 106068 8132
rect 106084 8188 106148 8192
rect 106084 8132 106088 8188
rect 106088 8132 106144 8188
rect 106144 8132 106148 8188
rect 106084 8128 106148 8132
rect 106164 8188 106228 8192
rect 106164 8132 106168 8188
rect 106168 8132 106224 8188
rect 106224 8132 106228 8188
rect 106164 8128 106228 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 66316 7644 66380 7648
rect 66316 7588 66320 7644
rect 66320 7588 66376 7644
rect 66376 7588 66380 7644
rect 66316 7584 66380 7588
rect 66396 7644 66460 7648
rect 66396 7588 66400 7644
rect 66400 7588 66456 7644
rect 66456 7588 66460 7644
rect 66396 7584 66460 7588
rect 66476 7644 66540 7648
rect 66476 7588 66480 7644
rect 66480 7588 66536 7644
rect 66536 7588 66540 7644
rect 66476 7584 66540 7588
rect 66556 7644 66620 7648
rect 66556 7588 66560 7644
rect 66560 7588 66616 7644
rect 66616 7588 66620 7644
rect 66556 7584 66620 7588
rect 97036 7644 97100 7648
rect 97036 7588 97040 7644
rect 97040 7588 97096 7644
rect 97096 7588 97100 7644
rect 97036 7584 97100 7588
rect 97116 7644 97180 7648
rect 97116 7588 97120 7644
rect 97120 7588 97176 7644
rect 97176 7588 97180 7644
rect 97116 7584 97180 7588
rect 97196 7644 97260 7648
rect 97196 7588 97200 7644
rect 97200 7588 97256 7644
rect 97256 7588 97260 7644
rect 97196 7584 97260 7588
rect 97276 7644 97340 7648
rect 97276 7588 97280 7644
rect 97280 7588 97336 7644
rect 97336 7588 97340 7644
rect 97276 7584 97340 7588
rect 106660 7644 106724 7648
rect 106660 7588 106664 7644
rect 106664 7588 106720 7644
rect 106720 7588 106724 7644
rect 106660 7584 106724 7588
rect 106740 7644 106804 7648
rect 106740 7588 106744 7644
rect 106744 7588 106800 7644
rect 106800 7588 106804 7644
rect 106740 7584 106804 7588
rect 106820 7644 106884 7648
rect 106820 7588 106824 7644
rect 106824 7588 106880 7644
rect 106880 7588 106884 7644
rect 106820 7584 106884 7588
rect 106900 7644 106964 7648
rect 106900 7588 106904 7644
rect 106904 7588 106960 7644
rect 106960 7588 106964 7644
rect 106900 7584 106964 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 96376 7100 96440 7104
rect 96376 7044 96380 7100
rect 96380 7044 96436 7100
rect 96436 7044 96440 7100
rect 96376 7040 96440 7044
rect 96456 7100 96520 7104
rect 96456 7044 96460 7100
rect 96460 7044 96516 7100
rect 96516 7044 96520 7100
rect 96456 7040 96520 7044
rect 96536 7100 96600 7104
rect 96536 7044 96540 7100
rect 96540 7044 96596 7100
rect 96596 7044 96600 7100
rect 96536 7040 96600 7044
rect 96616 7100 96680 7104
rect 96616 7044 96620 7100
rect 96620 7044 96676 7100
rect 96676 7044 96680 7100
rect 96616 7040 96680 7044
rect 105924 7100 105988 7104
rect 105924 7044 105928 7100
rect 105928 7044 105984 7100
rect 105984 7044 105988 7100
rect 105924 7040 105988 7044
rect 106004 7100 106068 7104
rect 106004 7044 106008 7100
rect 106008 7044 106064 7100
rect 106064 7044 106068 7100
rect 106004 7040 106068 7044
rect 106084 7100 106148 7104
rect 106084 7044 106088 7100
rect 106088 7044 106144 7100
rect 106144 7044 106148 7100
rect 106084 7040 106148 7044
rect 106164 7100 106228 7104
rect 106164 7044 106168 7100
rect 106168 7044 106224 7100
rect 106224 7044 106228 7100
rect 106164 7040 106228 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 66316 6556 66380 6560
rect 66316 6500 66320 6556
rect 66320 6500 66376 6556
rect 66376 6500 66380 6556
rect 66316 6496 66380 6500
rect 66396 6556 66460 6560
rect 66396 6500 66400 6556
rect 66400 6500 66456 6556
rect 66456 6500 66460 6556
rect 66396 6496 66460 6500
rect 66476 6556 66540 6560
rect 66476 6500 66480 6556
rect 66480 6500 66536 6556
rect 66536 6500 66540 6556
rect 66476 6496 66540 6500
rect 66556 6556 66620 6560
rect 66556 6500 66560 6556
rect 66560 6500 66616 6556
rect 66616 6500 66620 6556
rect 66556 6496 66620 6500
rect 97036 6556 97100 6560
rect 97036 6500 97040 6556
rect 97040 6500 97096 6556
rect 97096 6500 97100 6556
rect 97036 6496 97100 6500
rect 97116 6556 97180 6560
rect 97116 6500 97120 6556
rect 97120 6500 97176 6556
rect 97176 6500 97180 6556
rect 97116 6496 97180 6500
rect 97196 6556 97260 6560
rect 97196 6500 97200 6556
rect 97200 6500 97256 6556
rect 97256 6500 97260 6556
rect 97196 6496 97260 6500
rect 97276 6556 97340 6560
rect 97276 6500 97280 6556
rect 97280 6500 97336 6556
rect 97336 6500 97340 6556
rect 97276 6496 97340 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 96376 6012 96440 6016
rect 96376 5956 96380 6012
rect 96380 5956 96436 6012
rect 96436 5956 96440 6012
rect 96376 5952 96440 5956
rect 96456 6012 96520 6016
rect 96456 5956 96460 6012
rect 96460 5956 96516 6012
rect 96516 5956 96520 6012
rect 96456 5952 96520 5956
rect 96536 6012 96600 6016
rect 96536 5956 96540 6012
rect 96540 5956 96596 6012
rect 96596 5956 96600 6012
rect 96536 5952 96600 5956
rect 96616 6012 96680 6016
rect 96616 5956 96620 6012
rect 96620 5956 96676 6012
rect 96676 5956 96680 6012
rect 96616 5952 96680 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 66316 5468 66380 5472
rect 66316 5412 66320 5468
rect 66320 5412 66376 5468
rect 66376 5412 66380 5468
rect 66316 5408 66380 5412
rect 66396 5468 66460 5472
rect 66396 5412 66400 5468
rect 66400 5412 66456 5468
rect 66456 5412 66460 5468
rect 66396 5408 66460 5412
rect 66476 5468 66540 5472
rect 66476 5412 66480 5468
rect 66480 5412 66536 5468
rect 66536 5412 66540 5468
rect 66476 5408 66540 5412
rect 66556 5468 66620 5472
rect 66556 5412 66560 5468
rect 66560 5412 66616 5468
rect 66616 5412 66620 5468
rect 66556 5408 66620 5412
rect 97036 5468 97100 5472
rect 97036 5412 97040 5468
rect 97040 5412 97096 5468
rect 97096 5412 97100 5468
rect 97036 5408 97100 5412
rect 97116 5468 97180 5472
rect 97116 5412 97120 5468
rect 97120 5412 97176 5468
rect 97176 5412 97180 5468
rect 97116 5408 97180 5412
rect 97196 5468 97260 5472
rect 97196 5412 97200 5468
rect 97200 5412 97256 5468
rect 97256 5412 97260 5468
rect 97196 5408 97260 5412
rect 97276 5468 97340 5472
rect 97276 5412 97280 5468
rect 97280 5412 97336 5468
rect 97336 5412 97340 5468
rect 97276 5408 97340 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 96376 4924 96440 4928
rect 96376 4868 96380 4924
rect 96380 4868 96436 4924
rect 96436 4868 96440 4924
rect 96376 4864 96440 4868
rect 96456 4924 96520 4928
rect 96456 4868 96460 4924
rect 96460 4868 96516 4924
rect 96516 4868 96520 4924
rect 96456 4864 96520 4868
rect 96536 4924 96600 4928
rect 96536 4868 96540 4924
rect 96540 4868 96596 4924
rect 96596 4868 96600 4924
rect 96536 4864 96600 4868
rect 96616 4924 96680 4928
rect 96616 4868 96620 4924
rect 96620 4868 96676 4924
rect 96676 4868 96680 4924
rect 96616 4864 96680 4868
rect 39804 4524 39868 4588
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 66316 4380 66380 4384
rect 66316 4324 66320 4380
rect 66320 4324 66376 4380
rect 66376 4324 66380 4380
rect 66316 4320 66380 4324
rect 66396 4380 66460 4384
rect 66396 4324 66400 4380
rect 66400 4324 66456 4380
rect 66456 4324 66460 4380
rect 66396 4320 66460 4324
rect 66476 4380 66540 4384
rect 66476 4324 66480 4380
rect 66480 4324 66536 4380
rect 66536 4324 66540 4380
rect 66476 4320 66540 4324
rect 66556 4380 66620 4384
rect 66556 4324 66560 4380
rect 66560 4324 66616 4380
rect 66616 4324 66620 4380
rect 66556 4320 66620 4324
rect 97036 4380 97100 4384
rect 97036 4324 97040 4380
rect 97040 4324 97096 4380
rect 97096 4324 97100 4380
rect 97036 4320 97100 4324
rect 97116 4380 97180 4384
rect 97116 4324 97120 4380
rect 97120 4324 97176 4380
rect 97176 4324 97180 4380
rect 97116 4320 97180 4324
rect 97196 4380 97260 4384
rect 97196 4324 97200 4380
rect 97200 4324 97256 4380
rect 97256 4324 97260 4380
rect 97196 4320 97260 4324
rect 97276 4380 97340 4384
rect 97276 4324 97280 4380
rect 97280 4324 97336 4380
rect 97336 4324 97340 4380
rect 97276 4320 97340 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 96376 3836 96440 3840
rect 96376 3780 96380 3836
rect 96380 3780 96436 3836
rect 96436 3780 96440 3836
rect 96376 3776 96440 3780
rect 96456 3836 96520 3840
rect 96456 3780 96460 3836
rect 96460 3780 96516 3836
rect 96516 3780 96520 3836
rect 96456 3776 96520 3780
rect 96536 3836 96600 3840
rect 96536 3780 96540 3836
rect 96540 3780 96596 3836
rect 96596 3780 96600 3836
rect 96536 3776 96600 3780
rect 96616 3836 96680 3840
rect 96616 3780 96620 3836
rect 96620 3780 96676 3836
rect 96676 3780 96680 3836
rect 96616 3776 96680 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 66316 3292 66380 3296
rect 66316 3236 66320 3292
rect 66320 3236 66376 3292
rect 66376 3236 66380 3292
rect 66316 3232 66380 3236
rect 66396 3292 66460 3296
rect 66396 3236 66400 3292
rect 66400 3236 66456 3292
rect 66456 3236 66460 3292
rect 66396 3232 66460 3236
rect 66476 3292 66540 3296
rect 66476 3236 66480 3292
rect 66480 3236 66536 3292
rect 66536 3236 66540 3292
rect 66476 3232 66540 3236
rect 66556 3292 66620 3296
rect 66556 3236 66560 3292
rect 66560 3236 66616 3292
rect 66616 3236 66620 3292
rect 66556 3232 66620 3236
rect 97036 3292 97100 3296
rect 97036 3236 97040 3292
rect 97040 3236 97096 3292
rect 97096 3236 97100 3292
rect 97036 3232 97100 3236
rect 97116 3292 97180 3296
rect 97116 3236 97120 3292
rect 97120 3236 97176 3292
rect 97176 3236 97180 3292
rect 97116 3232 97180 3236
rect 97196 3292 97260 3296
rect 97196 3236 97200 3292
rect 97200 3236 97256 3292
rect 97256 3236 97260 3292
rect 97196 3232 97260 3236
rect 97276 3292 97340 3296
rect 97276 3236 97280 3292
rect 97280 3236 97336 3292
rect 97336 3236 97340 3292
rect 97276 3232 97340 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 96376 2748 96440 2752
rect 96376 2692 96380 2748
rect 96380 2692 96436 2748
rect 96436 2692 96440 2748
rect 96376 2688 96440 2692
rect 96456 2748 96520 2752
rect 96456 2692 96460 2748
rect 96460 2692 96516 2748
rect 96516 2692 96520 2748
rect 96456 2688 96520 2692
rect 96536 2748 96600 2752
rect 96536 2692 96540 2748
rect 96540 2692 96596 2748
rect 96596 2692 96600 2748
rect 96536 2688 96600 2692
rect 96616 2748 96680 2752
rect 96616 2692 96620 2748
rect 96620 2692 96676 2748
rect 96676 2692 96680 2748
rect 96616 2688 96680 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
rect 66316 2204 66380 2208
rect 66316 2148 66320 2204
rect 66320 2148 66376 2204
rect 66376 2148 66380 2204
rect 66316 2144 66380 2148
rect 66396 2204 66460 2208
rect 66396 2148 66400 2204
rect 66400 2148 66456 2204
rect 66456 2148 66460 2204
rect 66396 2144 66460 2148
rect 66476 2204 66540 2208
rect 66476 2148 66480 2204
rect 66480 2148 66536 2204
rect 66536 2148 66540 2204
rect 66476 2144 66540 2148
rect 66556 2204 66620 2208
rect 66556 2148 66560 2204
rect 66560 2148 66616 2204
rect 66616 2148 66620 2204
rect 66556 2144 66620 2148
rect 97036 2204 97100 2208
rect 97036 2148 97040 2204
rect 97040 2148 97096 2204
rect 97096 2148 97100 2204
rect 97036 2144 97100 2148
rect 97116 2204 97180 2208
rect 97116 2148 97120 2204
rect 97120 2148 97176 2204
rect 97176 2148 97180 2204
rect 97116 2144 97180 2148
rect 97196 2204 97260 2208
rect 97196 2148 97200 2204
rect 97200 2148 97256 2204
rect 97256 2148 97260 2204
rect 97196 2144 97260 2148
rect 97276 2204 97340 2208
rect 97276 2148 97280 2204
rect 97280 2148 97336 2204
rect 97336 2148 97340 2204
rect 97276 2144 97340 2148
<< metal4 >>
rect 4208 126784 4528 127344
rect 4208 126720 4216 126784
rect 4280 126720 4296 126784
rect 4360 126720 4376 126784
rect 4440 126720 4456 126784
rect 4520 126720 4528 126784
rect 4208 126258 4528 126720
rect 4208 126022 4250 126258
rect 4486 126022 4528 126258
rect 4208 125696 4528 126022
rect 4208 125632 4216 125696
rect 4280 125632 4296 125696
rect 4360 125632 4376 125696
rect 4440 125632 4456 125696
rect 4520 125632 4528 125696
rect 4208 124608 4528 125632
rect 4208 124544 4216 124608
rect 4280 124544 4296 124608
rect 4360 124544 4376 124608
rect 4440 124544 4456 124608
rect 4520 124544 4528 124608
rect 4208 123520 4528 124544
rect 4208 123456 4216 123520
rect 4280 123456 4296 123520
rect 4360 123456 4376 123520
rect 4440 123456 4456 123520
rect 4520 123456 4528 123520
rect 4208 122432 4528 123456
rect 4208 122368 4216 122432
rect 4280 122368 4296 122432
rect 4360 122368 4376 122432
rect 4440 122368 4456 122432
rect 4520 122368 4528 122432
rect 4208 121344 4528 122368
rect 4208 121280 4216 121344
rect 4280 121280 4296 121344
rect 4360 121280 4376 121344
rect 4440 121280 4456 121344
rect 4520 121280 4528 121344
rect 4208 120256 4528 121280
rect 4208 120192 4216 120256
rect 4280 120192 4296 120256
rect 4360 120192 4376 120256
rect 4440 120192 4456 120256
rect 4520 120192 4528 120256
rect 4208 119168 4528 120192
rect 4208 119104 4216 119168
rect 4280 119104 4296 119168
rect 4360 119104 4376 119168
rect 4440 119104 4456 119168
rect 4520 119104 4528 119168
rect 4208 118080 4528 119104
rect 4208 118016 4216 118080
rect 4280 118016 4296 118080
rect 4360 118016 4376 118080
rect 4440 118016 4456 118080
rect 4520 118016 4528 118080
rect 4208 116992 4528 118016
rect 4208 116928 4216 116992
rect 4280 116928 4296 116992
rect 4360 116928 4376 116992
rect 4440 116928 4456 116992
rect 4520 116928 4528 116992
rect 4208 115904 4528 116928
rect 4208 115840 4216 115904
rect 4280 115840 4296 115904
rect 4360 115840 4376 115904
rect 4440 115840 4456 115904
rect 4520 115840 4528 115904
rect 4208 114816 4528 115840
rect 4208 114752 4216 114816
rect 4280 114752 4296 114816
rect 4360 114752 4376 114816
rect 4440 114752 4456 114816
rect 4520 114752 4528 114816
rect 4208 113728 4528 114752
rect 4208 113664 4216 113728
rect 4280 113664 4296 113728
rect 4360 113664 4376 113728
rect 4440 113664 4456 113728
rect 4520 113664 4528 113728
rect 4208 112640 4528 113664
rect 4208 112576 4216 112640
rect 4280 112576 4296 112640
rect 4360 112576 4376 112640
rect 4440 112576 4456 112640
rect 4520 112576 4528 112640
rect 4208 111552 4528 112576
rect 4208 111488 4216 111552
rect 4280 111488 4296 111552
rect 4360 111488 4376 111552
rect 4440 111488 4456 111552
rect 4520 111488 4528 111552
rect 4208 110464 4528 111488
rect 4208 110400 4216 110464
rect 4280 110400 4296 110464
rect 4360 110400 4376 110464
rect 4440 110400 4456 110464
rect 4520 110400 4528 110464
rect 4208 109376 4528 110400
rect 4208 109312 4216 109376
rect 4280 109312 4296 109376
rect 4360 109312 4376 109376
rect 4440 109312 4456 109376
rect 4520 109312 4528 109376
rect 4208 108288 4528 109312
rect 4208 108224 4216 108288
rect 4280 108224 4296 108288
rect 4360 108224 4376 108288
rect 4440 108224 4456 108288
rect 4520 108224 4528 108288
rect 4208 107200 4528 108224
rect 4208 107136 4216 107200
rect 4280 107136 4296 107200
rect 4360 107136 4376 107200
rect 4440 107136 4456 107200
rect 4520 107136 4528 107200
rect 4208 106112 4528 107136
rect 4208 106048 4216 106112
rect 4280 106048 4296 106112
rect 4360 106048 4376 106112
rect 4440 106048 4456 106112
rect 4520 106048 4528 106112
rect 4208 105024 4528 106048
rect 4208 104960 4216 105024
rect 4280 104960 4296 105024
rect 4360 104960 4376 105024
rect 4440 104960 4456 105024
rect 4520 104960 4528 105024
rect 4208 103936 4528 104960
rect 4208 103872 4216 103936
rect 4280 103872 4296 103936
rect 4360 103872 4376 103936
rect 4440 103872 4456 103936
rect 4520 103872 4528 103936
rect 4208 102848 4528 103872
rect 4208 102784 4216 102848
rect 4280 102784 4296 102848
rect 4360 102784 4376 102848
rect 4440 102784 4456 102848
rect 4520 102784 4528 102848
rect 4208 101760 4528 102784
rect 4208 101696 4216 101760
rect 4280 101696 4296 101760
rect 4360 101696 4376 101760
rect 4440 101696 4456 101760
rect 4520 101696 4528 101760
rect 4208 100672 4528 101696
rect 4208 100608 4216 100672
rect 4280 100608 4296 100672
rect 4360 100608 4376 100672
rect 4440 100608 4456 100672
rect 4520 100608 4528 100672
rect 4208 99584 4528 100608
rect 4208 99520 4216 99584
rect 4280 99520 4296 99584
rect 4360 99520 4376 99584
rect 4440 99520 4456 99584
rect 4520 99520 4528 99584
rect 4208 98496 4528 99520
rect 4208 98432 4216 98496
rect 4280 98432 4296 98496
rect 4360 98432 4376 98496
rect 4440 98432 4456 98496
rect 4520 98432 4528 98496
rect 4208 97532 4528 98432
rect 4208 97408 4250 97532
rect 4486 97408 4528 97532
rect 4208 97344 4216 97408
rect 4520 97344 4528 97408
rect 4208 97296 4250 97344
rect 4486 97296 4528 97344
rect 4208 96320 4528 97296
rect 4208 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4528 96320
rect 4208 95232 4528 96256
rect 4208 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4528 95232
rect 4208 94144 4528 95168
rect 4208 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4528 94144
rect 4208 93056 4528 94080
rect 4208 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4528 93056
rect 4208 91968 4528 92992
rect 4208 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4528 91968
rect 4208 90880 4528 91904
rect 4208 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4528 90880
rect 4208 89792 4528 90816
rect 4208 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4528 89792
rect 4208 88704 4528 89728
rect 4208 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4528 88704
rect 4208 87616 4528 88640
rect 4208 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4528 87616
rect 4208 86528 4528 87552
rect 4208 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4528 86528
rect 4208 85440 4528 86464
rect 4208 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4528 85440
rect 4208 84352 4528 85376
rect 4208 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4528 84352
rect 4208 83264 4528 84288
rect 4208 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4528 83264
rect 4208 82176 4528 83200
rect 4208 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4528 82176
rect 4208 81088 4528 82112
rect 4208 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4528 81088
rect 4208 80000 4528 81024
rect 4208 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4528 80000
rect 4208 78912 4528 79936
rect 4208 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4528 78912
rect 4208 77824 4528 78848
rect 4208 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4528 77824
rect 4208 76736 4528 77760
rect 4208 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4528 76736
rect 4208 75648 4528 76672
rect 4208 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4528 75648
rect 4208 74560 4528 75584
rect 4208 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4528 74560
rect 4208 73472 4528 74496
rect 4208 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4528 73472
rect 4208 72384 4528 73408
rect 4208 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4528 72384
rect 4208 71296 4528 72320
rect 4208 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4528 71296
rect 4208 70208 4528 71232
rect 4208 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4528 70208
rect 4208 69120 4528 70144
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66896 4296 66944
rect 4360 66896 4376 66944
rect 4440 66896 4456 66944
rect 4520 66880 4528 66944
rect 4208 66660 4250 66880
rect 4486 66660 4528 66880
rect 4208 65856 4528 66660
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 127328 5188 127344
rect 4868 127264 4876 127328
rect 4940 127264 4956 127328
rect 5020 127264 5036 127328
rect 5100 127264 5116 127328
rect 5180 127264 5188 127328
rect 4868 126938 5188 127264
rect 4868 126702 4910 126938
rect 5146 126702 5188 126938
rect 4868 126240 5188 126702
rect 4868 126176 4876 126240
rect 4940 126176 4956 126240
rect 5020 126176 5036 126240
rect 5100 126176 5116 126240
rect 5180 126176 5188 126240
rect 4868 125152 5188 126176
rect 34928 126784 35248 127344
rect 34928 126720 34936 126784
rect 35000 126720 35016 126784
rect 35080 126720 35096 126784
rect 35160 126720 35176 126784
rect 35240 126720 35248 126784
rect 34928 126258 35248 126720
rect 34928 126022 34970 126258
rect 35206 126022 35248 126258
rect 34928 125650 35248 126022
rect 35588 127328 35908 127344
rect 35588 127264 35596 127328
rect 35660 127264 35676 127328
rect 35740 127264 35756 127328
rect 35820 127264 35836 127328
rect 35900 127264 35908 127328
rect 35588 126938 35908 127264
rect 35588 126702 35630 126938
rect 35866 126702 35908 126938
rect 35588 126240 35908 126702
rect 35588 126176 35596 126240
rect 35660 126176 35676 126240
rect 35740 126176 35756 126240
rect 35820 126176 35836 126240
rect 35900 126176 35908 126240
rect 35588 125650 35908 126176
rect 65648 126784 65968 127344
rect 65648 126720 65656 126784
rect 65720 126720 65736 126784
rect 65800 126720 65816 126784
rect 65880 126720 65896 126784
rect 65960 126720 65968 126784
rect 65648 126258 65968 126720
rect 46059 126036 46125 126037
rect 46059 125972 46060 126036
rect 46124 125972 46125 126036
rect 46059 125971 46125 125972
rect 53603 126036 53669 126037
rect 53603 125972 53604 126036
rect 53668 125972 53669 126036
rect 53603 125971 53669 125972
rect 65648 126022 65690 126258
rect 65926 126022 65968 126258
rect 4868 125088 4876 125152
rect 4940 125088 4956 125152
rect 5020 125088 5036 125152
rect 5100 125088 5116 125152
rect 5180 125088 5188 125152
rect 4868 124064 5188 125088
rect 36074 124268 36140 124269
rect 36074 124204 36075 124268
rect 36139 124204 36140 124268
rect 36074 124203 36140 124204
rect 38570 124268 38636 124269
rect 38570 124204 38571 124268
rect 38635 124204 38636 124268
rect 38570 124203 38636 124204
rect 41066 124268 41132 124269
rect 41066 124204 41067 124268
rect 41131 124204 41132 124268
rect 41066 124203 41132 124204
rect 4868 124000 4876 124064
rect 4940 124000 4956 124064
rect 5020 124000 5036 124064
rect 5100 124000 5116 124064
rect 5180 124000 5188 124064
rect 4868 122976 5188 124000
rect 36077 123676 36137 124203
rect 38573 123676 38633 124203
rect 41069 123676 41129 124203
rect 43562 124132 43628 124133
rect 43562 124068 43563 124132
rect 43627 124068 43628 124132
rect 43562 124067 43628 124068
rect 43565 123676 43625 124067
rect 46062 123676 46122 125971
rect 51027 125628 51093 125629
rect 51027 125564 51028 125628
rect 51092 125564 51093 125628
rect 51027 125563 51093 125564
rect 48543 124268 48609 124269
rect 48543 124204 48544 124268
rect 48608 124204 48609 124268
rect 48543 124203 48609 124204
rect 48546 123676 48606 124203
rect 51030 124130 51090 125563
rect 53606 124130 53666 125971
rect 65648 125834 65968 126022
rect 66308 127328 66628 127344
rect 66308 127264 66316 127328
rect 66380 127264 66396 127328
rect 66460 127264 66476 127328
rect 66540 127264 66556 127328
rect 66620 127264 66628 127328
rect 66308 126938 66628 127264
rect 66308 126702 66350 126938
rect 66586 126702 66628 126938
rect 66308 126240 66628 126702
rect 96368 126784 96688 127344
rect 96368 126720 96376 126784
rect 96440 126720 96456 126784
rect 96520 126720 96536 126784
rect 96600 126720 96616 126784
rect 96680 126720 96688 126784
rect 73475 126444 73541 126445
rect 73475 126380 73476 126444
rect 73540 126380 73541 126444
rect 73475 126379 73541 126380
rect 66308 126176 66316 126240
rect 66380 126176 66396 126240
rect 66460 126176 66476 126240
rect 66540 126176 66556 126240
rect 66620 126176 66628 126240
rect 58571 125764 58637 125765
rect 58571 125700 58572 125764
rect 58636 125700 58637 125764
rect 58571 125699 58637 125700
rect 55995 125628 56061 125629
rect 55995 125564 55996 125628
rect 56060 125564 56061 125628
rect 55995 125563 56061 125564
rect 51030 124070 51113 124130
rect 51053 123676 51113 124070
rect 53549 124070 53666 124130
rect 55998 124130 56058 125563
rect 58574 124130 58634 125699
rect 66308 125650 66628 126176
rect 61147 125628 61213 125629
rect 61147 125564 61148 125628
rect 61212 125564 61213 125628
rect 61147 125563 61213 125564
rect 61150 124130 61210 125563
rect 63539 125220 63605 125221
rect 63539 125156 63540 125220
rect 63604 125156 63605 125220
rect 63539 125155 63605 125156
rect 55998 124070 56105 124130
rect 53549 123676 53609 124070
rect 56045 123676 56105 124070
rect 58541 124070 58634 124130
rect 61058 124070 61210 124130
rect 58541 123676 58601 124070
rect 61058 123676 61118 124070
rect 63542 123676 63602 125155
rect 66026 124268 66092 124269
rect 66026 124204 66027 124268
rect 66091 124204 66092 124268
rect 66026 124203 66092 124204
rect 68522 124268 68588 124269
rect 68522 124204 68523 124268
rect 68587 124204 68588 124268
rect 68522 124203 68588 124204
rect 71018 124268 71084 124269
rect 71018 124204 71019 124268
rect 71083 124204 71084 124268
rect 71018 124203 71084 124204
rect 66029 123676 66089 124203
rect 68525 123676 68585 124203
rect 71021 123676 71081 124203
rect 73478 124130 73538 126379
rect 96368 126258 96688 126720
rect 96368 126022 96410 126258
rect 96646 126022 96688 126258
rect 96368 125650 96688 126022
rect 97028 127328 97348 127344
rect 97028 127264 97036 127328
rect 97100 127264 97116 127328
rect 97180 127264 97196 127328
rect 97260 127264 97276 127328
rect 97340 127264 97348 127328
rect 97028 126938 97348 127264
rect 97028 126702 97070 126938
rect 97306 126702 97348 126938
rect 97028 126240 97348 126702
rect 97028 126176 97036 126240
rect 97100 126176 97116 126240
rect 97180 126176 97196 126240
rect 97260 126176 97276 126240
rect 97340 126176 97348 126240
rect 97028 125650 97348 126176
rect 105916 126784 106236 126800
rect 105916 126720 105924 126784
rect 105988 126720 106004 126784
rect 106068 126720 106084 126784
rect 106148 126720 106164 126784
rect 106228 126720 106236 126784
rect 105916 126258 106236 126720
rect 105916 126022 105958 126258
rect 106194 126022 106236 126258
rect 105916 125696 106236 126022
rect 105916 125632 105924 125696
rect 105988 125632 106004 125696
rect 106068 125632 106084 125696
rect 106148 125632 106164 125696
rect 106228 125632 106236 125696
rect 105916 124608 106236 125632
rect 105916 124544 105924 124608
rect 105988 124544 106004 124608
rect 106068 124544 106084 124608
rect 106148 124544 106164 124608
rect 106228 124544 106236 124608
rect 73478 124070 73577 124130
rect 73517 123676 73577 124070
rect 95860 124070 96170 124130
rect 86141 123996 86207 123997
rect 86141 123932 86142 123996
rect 86206 123932 86207 123996
rect 86141 123931 86207 123932
rect 86144 123676 86204 123931
rect 87309 123860 87375 123861
rect 87309 123796 87310 123860
rect 87374 123796 87375 123860
rect 87309 123795 87375 123796
rect 87312 123676 87372 123795
rect 95860 123676 95920 124070
rect 96110 123861 96170 124070
rect 96107 123860 96173 123861
rect 96107 123796 96108 123860
rect 96172 123796 96173 123860
rect 96107 123795 96173 123796
rect 4868 122912 4876 122976
rect 4940 122912 4956 122976
rect 5020 122912 5036 122976
rect 5100 122912 5116 122976
rect 5180 122912 5188 122976
rect 4868 121888 5188 122912
rect 4868 121824 4876 121888
rect 4940 121824 4956 121888
rect 5020 121824 5036 121888
rect 5100 121824 5116 121888
rect 5180 121824 5188 121888
rect 4868 120800 5188 121824
rect 4868 120736 4876 120800
rect 4940 120736 4956 120800
rect 5020 120736 5036 120800
rect 5100 120736 5116 120800
rect 5180 120736 5188 120800
rect 4868 119712 5188 120736
rect 4868 119648 4876 119712
rect 4940 119648 4956 119712
rect 5020 119648 5036 119712
rect 5100 119648 5116 119712
rect 5180 119648 5188 119712
rect 4868 118624 5188 119648
rect 4868 118560 4876 118624
rect 4940 118560 4956 118624
rect 5020 118560 5036 118624
rect 5100 118560 5116 118624
rect 5180 118560 5188 118624
rect 4868 117536 5188 118560
rect 4868 117472 4876 117536
rect 4940 117472 4956 117536
rect 5020 117472 5036 117536
rect 5100 117472 5116 117536
rect 5180 117472 5188 117536
rect 4868 116448 5188 117472
rect 4868 116384 4876 116448
rect 4940 116384 4956 116448
rect 5020 116384 5036 116448
rect 5100 116384 5116 116448
rect 5180 116384 5188 116448
rect 4868 115360 5188 116384
rect 4868 115296 4876 115360
rect 4940 115296 4956 115360
rect 5020 115296 5036 115360
rect 5100 115296 5116 115360
rect 5180 115296 5188 115360
rect 4868 114272 5188 115296
rect 4868 114208 4876 114272
rect 4940 114208 4956 114272
rect 5020 114208 5036 114272
rect 5100 114208 5116 114272
rect 5180 114208 5188 114272
rect 4868 113184 5188 114208
rect 4868 113120 4876 113184
rect 4940 113120 4956 113184
rect 5020 113120 5036 113184
rect 5100 113120 5116 113184
rect 5180 113120 5188 113184
rect 4868 112096 5188 113120
rect 4868 112032 4876 112096
rect 4940 112032 4956 112096
rect 5020 112032 5036 112096
rect 5100 112032 5116 112096
rect 5180 112032 5188 112096
rect 4868 111008 5188 112032
rect 4868 110944 4876 111008
rect 4940 110944 4956 111008
rect 5020 110944 5036 111008
rect 5100 110944 5116 111008
rect 5180 110944 5188 111008
rect 4868 109920 5188 110944
rect 4868 109856 4876 109920
rect 4940 109856 4956 109920
rect 5020 109856 5036 109920
rect 5100 109856 5116 109920
rect 5180 109856 5188 109920
rect 4868 108832 5188 109856
rect 4868 108768 4876 108832
rect 4940 108768 4956 108832
rect 5020 108768 5036 108832
rect 5100 108768 5116 108832
rect 5180 108768 5188 108832
rect 4868 107744 5188 108768
rect 4868 107680 4876 107744
rect 4940 107680 4956 107744
rect 5020 107680 5036 107744
rect 5100 107680 5116 107744
rect 5180 107680 5188 107744
rect 4868 106656 5188 107680
rect 4868 106592 4876 106656
rect 4940 106592 4956 106656
rect 5020 106592 5036 106656
rect 5100 106592 5116 106656
rect 5180 106592 5188 106656
rect 4868 105568 5188 106592
rect 4868 105504 4876 105568
rect 4940 105504 4956 105568
rect 5020 105504 5036 105568
rect 5100 105504 5116 105568
rect 5180 105504 5188 105568
rect 4868 104480 5188 105504
rect 4868 104416 4876 104480
rect 4940 104416 4956 104480
rect 5020 104416 5036 104480
rect 5100 104416 5116 104480
rect 5180 104416 5188 104480
rect 4868 103392 5188 104416
rect 4868 103328 4876 103392
rect 4940 103328 4956 103392
rect 5020 103328 5036 103392
rect 5100 103328 5116 103392
rect 5180 103328 5188 103392
rect 4868 102304 5188 103328
rect 4868 102240 4876 102304
rect 4940 102240 4956 102304
rect 5020 102240 5036 102304
rect 5100 102240 5116 102304
rect 5180 102240 5188 102304
rect 4868 101216 5188 102240
rect 4868 101152 4876 101216
rect 4940 101152 4956 101216
rect 5020 101152 5036 101216
rect 5100 101152 5116 101216
rect 5180 101152 5188 101216
rect 4868 100128 5188 101152
rect 4868 100064 4876 100128
rect 4940 100064 4956 100128
rect 5020 100064 5036 100128
rect 5100 100064 5116 100128
rect 5180 100064 5188 100128
rect 4868 99040 5188 100064
rect 4868 98976 4876 99040
rect 4940 98976 4956 99040
rect 5020 98976 5036 99040
rect 5100 98976 5116 99040
rect 5180 98976 5188 99040
rect 4868 98192 5188 98976
rect 105916 123520 106236 124544
rect 105916 123456 105924 123520
rect 105988 123456 106004 123520
rect 106068 123456 106084 123520
rect 106148 123456 106164 123520
rect 106228 123456 106236 123520
rect 105916 122432 106236 123456
rect 105916 122368 105924 122432
rect 105988 122368 106004 122432
rect 106068 122368 106084 122432
rect 106148 122368 106164 122432
rect 106228 122368 106236 122432
rect 105916 121344 106236 122368
rect 105916 121280 105924 121344
rect 105988 121280 106004 121344
rect 106068 121280 106084 121344
rect 106148 121280 106164 121344
rect 106228 121280 106236 121344
rect 105916 120256 106236 121280
rect 105916 120192 105924 120256
rect 105988 120192 106004 120256
rect 106068 120192 106084 120256
rect 106148 120192 106164 120256
rect 106228 120192 106236 120256
rect 105916 119168 106236 120192
rect 105916 119104 105924 119168
rect 105988 119104 106004 119168
rect 106068 119104 106084 119168
rect 106148 119104 106164 119168
rect 106228 119104 106236 119168
rect 105916 118080 106236 119104
rect 105916 118016 105924 118080
rect 105988 118016 106004 118080
rect 106068 118016 106084 118080
rect 106148 118016 106164 118080
rect 106228 118016 106236 118080
rect 105916 116992 106236 118016
rect 105916 116928 105924 116992
rect 105988 116928 106004 116992
rect 106068 116928 106084 116992
rect 106148 116928 106164 116992
rect 106228 116928 106236 116992
rect 105916 115904 106236 116928
rect 105916 115840 105924 115904
rect 105988 115840 106004 115904
rect 106068 115840 106084 115904
rect 106148 115840 106164 115904
rect 106228 115840 106236 115904
rect 105916 114816 106236 115840
rect 105916 114752 105924 114816
rect 105988 114752 106004 114816
rect 106068 114752 106084 114816
rect 106148 114752 106164 114816
rect 106228 114752 106236 114816
rect 105916 113728 106236 114752
rect 105916 113664 105924 113728
rect 105988 113664 106004 113728
rect 106068 113664 106084 113728
rect 106148 113664 106164 113728
rect 106228 113664 106236 113728
rect 105916 112640 106236 113664
rect 105916 112576 105924 112640
rect 105988 112576 106004 112640
rect 106068 112576 106084 112640
rect 106148 112576 106164 112640
rect 106228 112576 106236 112640
rect 105916 111552 106236 112576
rect 105916 111488 105924 111552
rect 105988 111488 106004 111552
rect 106068 111488 106084 111552
rect 106148 111488 106164 111552
rect 106228 111488 106236 111552
rect 105916 110464 106236 111488
rect 105916 110400 105924 110464
rect 105988 110400 106004 110464
rect 106068 110400 106084 110464
rect 106148 110400 106164 110464
rect 106228 110400 106236 110464
rect 105916 109376 106236 110400
rect 105916 109312 105924 109376
rect 105988 109312 106004 109376
rect 106068 109312 106084 109376
rect 106148 109312 106164 109376
rect 106228 109312 106236 109376
rect 105916 108288 106236 109312
rect 105916 108224 105924 108288
rect 105988 108224 106004 108288
rect 106068 108224 106084 108288
rect 106148 108224 106164 108288
rect 106228 108224 106236 108288
rect 105916 107200 106236 108224
rect 105916 107136 105924 107200
rect 105988 107136 106004 107200
rect 106068 107136 106084 107200
rect 106148 107136 106164 107200
rect 106228 107136 106236 107200
rect 105916 106112 106236 107136
rect 105916 106048 105924 106112
rect 105988 106048 106004 106112
rect 106068 106048 106084 106112
rect 106148 106048 106164 106112
rect 106228 106048 106236 106112
rect 105916 105024 106236 106048
rect 105916 104960 105924 105024
rect 105988 104960 106004 105024
rect 106068 104960 106084 105024
rect 106148 104960 106164 105024
rect 106228 104960 106236 105024
rect 105916 103936 106236 104960
rect 105916 103872 105924 103936
rect 105988 103872 106004 103936
rect 106068 103872 106084 103936
rect 106148 103872 106164 103936
rect 106228 103872 106236 103936
rect 105916 102848 106236 103872
rect 105916 102784 105924 102848
rect 105988 102784 106004 102848
rect 106068 102784 106084 102848
rect 106148 102784 106164 102848
rect 106228 102784 106236 102848
rect 105916 101760 106236 102784
rect 105916 101696 105924 101760
rect 105988 101696 106004 101760
rect 106068 101696 106084 101760
rect 106148 101696 106164 101760
rect 106228 101696 106236 101760
rect 105916 100672 106236 101696
rect 105916 100608 105924 100672
rect 105988 100608 106004 100672
rect 106068 100608 106084 100672
rect 106148 100608 106164 100672
rect 106228 100608 106236 100672
rect 105916 99584 106236 100608
rect 105916 99520 105924 99584
rect 105988 99520 106004 99584
rect 106068 99520 106084 99584
rect 106148 99520 106164 99584
rect 106228 99520 106236 99584
rect 105916 98496 106236 99520
rect 105916 98432 105924 98496
rect 105988 98432 106004 98496
rect 106068 98432 106084 98496
rect 106148 98432 106164 98496
rect 106228 98432 106236 98496
rect 4868 97956 4910 98192
rect 5146 97956 5188 98192
rect 4868 97952 5188 97956
rect 4868 97888 4876 97952
rect 4940 97888 4956 97952
rect 5020 97888 5036 97952
rect 5100 97888 5116 97952
rect 5180 97888 5188 97952
rect 10696 98192 11044 98234
rect 10696 97956 10752 98192
rect 10988 97956 11044 98192
rect 10696 97914 11044 97956
rect 100936 98192 101284 98234
rect 100936 97956 100992 98192
rect 101228 97956 101284 98192
rect 100936 97914 101284 97956
rect 4868 96864 5188 97888
rect 10000 97532 10348 97574
rect 10000 97296 10056 97532
rect 10292 97296 10348 97532
rect 10000 97254 10348 97296
rect 101632 97532 101980 97574
rect 101632 97296 101688 97532
rect 101924 97296 101980 97532
rect 101632 97254 101980 97296
rect 105916 97532 106236 98432
rect 105916 97408 105958 97532
rect 106194 97408 106236 97532
rect 105916 97344 105924 97408
rect 106228 97344 106236 97408
rect 105916 97296 105958 97344
rect 106194 97296 106236 97344
rect 4868 96800 4876 96864
rect 4940 96800 4956 96864
rect 5020 96800 5036 96864
rect 5100 96800 5116 96864
rect 5180 96800 5188 96864
rect 4868 95776 5188 96800
rect 4868 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5188 95776
rect 4868 94688 5188 95712
rect 4868 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5188 94688
rect 4868 93600 5188 94624
rect 4868 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5188 93600
rect 4868 92512 5188 93536
rect 4868 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5188 92512
rect 4868 91424 5188 92448
rect 4868 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5188 91424
rect 4868 90336 5188 91360
rect 4868 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5188 90336
rect 4868 89248 5188 90272
rect 4868 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5188 89248
rect 4868 88160 5188 89184
rect 4868 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5188 88160
rect 4868 87072 5188 88096
rect 4868 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5188 87072
rect 4868 85984 5188 87008
rect 4868 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5188 85984
rect 4868 84896 5188 85920
rect 4868 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5188 84896
rect 4868 83808 5188 84832
rect 4868 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5188 83808
rect 4868 82720 5188 83744
rect 4868 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5188 82720
rect 4868 81632 5188 82656
rect 4868 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5188 81632
rect 4868 80544 5188 81568
rect 4868 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5188 80544
rect 4868 79456 5188 80480
rect 4868 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5188 79456
rect 4868 78368 5188 79392
rect 4868 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5188 78368
rect 4868 77280 5188 78304
rect 4868 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5188 77280
rect 4868 76192 5188 77216
rect 4868 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5188 76192
rect 4868 75104 5188 76128
rect 4868 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5188 75104
rect 4868 74016 5188 75040
rect 4868 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5188 74016
rect 4868 72928 5188 73952
rect 4868 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5188 72928
rect 4868 71840 5188 72864
rect 4868 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5188 71840
rect 4868 70752 5188 71776
rect 4868 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5188 70752
rect 4868 69664 5188 70688
rect 105916 96320 106236 97296
rect 105916 96256 105924 96320
rect 105988 96256 106004 96320
rect 106068 96256 106084 96320
rect 106148 96256 106164 96320
rect 106228 96256 106236 96320
rect 105916 95232 106236 96256
rect 105916 95168 105924 95232
rect 105988 95168 106004 95232
rect 106068 95168 106084 95232
rect 106148 95168 106164 95232
rect 106228 95168 106236 95232
rect 105916 94144 106236 95168
rect 105916 94080 105924 94144
rect 105988 94080 106004 94144
rect 106068 94080 106084 94144
rect 106148 94080 106164 94144
rect 106228 94080 106236 94144
rect 105916 93056 106236 94080
rect 105916 92992 105924 93056
rect 105988 92992 106004 93056
rect 106068 92992 106084 93056
rect 106148 92992 106164 93056
rect 106228 92992 106236 93056
rect 105916 91968 106236 92992
rect 105916 91904 105924 91968
rect 105988 91904 106004 91968
rect 106068 91904 106084 91968
rect 106148 91904 106164 91968
rect 106228 91904 106236 91968
rect 105916 90880 106236 91904
rect 105916 90816 105924 90880
rect 105988 90816 106004 90880
rect 106068 90816 106084 90880
rect 106148 90816 106164 90880
rect 106228 90816 106236 90880
rect 105916 89792 106236 90816
rect 105916 89728 105924 89792
rect 105988 89728 106004 89792
rect 106068 89728 106084 89792
rect 106148 89728 106164 89792
rect 106228 89728 106236 89792
rect 105916 88704 106236 89728
rect 105916 88640 105924 88704
rect 105988 88640 106004 88704
rect 106068 88640 106084 88704
rect 106148 88640 106164 88704
rect 106228 88640 106236 88704
rect 105916 87616 106236 88640
rect 105916 87552 105924 87616
rect 105988 87552 106004 87616
rect 106068 87552 106084 87616
rect 106148 87552 106164 87616
rect 106228 87552 106236 87616
rect 105916 86528 106236 87552
rect 105916 86464 105924 86528
rect 105988 86464 106004 86528
rect 106068 86464 106084 86528
rect 106148 86464 106164 86528
rect 106228 86464 106236 86528
rect 105916 85440 106236 86464
rect 105916 85376 105924 85440
rect 105988 85376 106004 85440
rect 106068 85376 106084 85440
rect 106148 85376 106164 85440
rect 106228 85376 106236 85440
rect 105916 84352 106236 85376
rect 105916 84288 105924 84352
rect 105988 84288 106004 84352
rect 106068 84288 106084 84352
rect 106148 84288 106164 84352
rect 106228 84288 106236 84352
rect 105916 83264 106236 84288
rect 105916 83200 105924 83264
rect 105988 83200 106004 83264
rect 106068 83200 106084 83264
rect 106148 83200 106164 83264
rect 106228 83200 106236 83264
rect 105916 82176 106236 83200
rect 105916 82112 105924 82176
rect 105988 82112 106004 82176
rect 106068 82112 106084 82176
rect 106148 82112 106164 82176
rect 106228 82112 106236 82176
rect 105916 81088 106236 82112
rect 105916 81024 105924 81088
rect 105988 81024 106004 81088
rect 106068 81024 106084 81088
rect 106148 81024 106164 81088
rect 106228 81024 106236 81088
rect 105916 80000 106236 81024
rect 105916 79936 105924 80000
rect 105988 79936 106004 80000
rect 106068 79936 106084 80000
rect 106148 79936 106164 80000
rect 106228 79936 106236 80000
rect 105916 78912 106236 79936
rect 105916 78848 105924 78912
rect 105988 78848 106004 78912
rect 106068 78848 106084 78912
rect 106148 78848 106164 78912
rect 106228 78848 106236 78912
rect 105916 77824 106236 78848
rect 105916 77760 105924 77824
rect 105988 77760 106004 77824
rect 106068 77760 106084 77824
rect 106148 77760 106164 77824
rect 106228 77760 106236 77824
rect 105916 76736 106236 77760
rect 105916 76672 105924 76736
rect 105988 76672 106004 76736
rect 106068 76672 106084 76736
rect 106148 76672 106164 76736
rect 106228 76672 106236 76736
rect 105916 75648 106236 76672
rect 105916 75584 105924 75648
rect 105988 75584 106004 75648
rect 106068 75584 106084 75648
rect 106148 75584 106164 75648
rect 106228 75584 106236 75648
rect 105916 74560 106236 75584
rect 105916 74496 105924 74560
rect 105988 74496 106004 74560
rect 106068 74496 106084 74560
rect 106148 74496 106164 74560
rect 106228 74496 106236 74560
rect 105916 73472 106236 74496
rect 105916 73408 105924 73472
rect 105988 73408 106004 73472
rect 106068 73408 106084 73472
rect 106148 73408 106164 73472
rect 106228 73408 106236 73472
rect 105916 72384 106236 73408
rect 105916 72320 105924 72384
rect 105988 72320 106004 72384
rect 106068 72320 106084 72384
rect 106148 72320 106164 72384
rect 106228 72320 106236 72384
rect 105916 71296 106236 72320
rect 105916 71232 105924 71296
rect 105988 71232 106004 71296
rect 106068 71232 106084 71296
rect 106148 71232 106164 71296
rect 106228 71232 106236 71296
rect 105916 70208 106236 71232
rect 105916 70144 105924 70208
rect 105988 70144 106004 70208
rect 106068 70144 106084 70208
rect 106148 70144 106164 70208
rect 106228 70144 106236 70208
rect 4868 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5188 69664
rect 4868 68576 5188 69600
rect 4868 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5188 68576
rect 4868 67556 5188 68512
rect 16070 67693 16130 70038
rect 23440 69597 23500 70038
rect 24626 69597 24686 70038
rect 25776 69597 25836 70038
rect 26944 69597 27004 70038
rect 28112 69597 28172 70038
rect 29280 69730 29340 70038
rect 29280 69670 29378 69730
rect 23437 69596 23503 69597
rect 23437 69532 23438 69596
rect 23502 69532 23503 69596
rect 23437 69531 23503 69532
rect 24623 69596 24689 69597
rect 24623 69532 24624 69596
rect 24688 69532 24689 69596
rect 24623 69531 24689 69532
rect 25773 69596 25839 69597
rect 25773 69532 25774 69596
rect 25838 69532 25839 69596
rect 25773 69531 25839 69532
rect 26941 69596 27007 69597
rect 26941 69532 26942 69596
rect 27006 69532 27007 69596
rect 26941 69531 27007 69532
rect 28109 69596 28175 69597
rect 28109 69532 28110 69596
rect 28174 69532 28175 69596
rect 28109 69531 28175 69532
rect 29318 69325 29378 69670
rect 30448 69597 30508 70038
rect 31616 69597 31676 70038
rect 32784 69597 32844 70038
rect 33952 69869 34012 70038
rect 33949 69868 34015 69869
rect 33949 69804 33950 69868
rect 34014 69804 34015 69868
rect 33949 69803 34015 69804
rect 33952 69597 34012 69803
rect 35120 69597 35180 70038
rect 36310 69597 36370 70040
rect 37456 69869 37516 70038
rect 38624 69869 38684 70038
rect 39792 69869 39852 70038
rect 40960 69869 41020 70038
rect 37453 69868 37519 69869
rect 37453 69804 37454 69868
rect 37518 69804 37519 69868
rect 37453 69803 37519 69804
rect 38621 69868 38687 69869
rect 38621 69804 38622 69868
rect 38686 69804 38687 69868
rect 38621 69803 38687 69804
rect 39789 69868 39855 69869
rect 39789 69804 39790 69868
rect 39854 69804 39855 69868
rect 39789 69803 39855 69804
rect 40957 69868 41023 69869
rect 40957 69804 40958 69868
rect 41022 69804 41023 69868
rect 40957 69803 41023 69804
rect 42128 69597 42188 70038
rect 43296 69869 43356 70038
rect 43293 69868 43359 69869
rect 43293 69804 43294 69868
rect 43358 69804 43359 69868
rect 43293 69803 43359 69804
rect 90529 69597 90589 70038
rect 90682 69869 90742 70038
rect 90679 69868 90745 69869
rect 90679 69804 90680 69868
rect 90744 69804 90745 69868
rect 90679 69803 90745 69804
rect 90816 69730 90876 70038
rect 90774 69670 90876 69730
rect 30445 69596 30511 69597
rect 30445 69532 30446 69596
rect 30510 69532 30511 69596
rect 30445 69531 30511 69532
rect 31613 69596 31679 69597
rect 31613 69532 31614 69596
rect 31678 69532 31679 69596
rect 32784 69596 32877 69597
rect 32784 69534 32812 69596
rect 31613 69531 31679 69532
rect 32811 69532 32812 69534
rect 32876 69532 32877 69596
rect 32811 69531 32877 69532
rect 33949 69596 34015 69597
rect 33949 69532 33950 69596
rect 34014 69532 34015 69596
rect 33949 69531 34015 69532
rect 35117 69596 35183 69597
rect 35117 69532 35118 69596
rect 35182 69532 35183 69596
rect 35117 69531 35183 69532
rect 36307 69596 36373 69597
rect 36307 69532 36308 69596
rect 36372 69532 36373 69596
rect 36307 69531 36373 69532
rect 42125 69596 42191 69597
rect 42125 69532 42126 69596
rect 42190 69532 42191 69596
rect 42125 69531 42191 69532
rect 90526 69596 90592 69597
rect 90526 69532 90527 69596
rect 90591 69532 90592 69596
rect 90526 69531 90592 69532
rect 29315 69324 29381 69325
rect 29315 69260 29316 69324
rect 29380 69260 29381 69324
rect 29315 69259 29381 69260
rect 90774 68781 90834 69670
rect 105916 69120 106236 70144
rect 105916 69056 105924 69120
rect 105988 69056 106004 69120
rect 106068 69056 106084 69120
rect 106148 69056 106164 69120
rect 106228 69056 106236 69120
rect 90771 68780 90837 68781
rect 90771 68716 90772 68780
rect 90836 68716 90837 68780
rect 90771 68715 90837 68716
rect 16067 67692 16133 67693
rect 16067 67628 16068 67692
rect 16132 67628 16133 67692
rect 16067 67627 16133 67628
rect 4868 67488 4910 67556
rect 5146 67488 5188 67556
rect 4868 67424 4876 67488
rect 5180 67424 5188 67488
rect 4868 67320 4910 67424
rect 5146 67320 5188 67424
rect 4868 66400 5188 67320
rect 4868 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5188 66400
rect 4868 65312 5188 66336
rect 34928 66944 35248 67880
rect 34928 66880 34936 66944
rect 35000 66896 35016 66944
rect 35080 66896 35096 66944
rect 35160 66896 35176 66944
rect 35240 66880 35248 66944
rect 34928 66660 34970 66880
rect 35206 66660 35248 66880
rect 34928 65856 35248 66660
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 65650 35248 65792
rect 35588 67556 35908 68064
rect 35588 67488 35630 67556
rect 35866 67488 35908 67556
rect 35588 67424 35596 67488
rect 35900 67424 35908 67488
rect 35588 67320 35630 67424
rect 35866 67320 35908 67424
rect 35588 66400 35908 67320
rect 65648 68032 65968 68064
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 66944 65968 67968
rect 65648 66880 65656 66944
rect 65720 66896 65736 66944
rect 65800 66896 65816 66944
rect 65880 66896 65896 66944
rect 65960 66880 65968 66944
rect 63539 66740 63605 66741
rect 63539 66676 63540 66740
rect 63604 66676 63605 66740
rect 63539 66675 63605 66676
rect 36123 66604 36189 66605
rect 36123 66540 36124 66604
rect 36188 66540 36189 66604
rect 36123 66539 36189 66540
rect 51027 66604 51093 66605
rect 51027 66540 51028 66604
rect 51092 66540 51093 66604
rect 51027 66539 51093 66540
rect 35588 66336 35596 66400
rect 35660 66336 35676 66400
rect 35740 66336 35756 66400
rect 35820 66336 35836 66400
rect 35900 66336 35908 66400
rect 35588 65650 35908 66336
rect 4868 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5188 65312
rect 4868 64224 5188 65248
rect 36126 64290 36186 66539
rect 41091 66332 41157 66333
rect 41091 66268 41092 66332
rect 41156 66268 41157 66332
rect 41091 66267 41157 66268
rect 41094 64290 41154 66267
rect 46059 66196 46125 66197
rect 46059 66132 46060 66196
rect 46124 66132 46125 66196
rect 46059 66131 46125 66132
rect 43483 65516 43549 65517
rect 43483 65452 43484 65516
rect 43548 65452 43549 65516
rect 43483 65451 43549 65452
rect 4868 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5188 64224
rect 4868 63136 5188 64160
rect 36077 64230 36186 64290
rect 41069 64230 41154 64290
rect 43486 64290 43546 65451
rect 43486 64230 43625 64290
rect 36077 63676 36137 64230
rect 38570 64156 38636 64157
rect 38570 64092 38571 64156
rect 38635 64092 38636 64156
rect 38570 64091 38636 64092
rect 38573 63676 38633 64091
rect 41069 63676 41129 64230
rect 43565 63676 43625 64230
rect 46062 63676 46122 66131
rect 51030 64290 51090 66539
rect 53603 65924 53669 65925
rect 53603 65860 53604 65924
rect 53668 65860 53669 65924
rect 53603 65859 53669 65860
rect 53606 64290 53666 65859
rect 51030 64230 51113 64290
rect 48543 64156 48609 64157
rect 48543 64092 48544 64156
rect 48608 64092 48609 64156
rect 48543 64091 48609 64092
rect 48546 63676 48606 64091
rect 51053 63676 51113 64230
rect 53549 64230 53666 64290
rect 53549 63676 53609 64230
rect 56042 64156 56108 64157
rect 56042 64092 56043 64156
rect 56107 64092 56108 64156
rect 56042 64091 56108 64092
rect 56045 63676 56105 64091
rect 58538 64020 58604 64021
rect 58538 63956 58539 64020
rect 58603 63956 58604 64020
rect 58538 63955 58604 63956
rect 58541 63676 58601 63955
rect 61055 63884 61121 63885
rect 61055 63820 61056 63884
rect 61120 63820 61121 63884
rect 61055 63819 61121 63820
rect 61058 63676 61118 63819
rect 63542 63676 63602 66675
rect 65648 66660 65690 66880
rect 65926 66660 65968 66880
rect 65648 65856 65968 66660
rect 66308 67556 66628 68064
rect 96368 68032 96688 68064
rect 96368 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96688 68032
rect 86171 67692 86237 67693
rect 86171 67628 86172 67692
rect 86236 67628 86237 67692
rect 86171 67627 86237 67628
rect 66308 67488 66350 67556
rect 66586 67488 66628 67556
rect 66308 67424 66316 67488
rect 66620 67424 66628 67488
rect 66308 67320 66350 67424
rect 66586 67320 66628 67424
rect 66115 66604 66181 66605
rect 66115 66540 66116 66604
rect 66180 66540 66181 66604
rect 66115 66539 66181 66540
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 65776 65968 65792
rect 66118 64290 66178 66539
rect 66308 66400 66628 67320
rect 66308 66336 66316 66400
rect 66380 66336 66396 66400
rect 66460 66336 66476 66400
rect 66540 66336 66556 66400
rect 66620 66336 66628 66400
rect 66308 65650 66628 66336
rect 71083 66332 71149 66333
rect 71083 66268 71084 66332
rect 71148 66268 71149 66332
rect 71083 66267 71149 66268
rect 71086 64290 71146 66267
rect 73475 65516 73541 65517
rect 73475 65452 73476 65516
rect 73540 65452 73541 65516
rect 73475 65451 73541 65452
rect 66029 64230 66178 64290
rect 71021 64230 71146 64290
rect 73478 64290 73538 65451
rect 86174 64290 86234 67627
rect 96368 66944 96688 67968
rect 96368 66880 96376 66944
rect 96440 66896 96456 66944
rect 96520 66896 96536 66944
rect 96600 66896 96616 66944
rect 96680 66880 96688 66944
rect 96368 66660 96410 66880
rect 96646 66660 96688 66880
rect 87275 66332 87341 66333
rect 87275 66268 87276 66332
rect 87340 66268 87341 66332
rect 87275 66267 87341 66268
rect 73478 64230 73577 64290
rect 66029 63676 66089 64230
rect 68522 64156 68588 64157
rect 68522 64092 68523 64156
rect 68587 64092 68588 64156
rect 68522 64091 68588 64092
rect 68525 63676 68585 64091
rect 71021 63676 71081 64230
rect 73517 63676 73577 64230
rect 86144 64230 86234 64290
rect 87278 64290 87338 66267
rect 96368 65856 96688 66660
rect 96368 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96688 65856
rect 96368 65650 96688 65792
rect 97028 67556 97348 68064
rect 97028 67488 97070 67556
rect 97306 67488 97348 67556
rect 97028 67424 97036 67488
rect 97340 67424 97348 67488
rect 97028 67320 97070 67424
rect 97306 67320 97348 67424
rect 105916 68032 106236 69056
rect 105916 67968 105924 68032
rect 105988 67968 106004 68032
rect 106068 67968 106084 68032
rect 106148 67968 106164 68032
rect 106228 67968 106236 68032
rect 105916 67408 106236 67968
rect 106652 126240 106972 126800
rect 106652 126176 106660 126240
rect 106724 126176 106740 126240
rect 106804 126176 106820 126240
rect 106884 126176 106900 126240
rect 106964 126176 106972 126240
rect 106652 125152 106972 126176
rect 106652 125088 106660 125152
rect 106724 125088 106740 125152
rect 106804 125088 106820 125152
rect 106884 125088 106900 125152
rect 106964 125088 106972 125152
rect 106652 124064 106972 125088
rect 106652 124000 106660 124064
rect 106724 124000 106740 124064
rect 106804 124000 106820 124064
rect 106884 124000 106900 124064
rect 106964 124000 106972 124064
rect 106652 122976 106972 124000
rect 106652 122912 106660 122976
rect 106724 122912 106740 122976
rect 106804 122912 106820 122976
rect 106884 122912 106900 122976
rect 106964 122912 106972 122976
rect 106652 121888 106972 122912
rect 106652 121824 106660 121888
rect 106724 121824 106740 121888
rect 106804 121824 106820 121888
rect 106884 121824 106900 121888
rect 106964 121824 106972 121888
rect 106652 120800 106972 121824
rect 106652 120736 106660 120800
rect 106724 120736 106740 120800
rect 106804 120736 106820 120800
rect 106884 120736 106900 120800
rect 106964 120736 106972 120800
rect 106652 119712 106972 120736
rect 106652 119648 106660 119712
rect 106724 119648 106740 119712
rect 106804 119648 106820 119712
rect 106884 119648 106900 119712
rect 106964 119648 106972 119712
rect 106652 118624 106972 119648
rect 106652 118560 106660 118624
rect 106724 118560 106740 118624
rect 106804 118560 106820 118624
rect 106884 118560 106900 118624
rect 106964 118560 106972 118624
rect 106652 117536 106972 118560
rect 106652 117472 106660 117536
rect 106724 117472 106740 117536
rect 106804 117472 106820 117536
rect 106884 117472 106900 117536
rect 106964 117472 106972 117536
rect 106652 116448 106972 117472
rect 106652 116384 106660 116448
rect 106724 116384 106740 116448
rect 106804 116384 106820 116448
rect 106884 116384 106900 116448
rect 106964 116384 106972 116448
rect 106652 115360 106972 116384
rect 106652 115296 106660 115360
rect 106724 115296 106740 115360
rect 106804 115296 106820 115360
rect 106884 115296 106900 115360
rect 106964 115296 106972 115360
rect 106652 114272 106972 115296
rect 106652 114208 106660 114272
rect 106724 114208 106740 114272
rect 106804 114208 106820 114272
rect 106884 114208 106900 114272
rect 106964 114208 106972 114272
rect 106652 113184 106972 114208
rect 106652 113120 106660 113184
rect 106724 113120 106740 113184
rect 106804 113120 106820 113184
rect 106884 113120 106900 113184
rect 106964 113120 106972 113184
rect 106652 112096 106972 113120
rect 106652 112032 106660 112096
rect 106724 112032 106740 112096
rect 106804 112032 106820 112096
rect 106884 112032 106900 112096
rect 106964 112032 106972 112096
rect 106652 111008 106972 112032
rect 106652 110944 106660 111008
rect 106724 110944 106740 111008
rect 106804 110944 106820 111008
rect 106884 110944 106900 111008
rect 106964 110944 106972 111008
rect 106652 109920 106972 110944
rect 106652 109856 106660 109920
rect 106724 109856 106740 109920
rect 106804 109856 106820 109920
rect 106884 109856 106900 109920
rect 106964 109856 106972 109920
rect 106652 108832 106972 109856
rect 106652 108768 106660 108832
rect 106724 108768 106740 108832
rect 106804 108768 106820 108832
rect 106884 108768 106900 108832
rect 106964 108768 106972 108832
rect 106652 107744 106972 108768
rect 106652 107680 106660 107744
rect 106724 107680 106740 107744
rect 106804 107680 106820 107744
rect 106884 107680 106900 107744
rect 106964 107680 106972 107744
rect 106652 106656 106972 107680
rect 106652 106592 106660 106656
rect 106724 106592 106740 106656
rect 106804 106592 106820 106656
rect 106884 106592 106900 106656
rect 106964 106592 106972 106656
rect 106652 105568 106972 106592
rect 106652 105504 106660 105568
rect 106724 105504 106740 105568
rect 106804 105504 106820 105568
rect 106884 105504 106900 105568
rect 106964 105504 106972 105568
rect 106652 104480 106972 105504
rect 106652 104416 106660 104480
rect 106724 104416 106740 104480
rect 106804 104416 106820 104480
rect 106884 104416 106900 104480
rect 106964 104416 106972 104480
rect 106652 103392 106972 104416
rect 106652 103328 106660 103392
rect 106724 103328 106740 103392
rect 106804 103328 106820 103392
rect 106884 103328 106900 103392
rect 106964 103328 106972 103392
rect 106652 102304 106972 103328
rect 106652 102240 106660 102304
rect 106724 102240 106740 102304
rect 106804 102240 106820 102304
rect 106884 102240 106900 102304
rect 106964 102240 106972 102304
rect 106652 101216 106972 102240
rect 106652 101152 106660 101216
rect 106724 101152 106740 101216
rect 106804 101152 106820 101216
rect 106884 101152 106900 101216
rect 106964 101152 106972 101216
rect 106652 100128 106972 101152
rect 106652 100064 106660 100128
rect 106724 100064 106740 100128
rect 106804 100064 106820 100128
rect 106884 100064 106900 100128
rect 106964 100064 106972 100128
rect 106652 99040 106972 100064
rect 106652 98976 106660 99040
rect 106724 98976 106740 99040
rect 106804 98976 106820 99040
rect 106884 98976 106900 99040
rect 106964 98976 106972 99040
rect 106652 98192 106972 98976
rect 106652 97956 106694 98192
rect 106930 97956 106972 98192
rect 106652 97952 106972 97956
rect 106652 97888 106660 97952
rect 106724 97888 106740 97952
rect 106804 97888 106820 97952
rect 106884 97888 106900 97952
rect 106964 97888 106972 97952
rect 106652 96864 106972 97888
rect 106652 96800 106660 96864
rect 106724 96800 106740 96864
rect 106804 96800 106820 96864
rect 106884 96800 106900 96864
rect 106964 96800 106972 96864
rect 106652 95776 106972 96800
rect 106652 95712 106660 95776
rect 106724 95712 106740 95776
rect 106804 95712 106820 95776
rect 106884 95712 106900 95776
rect 106964 95712 106972 95776
rect 106652 94688 106972 95712
rect 106652 94624 106660 94688
rect 106724 94624 106740 94688
rect 106804 94624 106820 94688
rect 106884 94624 106900 94688
rect 106964 94624 106972 94688
rect 106652 93600 106972 94624
rect 106652 93536 106660 93600
rect 106724 93536 106740 93600
rect 106804 93536 106820 93600
rect 106884 93536 106900 93600
rect 106964 93536 106972 93600
rect 106652 92512 106972 93536
rect 106652 92448 106660 92512
rect 106724 92448 106740 92512
rect 106804 92448 106820 92512
rect 106884 92448 106900 92512
rect 106964 92448 106972 92512
rect 106652 91424 106972 92448
rect 106652 91360 106660 91424
rect 106724 91360 106740 91424
rect 106804 91360 106820 91424
rect 106884 91360 106900 91424
rect 106964 91360 106972 91424
rect 106652 90336 106972 91360
rect 106652 90272 106660 90336
rect 106724 90272 106740 90336
rect 106804 90272 106820 90336
rect 106884 90272 106900 90336
rect 106964 90272 106972 90336
rect 106652 89248 106972 90272
rect 106652 89184 106660 89248
rect 106724 89184 106740 89248
rect 106804 89184 106820 89248
rect 106884 89184 106900 89248
rect 106964 89184 106972 89248
rect 106652 88160 106972 89184
rect 106652 88096 106660 88160
rect 106724 88096 106740 88160
rect 106804 88096 106820 88160
rect 106884 88096 106900 88160
rect 106964 88096 106972 88160
rect 106652 87072 106972 88096
rect 106652 87008 106660 87072
rect 106724 87008 106740 87072
rect 106804 87008 106820 87072
rect 106884 87008 106900 87072
rect 106964 87008 106972 87072
rect 106652 85984 106972 87008
rect 106652 85920 106660 85984
rect 106724 85920 106740 85984
rect 106804 85920 106820 85984
rect 106884 85920 106900 85984
rect 106964 85920 106972 85984
rect 106652 84896 106972 85920
rect 106652 84832 106660 84896
rect 106724 84832 106740 84896
rect 106804 84832 106820 84896
rect 106884 84832 106900 84896
rect 106964 84832 106972 84896
rect 106652 83808 106972 84832
rect 106652 83744 106660 83808
rect 106724 83744 106740 83808
rect 106804 83744 106820 83808
rect 106884 83744 106900 83808
rect 106964 83744 106972 83808
rect 106652 82720 106972 83744
rect 106652 82656 106660 82720
rect 106724 82656 106740 82720
rect 106804 82656 106820 82720
rect 106884 82656 106900 82720
rect 106964 82656 106972 82720
rect 106652 81632 106972 82656
rect 106652 81568 106660 81632
rect 106724 81568 106740 81632
rect 106804 81568 106820 81632
rect 106884 81568 106900 81632
rect 106964 81568 106972 81632
rect 106652 80544 106972 81568
rect 106652 80480 106660 80544
rect 106724 80480 106740 80544
rect 106804 80480 106820 80544
rect 106884 80480 106900 80544
rect 106964 80480 106972 80544
rect 106652 79456 106972 80480
rect 106652 79392 106660 79456
rect 106724 79392 106740 79456
rect 106804 79392 106820 79456
rect 106884 79392 106900 79456
rect 106964 79392 106972 79456
rect 106652 78368 106972 79392
rect 106652 78304 106660 78368
rect 106724 78304 106740 78368
rect 106804 78304 106820 78368
rect 106884 78304 106900 78368
rect 106964 78304 106972 78368
rect 106652 77280 106972 78304
rect 106652 77216 106660 77280
rect 106724 77216 106740 77280
rect 106804 77216 106820 77280
rect 106884 77216 106900 77280
rect 106964 77216 106972 77280
rect 106652 76192 106972 77216
rect 106652 76128 106660 76192
rect 106724 76128 106740 76192
rect 106804 76128 106820 76192
rect 106884 76128 106900 76192
rect 106964 76128 106972 76192
rect 106652 75104 106972 76128
rect 106652 75040 106660 75104
rect 106724 75040 106740 75104
rect 106804 75040 106820 75104
rect 106884 75040 106900 75104
rect 106964 75040 106972 75104
rect 106652 74016 106972 75040
rect 106652 73952 106660 74016
rect 106724 73952 106740 74016
rect 106804 73952 106820 74016
rect 106884 73952 106900 74016
rect 106964 73952 106972 74016
rect 106652 72928 106972 73952
rect 106652 72864 106660 72928
rect 106724 72864 106740 72928
rect 106804 72864 106820 72928
rect 106884 72864 106900 72928
rect 106964 72864 106972 72928
rect 106652 71840 106972 72864
rect 106652 71776 106660 71840
rect 106724 71776 106740 71840
rect 106804 71776 106820 71840
rect 106884 71776 106900 71840
rect 106964 71776 106972 71840
rect 106652 70752 106972 71776
rect 106652 70688 106660 70752
rect 106724 70688 106740 70752
rect 106804 70688 106820 70752
rect 106884 70688 106900 70752
rect 106964 70688 106972 70752
rect 106652 69664 106972 70688
rect 106652 69600 106660 69664
rect 106724 69600 106740 69664
rect 106804 69600 106820 69664
rect 106884 69600 106900 69664
rect 106964 69600 106972 69664
rect 106652 68576 106972 69600
rect 106652 68512 106660 68576
rect 106724 68512 106740 68576
rect 106804 68512 106820 68576
rect 106884 68512 106900 68576
rect 106964 68512 106972 68576
rect 106652 67488 106972 68512
rect 106652 67424 106660 67488
rect 106724 67424 106740 67488
rect 106804 67424 106820 67488
rect 106884 67424 106900 67488
rect 106964 67424 106972 67488
rect 106652 67408 106972 67424
rect 97028 66400 97348 67320
rect 97028 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97348 66400
rect 97028 65650 97348 66336
rect 105916 65856 106236 66416
rect 105916 65792 105924 65856
rect 105988 65792 106004 65856
rect 106068 65792 106084 65856
rect 106148 65792 106164 65856
rect 106228 65792 106236 65856
rect 105916 64768 106236 65792
rect 105916 64704 105924 64768
rect 105988 64704 106004 64768
rect 106068 64704 106084 64768
rect 106148 64704 106164 64768
rect 106228 64704 106236 64768
rect 87278 64230 87372 64290
rect 86144 63676 86204 64230
rect 87312 63676 87372 64230
rect 95857 63884 95923 63885
rect 95857 63820 95858 63884
rect 95922 63820 95923 63884
rect 95857 63819 95923 63820
rect 95860 63676 95920 63819
rect 105916 63680 106236 64704
rect 4868 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5188 63136
rect 4868 62048 5188 63072
rect 4868 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5188 62048
rect 4868 60960 5188 61984
rect 4868 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5188 60960
rect 4868 59872 5188 60896
rect 4868 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5188 59872
rect 4868 58784 5188 59808
rect 4868 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5188 58784
rect 4868 57696 5188 58720
rect 4868 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5188 57696
rect 4868 56608 5188 57632
rect 4868 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5188 56608
rect 4868 55520 5188 56544
rect 4868 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5188 55520
rect 4868 54432 5188 55456
rect 4868 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5188 54432
rect 4868 53344 5188 54368
rect 4868 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5188 53344
rect 4868 52256 5188 53280
rect 4868 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5188 52256
rect 4868 51168 5188 52192
rect 4868 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5188 51168
rect 4868 50080 5188 51104
rect 4868 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5188 50080
rect 4868 48992 5188 50016
rect 4868 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5188 48992
rect 4868 47904 5188 48928
rect 4868 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5188 47904
rect 4868 46816 5188 47840
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 105916 63616 105924 63680
rect 105988 63616 106004 63680
rect 106068 63616 106084 63680
rect 106148 63616 106164 63680
rect 106228 63616 106236 63680
rect 105916 62592 106236 63616
rect 105916 62528 105924 62592
rect 105988 62528 106004 62592
rect 106068 62528 106084 62592
rect 106148 62528 106164 62592
rect 106228 62528 106236 62592
rect 105916 61504 106236 62528
rect 105916 61440 105924 61504
rect 105988 61440 106004 61504
rect 106068 61440 106084 61504
rect 106148 61440 106164 61504
rect 106228 61440 106236 61504
rect 105916 60416 106236 61440
rect 105916 60352 105924 60416
rect 105988 60352 106004 60416
rect 106068 60352 106084 60416
rect 106148 60352 106164 60416
rect 106228 60352 106236 60416
rect 105916 59328 106236 60352
rect 105916 59264 105924 59328
rect 105988 59264 106004 59328
rect 106068 59264 106084 59328
rect 106148 59264 106164 59328
rect 106228 59264 106236 59328
rect 105916 58240 106236 59264
rect 105916 58176 105924 58240
rect 105988 58176 106004 58240
rect 106068 58176 106084 58240
rect 106148 58176 106164 58240
rect 106228 58176 106236 58240
rect 105916 57152 106236 58176
rect 105916 57088 105924 57152
rect 105988 57088 106004 57152
rect 106068 57088 106084 57152
rect 106148 57088 106164 57152
rect 106228 57088 106236 57152
rect 105916 56064 106236 57088
rect 105916 56000 105924 56064
rect 105988 56000 106004 56064
rect 106068 56000 106084 56064
rect 106148 56000 106164 56064
rect 106228 56000 106236 56064
rect 105916 54976 106236 56000
rect 105916 54912 105924 54976
rect 105988 54912 106004 54976
rect 106068 54912 106084 54976
rect 106148 54912 106164 54976
rect 106228 54912 106236 54976
rect 105916 53888 106236 54912
rect 105916 53824 105924 53888
rect 105988 53824 106004 53888
rect 106068 53824 106084 53888
rect 106148 53824 106164 53888
rect 106228 53824 106236 53888
rect 105916 52800 106236 53824
rect 105916 52736 105924 52800
rect 105988 52736 106004 52800
rect 106068 52736 106084 52800
rect 106148 52736 106164 52800
rect 106228 52736 106236 52800
rect 105916 51712 106236 52736
rect 105916 51648 105924 51712
rect 105988 51648 106004 51712
rect 106068 51648 106084 51712
rect 106148 51648 106164 51712
rect 106228 51648 106236 51712
rect 105916 50624 106236 51648
rect 105916 50560 105924 50624
rect 105988 50560 106004 50624
rect 106068 50560 106084 50624
rect 106148 50560 106164 50624
rect 106228 50560 106236 50624
rect 105916 49536 106236 50560
rect 105916 49472 105924 49536
rect 105988 49472 106004 49536
rect 106068 49472 106084 49536
rect 106148 49472 106164 49536
rect 106228 49472 106236 49536
rect 105916 48448 106236 49472
rect 105916 48384 105924 48448
rect 105988 48384 106004 48448
rect 106068 48384 106084 48448
rect 106148 48384 106164 48448
rect 106228 48384 106236 48448
rect 105916 47360 106236 48384
rect 105916 47296 105924 47360
rect 105988 47296 106004 47360
rect 106068 47296 106084 47360
rect 106148 47296 106164 47360
rect 106228 47296 106236 47360
rect 105916 46272 106236 47296
rect 105916 46208 105924 46272
rect 105988 46208 106004 46272
rect 106068 46208 106084 46272
rect 106148 46208 106164 46272
rect 106228 46208 106236 46272
rect 105916 45184 106236 46208
rect 105916 45120 105924 45184
rect 105988 45120 106004 45184
rect 106068 45120 106084 45184
rect 106148 45120 106164 45184
rect 106228 45120 106236 45184
rect 105916 44096 106236 45120
rect 105916 44032 105924 44096
rect 105988 44032 106004 44096
rect 106068 44032 106084 44096
rect 106148 44032 106164 44096
rect 106228 44032 106236 44096
rect 105916 43008 106236 44032
rect 105916 42944 105924 43008
rect 105988 42944 106004 43008
rect 106068 42944 106084 43008
rect 106148 42944 106164 43008
rect 106228 42944 106236 43008
rect 105916 41920 106236 42944
rect 105916 41856 105924 41920
rect 105988 41856 106004 41920
rect 106068 41856 106084 41920
rect 106148 41856 106164 41920
rect 106228 41856 106236 41920
rect 105916 40832 106236 41856
rect 105916 40768 105924 40832
rect 105988 40768 106004 40832
rect 106068 40768 106084 40832
rect 106148 40768 106164 40832
rect 106228 40768 106236 40832
rect 105916 39744 106236 40768
rect 105916 39680 105924 39744
rect 105988 39680 106004 39744
rect 106068 39680 106084 39744
rect 106148 39680 106164 39744
rect 106228 39680 106236 39744
rect 105916 38656 106236 39680
rect 105916 38592 105924 38656
rect 105988 38592 106004 38656
rect 106068 38592 106084 38656
rect 106148 38592 106164 38656
rect 106228 38592 106236 38656
rect 105916 37568 106236 38592
rect 105916 37504 105924 37568
rect 105988 37504 106004 37568
rect 106068 37504 106084 37568
rect 106148 37504 106164 37568
rect 106228 37504 106236 37568
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 10696 36920 11044 36962
rect 10696 36684 10752 36920
rect 10988 36684 11044 36920
rect 10696 36642 11044 36684
rect 100936 36920 101284 36962
rect 100936 36684 100992 36920
rect 101228 36684 101284 36920
rect 100936 36642 101284 36684
rect 105916 36480 106236 37504
rect 105916 36416 105924 36480
rect 105988 36416 106004 36480
rect 106068 36416 106084 36480
rect 106148 36416 106164 36480
rect 106228 36416 106236 36480
rect 10000 36260 10348 36302
rect 10000 36024 10056 36260
rect 10292 36024 10348 36260
rect 10000 35982 10348 36024
rect 101632 36260 101980 36302
rect 101632 36024 101688 36260
rect 101924 36024 101980 36260
rect 101632 35982 101980 36024
rect 105916 36260 106236 36416
rect 105916 36024 105958 36260
rect 106194 36024 106236 36260
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 105916 35392 106236 36024
rect 105916 35328 105924 35392
rect 105988 35328 106004 35392
rect 106068 35328 106084 35392
rect 106148 35328 106164 35392
rect 106228 35328 106236 35392
rect 105916 34304 106236 35328
rect 105916 34240 105924 34304
rect 105988 34240 106004 34304
rect 106068 34240 106084 34304
rect 106148 34240 106164 34304
rect 106228 34240 106236 34304
rect 105916 33216 106236 34240
rect 105916 33152 105924 33216
rect 105988 33152 106004 33216
rect 106068 33152 106084 33216
rect 106148 33152 106164 33216
rect 106228 33152 106236 33216
rect 105916 32128 106236 33152
rect 105916 32064 105924 32128
rect 105988 32064 106004 32128
rect 106068 32064 106084 32128
rect 106148 32064 106164 32128
rect 106228 32064 106236 32128
rect 105916 31040 106236 32064
rect 105916 30976 105924 31040
rect 105988 30976 106004 31040
rect 106068 30976 106084 31040
rect 106148 30976 106164 31040
rect 106228 30976 106236 31040
rect 105916 29952 106236 30976
rect 105916 29888 105924 29952
rect 105988 29888 106004 29952
rect 106068 29888 106084 29952
rect 106148 29888 106164 29952
rect 106228 29888 106236 29952
rect 105916 28864 106236 29888
rect 105916 28800 105924 28864
rect 105988 28800 106004 28864
rect 106068 28800 106084 28864
rect 106148 28800 106164 28864
rect 106228 28800 106236 28864
rect 105916 27776 106236 28800
rect 105916 27712 105924 27776
rect 105988 27712 106004 27776
rect 106068 27712 106084 27776
rect 106148 27712 106164 27776
rect 106228 27712 106236 27776
rect 105916 26688 106236 27712
rect 105916 26624 105924 26688
rect 105988 26624 106004 26688
rect 106068 26624 106084 26688
rect 106148 26624 106164 26688
rect 106228 26624 106236 26688
rect 105916 25600 106236 26624
rect 105916 25536 105924 25600
rect 105988 25536 106004 25600
rect 106068 25536 106084 25600
rect 106148 25536 106164 25600
rect 106228 25536 106236 25600
rect 105916 24512 106236 25536
rect 105916 24448 105924 24512
rect 105988 24448 106004 24512
rect 106068 24448 106084 24512
rect 106148 24448 106164 24512
rect 106228 24448 106236 24512
rect 105916 23424 106236 24448
rect 105916 23360 105924 23424
rect 105988 23360 106004 23424
rect 106068 23360 106084 23424
rect 106148 23360 106164 23424
rect 106228 23360 106236 23424
rect 105916 22336 106236 23360
rect 105916 22272 105924 22336
rect 105988 22272 106004 22336
rect 106068 22272 106084 22336
rect 106148 22272 106164 22336
rect 106228 22272 106236 22336
rect 105916 21248 106236 22272
rect 105916 21184 105924 21248
rect 105988 21184 106004 21248
rect 106068 21184 106084 21248
rect 106148 21184 106164 21248
rect 106228 21184 106236 21248
rect 105916 20160 106236 21184
rect 105916 20096 105924 20160
rect 105988 20096 106004 20160
rect 106068 20096 106084 20160
rect 106148 20096 106164 20160
rect 106228 20096 106236 20160
rect 105916 19072 106236 20096
rect 105916 19008 105924 19072
rect 105988 19008 106004 19072
rect 106068 19008 106084 19072
rect 106148 19008 106164 19072
rect 106228 19008 106236 19072
rect 105916 17984 106236 19008
rect 105916 17920 105924 17984
rect 105988 17920 106004 17984
rect 106068 17920 106084 17984
rect 106148 17920 106164 17984
rect 106228 17920 106236 17984
rect 105916 16896 106236 17920
rect 105916 16832 105924 16896
rect 105988 16832 106004 16896
rect 106068 16832 106084 16896
rect 106148 16832 106164 16896
rect 106228 16832 106236 16896
rect 105916 15808 106236 16832
rect 105916 15744 105924 15808
rect 105988 15744 106004 15808
rect 106068 15744 106084 15808
rect 106148 15744 106164 15808
rect 106228 15744 106236 15808
rect 105916 14720 106236 15744
rect 105916 14656 105924 14720
rect 105988 14656 106004 14720
rect 106068 14656 106084 14720
rect 106148 14656 106164 14720
rect 106228 14656 106236 14720
rect 105916 13632 106236 14656
rect 105916 13568 105924 13632
rect 105988 13568 106004 13632
rect 106068 13568 106084 13632
rect 106148 13568 106164 13632
rect 106228 13568 106236 13632
rect 105916 12544 106236 13568
rect 105916 12480 105924 12544
rect 105988 12480 106004 12544
rect 106068 12480 106084 12544
rect 106148 12480 106164 12544
rect 106228 12480 106236 12544
rect 105916 11456 106236 12480
rect 105916 11392 105924 11456
rect 105988 11392 106004 11456
rect 106068 11392 106084 11456
rect 106148 11392 106164 11456
rect 106228 11392 106236 11456
rect 105916 10368 106236 11392
rect 105916 10304 105924 10368
rect 105988 10304 106004 10368
rect 106068 10304 106084 10368
rect 106148 10304 106164 10368
rect 106228 10304 106236 10368
rect 16060 9893 16120 10038
rect 16057 9892 16123 9893
rect 16057 9828 16058 9892
rect 16122 9828 16123 9892
rect 16057 9827 16123 9828
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 23430 8261 23490 10038
rect 24626 9890 24686 10038
rect 25776 9890 25836 10038
rect 24626 9830 24778 9890
rect 25776 9830 25882 9890
rect 24718 8261 24778 9830
rect 25822 8261 25882 9830
rect 26926 8261 26986 10038
rect 28122 9890 28182 10038
rect 29280 9890 29340 10038
rect 30448 9890 30508 10038
rect 28122 9830 28274 9890
rect 29280 9830 29378 9890
rect 28214 8261 28274 9830
rect 29318 8261 29378 9830
rect 30422 9830 30508 9890
rect 31618 9890 31678 10038
rect 32784 9890 32844 10038
rect 33952 9890 34012 10038
rect 31618 9830 31770 9890
rect 32784 9830 32874 9890
rect 30422 8261 30482 9830
rect 31710 8261 31770 9830
rect 32814 8261 32874 9830
rect 33918 9830 34012 9890
rect 35120 9890 35180 10038
rect 36288 9890 36348 10038
rect 37456 9890 37516 10038
rect 35120 9830 35266 9890
rect 36288 9830 36370 9890
rect 33918 8261 33978 9830
rect 35206 8261 35266 9830
rect 36310 8261 36370 9830
rect 37414 9830 37516 9890
rect 38624 9890 38684 10038
rect 38624 9830 38762 9890
rect 37414 8261 37474 9830
rect 38702 8261 38762 9830
rect 23427 8260 23493 8261
rect 23427 8196 23428 8260
rect 23492 8196 23493 8260
rect 23427 8195 23493 8196
rect 24715 8260 24781 8261
rect 24715 8196 24716 8260
rect 24780 8196 24781 8260
rect 24715 8195 24781 8196
rect 25819 8260 25885 8261
rect 25819 8196 25820 8260
rect 25884 8196 25885 8260
rect 25819 8195 25885 8196
rect 26923 8260 26989 8261
rect 26923 8196 26924 8260
rect 26988 8196 26989 8260
rect 26923 8195 26989 8196
rect 28211 8260 28277 8261
rect 28211 8196 28212 8260
rect 28276 8196 28277 8260
rect 28211 8195 28277 8196
rect 29315 8260 29381 8261
rect 29315 8196 29316 8260
rect 29380 8196 29381 8260
rect 29315 8195 29381 8196
rect 30419 8260 30485 8261
rect 30419 8196 30420 8260
rect 30484 8196 30485 8260
rect 30419 8195 30485 8196
rect 31707 8260 31773 8261
rect 31707 8196 31708 8260
rect 31772 8196 31773 8260
rect 31707 8195 31773 8196
rect 32811 8260 32877 8261
rect 32811 8196 32812 8260
rect 32876 8196 32877 8260
rect 32811 8195 32877 8196
rect 33915 8260 33981 8261
rect 33915 8196 33916 8260
rect 33980 8196 33981 8260
rect 33915 8195 33981 8196
rect 35203 8260 35269 8261
rect 35203 8196 35204 8260
rect 35268 8196 35269 8260
rect 35203 8195 35269 8196
rect 36307 8260 36373 8261
rect 36307 8196 36308 8260
rect 36372 8196 36373 8260
rect 36307 8195 36373 8196
rect 37411 8260 37477 8261
rect 37411 8196 37412 8260
rect 37476 8196 37477 8260
rect 37411 8195 37477 8196
rect 38699 8260 38765 8261
rect 38699 8196 38700 8260
rect 38764 8196 38765 8260
rect 38699 8195 38765 8196
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 7104 35248 7880
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 7648 35908 8064
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 39806 4589 39866 10038
rect 40960 9890 41020 10038
rect 40910 9830 41020 9890
rect 42128 9890 42188 10038
rect 42128 9830 42258 9890
rect 40910 8261 40970 9830
rect 42198 8261 42258 9830
rect 43302 8261 43362 10038
rect 90529 9893 90589 10038
rect 90526 9892 90592 9893
rect 90526 9828 90527 9892
rect 90591 9828 90592 9892
rect 90526 9827 90592 9828
rect 90529 9210 90589 9827
rect 90682 9757 90742 10038
rect 90816 9890 90876 10038
rect 90955 9892 91021 9893
rect 90955 9890 90956 9892
rect 90816 9830 90956 9890
rect 90955 9828 90956 9830
rect 91020 9828 91021 9892
rect 90955 9827 91021 9828
rect 90679 9756 90745 9757
rect 90679 9692 90680 9756
rect 90744 9692 90745 9756
rect 90679 9691 90745 9692
rect 90529 9150 90650 9210
rect 90590 8261 90650 9150
rect 90958 8261 91018 9827
rect 105916 9280 106236 10304
rect 105916 9216 105924 9280
rect 105988 9216 106004 9280
rect 106068 9216 106084 9280
rect 106148 9216 106164 9280
rect 106228 9216 106236 9280
rect 40907 8260 40973 8261
rect 40907 8196 40908 8260
rect 40972 8196 40973 8260
rect 40907 8195 40973 8196
rect 42195 8260 42261 8261
rect 42195 8196 42196 8260
rect 42260 8196 42261 8260
rect 42195 8195 42261 8196
rect 43299 8260 43365 8261
rect 43299 8196 43300 8260
rect 43364 8196 43365 8260
rect 43299 8195 43365 8196
rect 90587 8260 90653 8261
rect 90587 8196 90588 8260
rect 90652 8196 90653 8260
rect 90587 8195 90653 8196
rect 90955 8260 91021 8261
rect 90955 8196 90956 8260
rect 91020 8196 91021 8260
rect 90955 8195 91021 8196
rect 105916 8192 106236 9216
rect 105916 8128 105924 8192
rect 105988 8128 106004 8192
rect 106068 8128 106084 8192
rect 106148 8128 106164 8192
rect 106228 8128 106236 8192
rect 65648 7104 65968 8064
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 5624 65968 5952
rect 65648 5388 65690 5624
rect 65926 5388 65968 5624
rect 65648 4928 65968 5388
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 39803 4588 39869 4589
rect 39803 4524 39804 4588
rect 39868 4524 39869 4588
rect 39803 4523 39869 4524
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
rect 66308 7648 66628 8064
rect 66308 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66628 7648
rect 66308 6560 66628 7584
rect 66308 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66628 6560
rect 66308 6284 66628 6496
rect 66308 6048 66350 6284
rect 66586 6048 66628 6284
rect 66308 5472 66628 6048
rect 66308 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66628 5472
rect 66308 4384 66628 5408
rect 66308 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66628 4384
rect 66308 3296 66628 4320
rect 66308 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66628 3296
rect 66308 2208 66628 3232
rect 66308 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66628 2208
rect 66308 2128 66628 2144
rect 96368 7104 96688 8064
rect 96368 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96688 7104
rect 96368 6016 96688 7040
rect 96368 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96688 6016
rect 96368 5624 96688 5952
rect 96368 5388 96410 5624
rect 96646 5388 96688 5624
rect 96368 4928 96688 5388
rect 96368 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96688 4928
rect 96368 3840 96688 4864
rect 96368 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96688 3840
rect 96368 2752 96688 3776
rect 96368 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96688 2752
rect 96368 2128 96688 2688
rect 97028 7648 97348 8064
rect 97028 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97348 7648
rect 97028 6560 97348 7584
rect 105916 7104 106236 8128
rect 105916 7040 105924 7104
rect 105988 7040 106004 7104
rect 106068 7040 106084 7104
rect 106148 7040 106164 7104
rect 106228 7040 106236 7104
rect 105916 7024 106236 7040
rect 106652 66400 106972 66416
rect 106652 66336 106660 66400
rect 106724 66336 106740 66400
rect 106804 66336 106820 66400
rect 106884 66336 106900 66400
rect 106964 66336 106972 66400
rect 106652 65312 106972 66336
rect 106652 65248 106660 65312
rect 106724 65248 106740 65312
rect 106804 65248 106820 65312
rect 106884 65248 106900 65312
rect 106964 65248 106972 65312
rect 106652 64224 106972 65248
rect 106652 64160 106660 64224
rect 106724 64160 106740 64224
rect 106804 64160 106820 64224
rect 106884 64160 106900 64224
rect 106964 64160 106972 64224
rect 106652 63136 106972 64160
rect 106652 63072 106660 63136
rect 106724 63072 106740 63136
rect 106804 63072 106820 63136
rect 106884 63072 106900 63136
rect 106964 63072 106972 63136
rect 106652 62048 106972 63072
rect 106652 61984 106660 62048
rect 106724 61984 106740 62048
rect 106804 61984 106820 62048
rect 106884 61984 106900 62048
rect 106964 61984 106972 62048
rect 106652 60960 106972 61984
rect 106652 60896 106660 60960
rect 106724 60896 106740 60960
rect 106804 60896 106820 60960
rect 106884 60896 106900 60960
rect 106964 60896 106972 60960
rect 106652 59872 106972 60896
rect 106652 59808 106660 59872
rect 106724 59808 106740 59872
rect 106804 59808 106820 59872
rect 106884 59808 106900 59872
rect 106964 59808 106972 59872
rect 106652 58784 106972 59808
rect 106652 58720 106660 58784
rect 106724 58720 106740 58784
rect 106804 58720 106820 58784
rect 106884 58720 106900 58784
rect 106964 58720 106972 58784
rect 106652 57696 106972 58720
rect 106652 57632 106660 57696
rect 106724 57632 106740 57696
rect 106804 57632 106820 57696
rect 106884 57632 106900 57696
rect 106964 57632 106972 57696
rect 106652 56608 106972 57632
rect 106652 56544 106660 56608
rect 106724 56544 106740 56608
rect 106804 56544 106820 56608
rect 106884 56544 106900 56608
rect 106964 56544 106972 56608
rect 106652 55520 106972 56544
rect 106652 55456 106660 55520
rect 106724 55456 106740 55520
rect 106804 55456 106820 55520
rect 106884 55456 106900 55520
rect 106964 55456 106972 55520
rect 106652 54432 106972 55456
rect 106652 54368 106660 54432
rect 106724 54368 106740 54432
rect 106804 54368 106820 54432
rect 106884 54368 106900 54432
rect 106964 54368 106972 54432
rect 106652 53344 106972 54368
rect 106652 53280 106660 53344
rect 106724 53280 106740 53344
rect 106804 53280 106820 53344
rect 106884 53280 106900 53344
rect 106964 53280 106972 53344
rect 106652 52256 106972 53280
rect 106652 52192 106660 52256
rect 106724 52192 106740 52256
rect 106804 52192 106820 52256
rect 106884 52192 106900 52256
rect 106964 52192 106972 52256
rect 106652 51168 106972 52192
rect 106652 51104 106660 51168
rect 106724 51104 106740 51168
rect 106804 51104 106820 51168
rect 106884 51104 106900 51168
rect 106964 51104 106972 51168
rect 106652 50080 106972 51104
rect 106652 50016 106660 50080
rect 106724 50016 106740 50080
rect 106804 50016 106820 50080
rect 106884 50016 106900 50080
rect 106964 50016 106972 50080
rect 106652 48992 106972 50016
rect 106652 48928 106660 48992
rect 106724 48928 106740 48992
rect 106804 48928 106820 48992
rect 106884 48928 106900 48992
rect 106964 48928 106972 48992
rect 106652 47904 106972 48928
rect 106652 47840 106660 47904
rect 106724 47840 106740 47904
rect 106804 47840 106820 47904
rect 106884 47840 106900 47904
rect 106964 47840 106972 47904
rect 106652 46816 106972 47840
rect 106652 46752 106660 46816
rect 106724 46752 106740 46816
rect 106804 46752 106820 46816
rect 106884 46752 106900 46816
rect 106964 46752 106972 46816
rect 106652 45728 106972 46752
rect 106652 45664 106660 45728
rect 106724 45664 106740 45728
rect 106804 45664 106820 45728
rect 106884 45664 106900 45728
rect 106964 45664 106972 45728
rect 106652 44640 106972 45664
rect 106652 44576 106660 44640
rect 106724 44576 106740 44640
rect 106804 44576 106820 44640
rect 106884 44576 106900 44640
rect 106964 44576 106972 44640
rect 106652 43552 106972 44576
rect 106652 43488 106660 43552
rect 106724 43488 106740 43552
rect 106804 43488 106820 43552
rect 106884 43488 106900 43552
rect 106964 43488 106972 43552
rect 106652 42464 106972 43488
rect 106652 42400 106660 42464
rect 106724 42400 106740 42464
rect 106804 42400 106820 42464
rect 106884 42400 106900 42464
rect 106964 42400 106972 42464
rect 106652 41376 106972 42400
rect 106652 41312 106660 41376
rect 106724 41312 106740 41376
rect 106804 41312 106820 41376
rect 106884 41312 106900 41376
rect 106964 41312 106972 41376
rect 106652 40288 106972 41312
rect 106652 40224 106660 40288
rect 106724 40224 106740 40288
rect 106804 40224 106820 40288
rect 106884 40224 106900 40288
rect 106964 40224 106972 40288
rect 106652 39200 106972 40224
rect 106652 39136 106660 39200
rect 106724 39136 106740 39200
rect 106804 39136 106820 39200
rect 106884 39136 106900 39200
rect 106964 39136 106972 39200
rect 106652 38112 106972 39136
rect 106652 38048 106660 38112
rect 106724 38048 106740 38112
rect 106804 38048 106820 38112
rect 106884 38048 106900 38112
rect 106964 38048 106972 38112
rect 106652 37024 106972 38048
rect 106652 36960 106660 37024
rect 106724 36960 106740 37024
rect 106804 36960 106820 37024
rect 106884 36960 106900 37024
rect 106964 36960 106972 37024
rect 106652 36920 106972 36960
rect 106652 36684 106694 36920
rect 106930 36684 106972 36920
rect 106652 35936 106972 36684
rect 106652 35872 106660 35936
rect 106724 35872 106740 35936
rect 106804 35872 106820 35936
rect 106884 35872 106900 35936
rect 106964 35872 106972 35936
rect 106652 34848 106972 35872
rect 106652 34784 106660 34848
rect 106724 34784 106740 34848
rect 106804 34784 106820 34848
rect 106884 34784 106900 34848
rect 106964 34784 106972 34848
rect 106652 33760 106972 34784
rect 106652 33696 106660 33760
rect 106724 33696 106740 33760
rect 106804 33696 106820 33760
rect 106884 33696 106900 33760
rect 106964 33696 106972 33760
rect 106652 32672 106972 33696
rect 106652 32608 106660 32672
rect 106724 32608 106740 32672
rect 106804 32608 106820 32672
rect 106884 32608 106900 32672
rect 106964 32608 106972 32672
rect 106652 31584 106972 32608
rect 106652 31520 106660 31584
rect 106724 31520 106740 31584
rect 106804 31520 106820 31584
rect 106884 31520 106900 31584
rect 106964 31520 106972 31584
rect 106652 30496 106972 31520
rect 106652 30432 106660 30496
rect 106724 30432 106740 30496
rect 106804 30432 106820 30496
rect 106884 30432 106900 30496
rect 106964 30432 106972 30496
rect 106652 29408 106972 30432
rect 106652 29344 106660 29408
rect 106724 29344 106740 29408
rect 106804 29344 106820 29408
rect 106884 29344 106900 29408
rect 106964 29344 106972 29408
rect 106652 28320 106972 29344
rect 106652 28256 106660 28320
rect 106724 28256 106740 28320
rect 106804 28256 106820 28320
rect 106884 28256 106900 28320
rect 106964 28256 106972 28320
rect 106652 27232 106972 28256
rect 106652 27168 106660 27232
rect 106724 27168 106740 27232
rect 106804 27168 106820 27232
rect 106884 27168 106900 27232
rect 106964 27168 106972 27232
rect 106652 26144 106972 27168
rect 106652 26080 106660 26144
rect 106724 26080 106740 26144
rect 106804 26080 106820 26144
rect 106884 26080 106900 26144
rect 106964 26080 106972 26144
rect 106652 25056 106972 26080
rect 106652 24992 106660 25056
rect 106724 24992 106740 25056
rect 106804 24992 106820 25056
rect 106884 24992 106900 25056
rect 106964 24992 106972 25056
rect 106652 23968 106972 24992
rect 106652 23904 106660 23968
rect 106724 23904 106740 23968
rect 106804 23904 106820 23968
rect 106884 23904 106900 23968
rect 106964 23904 106972 23968
rect 106652 22880 106972 23904
rect 106652 22816 106660 22880
rect 106724 22816 106740 22880
rect 106804 22816 106820 22880
rect 106884 22816 106900 22880
rect 106964 22816 106972 22880
rect 106652 21792 106972 22816
rect 106652 21728 106660 21792
rect 106724 21728 106740 21792
rect 106804 21728 106820 21792
rect 106884 21728 106900 21792
rect 106964 21728 106972 21792
rect 106652 20704 106972 21728
rect 106652 20640 106660 20704
rect 106724 20640 106740 20704
rect 106804 20640 106820 20704
rect 106884 20640 106900 20704
rect 106964 20640 106972 20704
rect 106652 19616 106972 20640
rect 106652 19552 106660 19616
rect 106724 19552 106740 19616
rect 106804 19552 106820 19616
rect 106884 19552 106900 19616
rect 106964 19552 106972 19616
rect 106652 18528 106972 19552
rect 106652 18464 106660 18528
rect 106724 18464 106740 18528
rect 106804 18464 106820 18528
rect 106884 18464 106900 18528
rect 106964 18464 106972 18528
rect 106652 17440 106972 18464
rect 106652 17376 106660 17440
rect 106724 17376 106740 17440
rect 106804 17376 106820 17440
rect 106884 17376 106900 17440
rect 106964 17376 106972 17440
rect 106652 16352 106972 17376
rect 106652 16288 106660 16352
rect 106724 16288 106740 16352
rect 106804 16288 106820 16352
rect 106884 16288 106900 16352
rect 106964 16288 106972 16352
rect 106652 15264 106972 16288
rect 106652 15200 106660 15264
rect 106724 15200 106740 15264
rect 106804 15200 106820 15264
rect 106884 15200 106900 15264
rect 106964 15200 106972 15264
rect 106652 14176 106972 15200
rect 106652 14112 106660 14176
rect 106724 14112 106740 14176
rect 106804 14112 106820 14176
rect 106884 14112 106900 14176
rect 106964 14112 106972 14176
rect 106652 13088 106972 14112
rect 106652 13024 106660 13088
rect 106724 13024 106740 13088
rect 106804 13024 106820 13088
rect 106884 13024 106900 13088
rect 106964 13024 106972 13088
rect 106652 12000 106972 13024
rect 106652 11936 106660 12000
rect 106724 11936 106740 12000
rect 106804 11936 106820 12000
rect 106884 11936 106900 12000
rect 106964 11936 106972 12000
rect 106652 10912 106972 11936
rect 106652 10848 106660 10912
rect 106724 10848 106740 10912
rect 106804 10848 106820 10912
rect 106884 10848 106900 10912
rect 106964 10848 106972 10912
rect 106652 9824 106972 10848
rect 106652 9760 106660 9824
rect 106724 9760 106740 9824
rect 106804 9760 106820 9824
rect 106884 9760 106900 9824
rect 106964 9760 106972 9824
rect 106652 8736 106972 9760
rect 106652 8672 106660 8736
rect 106724 8672 106740 8736
rect 106804 8672 106820 8736
rect 106884 8672 106900 8736
rect 106964 8672 106972 8736
rect 106652 7648 106972 8672
rect 106652 7584 106660 7648
rect 106724 7584 106740 7648
rect 106804 7584 106820 7648
rect 106884 7584 106900 7648
rect 106964 7584 106972 7648
rect 106652 7024 106972 7584
rect 97028 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97348 6560
rect 97028 6284 97348 6496
rect 97028 6048 97070 6284
rect 97306 6048 97348 6284
rect 97028 5472 97348 6048
rect 97028 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97348 5472
rect 97028 4384 97348 5408
rect 97028 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97348 4384
rect 97028 3296 97348 4320
rect 97028 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97348 3296
rect 97028 2208 97348 3232
rect 97028 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97348 2208
rect 97028 2128 97348 2144
<< via4 >>
rect 4250 126022 4486 126258
rect 4250 97408 4486 97532
rect 4250 97344 4280 97408
rect 4280 97344 4296 97408
rect 4296 97344 4360 97408
rect 4360 97344 4376 97408
rect 4376 97344 4440 97408
rect 4440 97344 4456 97408
rect 4456 97344 4486 97408
rect 4250 97296 4486 97344
rect 4250 66880 4280 66896
rect 4280 66880 4296 66896
rect 4296 66880 4360 66896
rect 4360 66880 4376 66896
rect 4376 66880 4440 66896
rect 4440 66880 4456 66896
rect 4456 66880 4486 66896
rect 4250 66660 4486 66880
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 126702 5146 126938
rect 34970 126022 35206 126258
rect 35630 126702 35866 126938
rect 65690 126022 65926 126258
rect 66350 126702 66586 126938
rect 96410 126022 96646 126258
rect 97070 126702 97306 126938
rect 105958 126022 106194 126258
rect 4910 97956 5146 98192
rect 10752 97956 10988 98192
rect 100992 97956 101228 98192
rect 10056 97296 10292 97532
rect 101688 97296 101924 97532
rect 105958 97408 106194 97532
rect 105958 97344 105988 97408
rect 105988 97344 106004 97408
rect 106004 97344 106068 97408
rect 106068 97344 106084 97408
rect 106084 97344 106148 97408
rect 106148 97344 106164 97408
rect 106164 97344 106194 97408
rect 105958 97296 106194 97344
rect 4910 67488 5146 67556
rect 4910 67424 4940 67488
rect 4940 67424 4956 67488
rect 4956 67424 5020 67488
rect 5020 67424 5036 67488
rect 5036 67424 5100 67488
rect 5100 67424 5116 67488
rect 5116 67424 5146 67488
rect 4910 67320 5146 67424
rect 34970 66880 35000 66896
rect 35000 66880 35016 66896
rect 35016 66880 35080 66896
rect 35080 66880 35096 66896
rect 35096 66880 35160 66896
rect 35160 66880 35176 66896
rect 35176 66880 35206 66896
rect 34970 66660 35206 66880
rect 35630 67488 35866 67556
rect 35630 67424 35660 67488
rect 35660 67424 35676 67488
rect 35676 67424 35740 67488
rect 35740 67424 35756 67488
rect 35756 67424 35820 67488
rect 35820 67424 35836 67488
rect 35836 67424 35866 67488
rect 35630 67320 35866 67424
rect 65690 66880 65720 66896
rect 65720 66880 65736 66896
rect 65736 66880 65800 66896
rect 65800 66880 65816 66896
rect 65816 66880 65880 66896
rect 65880 66880 65896 66896
rect 65896 66880 65926 66896
rect 65690 66660 65926 66880
rect 66350 67488 66586 67556
rect 66350 67424 66380 67488
rect 66380 67424 66396 67488
rect 66396 67424 66460 67488
rect 66460 67424 66476 67488
rect 66476 67424 66540 67488
rect 66540 67424 66556 67488
rect 66556 67424 66586 67488
rect 66350 67320 66586 67424
rect 96410 66880 96440 66896
rect 96440 66880 96456 66896
rect 96456 66880 96520 66896
rect 96520 66880 96536 66896
rect 96536 66880 96600 66896
rect 96600 66880 96616 66896
rect 96616 66880 96646 66896
rect 96410 66660 96646 66880
rect 97070 67488 97306 67556
rect 97070 67424 97100 67488
rect 97100 67424 97116 67488
rect 97116 67424 97180 67488
rect 97180 67424 97196 67488
rect 97196 67424 97260 67488
rect 97260 67424 97276 67488
rect 97276 67424 97306 67488
rect 97070 67320 97306 67424
rect 106694 97956 106930 98192
rect 4910 36684 5146 36920
rect 10752 36684 10988 36920
rect 100992 36684 101228 36920
rect 10056 36024 10292 36260
rect 101688 36024 101924 36260
rect 105958 36024 106194 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 6048 35866 6284
rect 65690 5388 65926 5624
rect 66350 6048 66586 6284
rect 96410 5388 96646 5624
rect 106694 36684 106930 36920
rect 97070 6048 97306 6284
<< metal5 >>
rect 4208 126938 108884 126980
rect 4208 126702 4910 126938
rect 5146 126702 35630 126938
rect 35866 126702 66350 126938
rect 66586 126702 97070 126938
rect 97306 126702 108884 126938
rect 4208 126660 108884 126702
rect 4208 126258 108884 126300
rect 4208 126022 4250 126258
rect 4486 126022 34970 126258
rect 35206 126022 65690 126258
rect 65926 126022 96410 126258
rect 96646 126022 105958 126258
rect 106194 126022 108884 126258
rect 4208 125980 108884 126022
rect 1056 98192 108884 98234
rect 1056 97956 4910 98192
rect 5146 97956 10752 98192
rect 10988 97956 100992 98192
rect 101228 97956 106694 98192
rect 106930 97956 108884 98192
rect 1056 97914 108884 97956
rect 1056 97532 108884 97574
rect 1056 97296 4250 97532
rect 4486 97296 10056 97532
rect 10292 97296 101688 97532
rect 101924 97296 105958 97532
rect 106194 97296 108884 97532
rect 1056 97254 108884 97296
rect 1056 67556 108884 67598
rect 1056 67320 4910 67556
rect 5146 67320 35630 67556
rect 35866 67320 66350 67556
rect 66586 67320 97070 67556
rect 97306 67320 108884 67556
rect 1056 67278 108884 67320
rect 1056 66896 108884 66938
rect 1056 66660 4250 66896
rect 4486 66660 34970 66896
rect 35206 66660 65690 66896
rect 65926 66660 96410 66896
rect 96646 66660 108884 66896
rect 1056 66618 108884 66660
rect 1056 36920 108884 36962
rect 1056 36684 4910 36920
rect 5146 36684 10752 36920
rect 10988 36684 100992 36920
rect 101228 36684 106694 36920
rect 106930 36684 108884 36920
rect 1056 36642 108884 36684
rect 1056 36260 108884 36302
rect 1056 36024 4250 36260
rect 4486 36024 10056 36260
rect 10292 36024 101688 36260
rect 101924 36024 105958 36260
rect 106194 36024 108884 36260
rect 1056 35982 108884 36024
rect 1056 6284 108884 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 66350 6284
rect 66586 6048 97070 6284
rect 97306 6048 108884 6284
rect 1056 6006 108884 6048
rect 1056 5624 108884 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 65690 5624
rect 65926 5388 96410 5624
rect 96646 5388 108884 5624
rect 1056 5346 108884 5388
use sky130_fd_sc_hd__inv_2  _061_
timestamp 1
transform -1 0 93840 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1
transform -1 0 87584 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _063_
timestamp 1
transform 1 0 34960 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _064_
timestamp 1
transform 1 0 33120 0 1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _065_
timestamp 1
transform 1 0 38640 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _066_
timestamp 1
transform 1 0 33212 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _067_
timestamp 1
transform 1 0 39928 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _068_
timestamp 1
transform 1 0 46184 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _069_
timestamp 1
transform 1 0 43976 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _070_
timestamp 1
transform -1 0 69000 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _071_
timestamp 1
transform -1 0 67528 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _072_
timestamp 1
transform -1 0 70656 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _073_
timestamp 1
transform -1 0 72312 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _074_
timestamp 1
transform -1 0 71484 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _075_
timestamp 1
transform -1 0 69828 0 1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _076_
timestamp 1
transform -1 0 75900 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _077_
timestamp 1
transform -1 0 74152 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _078_
timestamp 1
transform -1 0 85928 0 1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _079_
timestamp 1
transform 1 0 104328 0 -1 85952
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _080_
timestamp 1
transform 1 0 90436 0 1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _081_
timestamp 1
transform 1 0 104328 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _082_
timestamp 1
transform -1 0 96232 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _083_
timestamp 1
transform 1 0 95404 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _084_
timestamp 1
transform 1 0 102028 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _085_
timestamp 1
transform -1 0 100464 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _086_
timestamp 1
transform 1 0 91356 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _087_
timestamp 1
transform 1 0 104328 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _088_
timestamp 1
transform 1 0 98348 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _089_
timestamp 1
transform 1 0 104328 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _090_
timestamp 1
transform -1 0 104972 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _091_
timestamp 1
transform 1 0 104328 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _092_
timestamp 1
transform 1 0 104328 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _093_
timestamp 1
transform -1 0 105064 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _094_
timestamp 1
transform 1 0 92368 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _095_
timestamp 1
transform -1 0 80040 0 1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1
transform -1 0 91908 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 1
transform -1 0 90160 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098_
timestamp 1
transform 1 0 90160 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1
transform 1 0 88044 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1
transform -1 0 86480 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1
transform 1 0 88228 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1
transform -1 0 95680 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1
transform 1 0 87124 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1
transform 1 0 104328 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105_
timestamp 1
transform 1 0 89056 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1
transform 1 0 105708 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp 1
transform 1 0 87676 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1
transform 1 0 93932 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _109_
timestamp 1
transform -1 0 105156 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp 1
transform 1 0 88780 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 1
transform 1 0 76176 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1
transform -1 0 17480 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113_
timestamp 1
transform -1 0 30728 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 1
transform -1 0 29164 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1
transform -1 0 30452 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 1
transform -1 0 29072 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 1
transform -1 0 33120 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1
transform -1 0 31188 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1
transform 1 0 76912 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _120_
timestamp 1
transform 1 0 82708 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _121_
timestamp 1
transform 1 0 86664 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _122_
timestamp 1
transform 1 0 86204 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _123_
timestamp 1
transform 1 0 83628 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _124_
timestamp 1
transform 1 0 89424 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _125_
timestamp 1
transform 1 0 88044 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _126_
timestamp 1
transform 1 0 94116 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _127_
timestamp 1
transform 1 0 91356 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _128_
timestamp 1
transform -1 0 91264 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _129_
timestamp 1
transform -1 0 106168 0 -1 76160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _130_
timestamp 1
transform 1 0 96508 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _131_
timestamp 1
transform -1 0 98992 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _132_
timestamp 1
transform 1 0 92000 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _133_
timestamp 1
transform -1 0 96416 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _134_
timestamp 1
transform -1 0 106168 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _135_
timestamp 1
transform 1 0 93196 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _136_
timestamp 1
transform -1 0 79396 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _137_
timestamp 1
transform -1 0 20700 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _138_
timestamp 1
transform 1 0 21988 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _139_
timestamp 1
transform -1 0 25116 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _140_
timestamp 1
transform 1 0 24380 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _141_
timestamp 1
transform -1 0 22264 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _142_
timestamp 1
transform -1 0 28888 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _143_
timestamp 1
transform -1 0 31924 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _144_
timestamp 1
transform 1 0 85284 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform 1 0 86480 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform -1 0 72496 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform 1 0 69644 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform -1 0 85100 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform -1 0 33212 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform 1 0 66516 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform 1 0 69460 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform -1 0 21988 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1
transform 1 0 95220 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A1
timestamp 1
transform -1 0 35972 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__S
timestamp 1
transform 1 0 35972 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A1
timestamp 1
transform 1 0 33948 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__S
timestamp 1
transform 1 0 34132 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A1
timestamp 1
transform -1 0 39652 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__S
timestamp 1
transform 1 0 39652 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A1
timestamp 1
transform -1 0 34224 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__S
timestamp 1
transform 1 0 34224 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A1
timestamp 1
transform -1 0 41124 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__S
timestamp 1
transform 1 0 41124 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__X
timestamp 1
transform -1 0 40940 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A1
timestamp 1
transform -1 0 47380 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__S
timestamp 1
transform 1 0 47564 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__X
timestamp 1
transform -1 0 47196 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A1
timestamp 1
transform -1 0 44988 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__S
timestamp 1
transform 1 0 44988 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A0
timestamp 1
transform 1 0 67988 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A1
timestamp 1
transform -1 0 67988 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__S
timestamp 1
transform 1 0 68632 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A1
timestamp 1
transform -1 0 66516 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__S
timestamp 1
transform 1 0 67528 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A1
timestamp 1
transform 1 0 69644 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__S
timestamp 1
transform -1 0 69644 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A1
timestamp 1
transform -1 0 71484 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A1
timestamp 1
transform -1 0 70932 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A1
timestamp 1
transform 1 0 68816 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__X
timestamp 1
transform -1 0 70012 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A1
timestamp 1
transform -1 0 75072 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A1
timestamp 1
transform -1 0 73232 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__X
timestamp 1
transform 1 0 74152 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A1
timestamp 1
transform 1 0 84732 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__B
timestamp 1
transform -1 0 90252 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A1
timestamp 1
transform -1 0 104512 0 -1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__B1
timestamp 1
transform -1 0 104696 0 -1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__Y
timestamp 1
transform -1 0 105708 0 1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__B
timestamp 1
transform -1 0 96600 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__B
timestamp 1
transform 1 0 96876 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__X
timestamp 1
transform -1 0 96876 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1
transform 1 0 100464 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B
timestamp 1
transform 1 0 92184 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1
transform -1 0 104512 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__B
timestamp 1
transform 1 0 104328 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__C
timestamp 1
transform -1 0 104696 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A2
timestamp 1
transform 1 0 98716 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__B
timestamp 1
transform -1 0 104512 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1
transform 1 0 104328 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__B
timestamp 1
transform 1 0 104512 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__C
timestamp 1
transform -1 0 105248 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__X
timestamp 1
transform -1 0 105432 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A1
timestamp 1
transform 1 0 104328 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A2
timestamp 1
transform 1 0 104512 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A4
timestamp 1
transform 1 0 104696 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__B1
timestamp 1
transform 1 0 105064 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__X
timestamp 1
transform -1 0 105432 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A_N
timestamp 1
transform 1 0 92920 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__B
timestamp 1
transform -1 0 93564 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__B
timestamp 1
transform -1 0 80224 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1
transform 1 0 93380 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1
transform 1 0 96048 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1
transform 1 0 104604 0 -1 80512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1
transform 1 0 105524 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1
transform 1 0 94392 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1
transform -1 0 105340 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1
transform 1 0 76452 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1
transform 1 0 17480 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1
transform 1 0 30728 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1
transform 1 0 29532 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1
transform 1 0 30912 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1
transform -1 0 29256 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1
transform 1 0 32660 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1
transform 1 0 31188 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1
transform 1 0 77188 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__CLK
timestamp 1
transform -1 0 82708 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__Q
timestamp 1
transform 1 0 84548 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__CLK
timestamp 1
transform 1 0 88780 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__Q
timestamp 1
transform 1 0 88504 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__CLK
timestamp 1
transform 1 0 88504 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__Q
timestamp 1
transform -1 0 88504 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__CLK
timestamp 1
transform -1 0 83536 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__Q
timestamp 1
transform -1 0 85652 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__CLK
timestamp 1
transform 1 0 92000 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__D
timestamp 1
transform 1 0 89240 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__CLK
timestamp 1
transform 1 0 90804 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__Q
timestamp 1
transform -1 0 90620 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__CLK
timestamp 1
transform 1 0 96232 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__D
timestamp 1
transform -1 0 94392 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__CLK
timestamp 1
transform 1 0 93196 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__CLK
timestamp 1
transform 1 0 91264 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__CLK
timestamp 1
transform -1 0 106352 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__CLK
timestamp 1
transform -1 0 100188 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__CLK
timestamp 1
transform 1 0 99728 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__CLK
timestamp 1
transform 1 0 93932 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__CLK
timestamp 1
transform 1 0 96876 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__CLK
timestamp 1
transform -1 0 106352 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__CLK
timestamp 1
transform 1 0 95680 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__CLK
timestamp 1
transform -1 0 77556 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__CLK
timestamp 1
transform 1 0 20884 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__Q
timestamp 1
transform -1 0 20884 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__CLK
timestamp 1
transform 1 0 21528 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__Q
timestamp 1
transform -1 0 24012 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__CLK
timestamp 1
transform 1 0 23092 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__Q
timestamp 1
transform -1 0 25300 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__CLK
timestamp 1
transform 1 0 24104 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__Q
timestamp 1
transform -1 0 26404 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__CLK
timestamp 1
transform 1 0 20240 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__D
timestamp 1
transform -1 0 22448 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__Q
timestamp 1
transform -1 0 22632 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__CLK
timestamp 1
transform -1 0 29440 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__D
timestamp 1
transform -1 0 29072 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__Q
timestamp 1
transform -1 0 29900 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__CLK
timestamp 1
transform -1 0 32292 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__Q
timestamp 1
transform -1 0 32108 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__CLK
timestamp 1
transform -1 0 87768 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__Q
timestamp 1
transform 1 0 87400 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1
transform -1 0 62468 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 1
transform 1 0 62100 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_A
timestamp 1
transform 1 0 21252 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_X
timestamp 1
transform 1 0 21344 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_A
timestamp 1
transform 1 0 57868 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_X
timestamp 1
transform -1 0 58236 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_A
timestamp 1
transform -1 0 104512 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_X
timestamp 1
transform -1 0 106352 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_A
timestamp 1
transform -1 0 105064 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_X
timestamp 1
transform -1 0 106352 0 -1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload0_A
timestamp 1
transform 1 0 19228 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload1_A
timestamp 1
transform -1 0 57132 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload2_A
timestamp 1
transform 1 0 105064 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout84_X
timestamp 1
transform -1 0 70564 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout112_A
timestamp 1
transform 1 0 90620 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_A
timestamp 1
transform -1 0 105708 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_X
timestamp 1
transform -1 0 105524 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout114_X
timestamp 1
transform 1 0 105156 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1
transform -1 0 23276 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1
transform -1 0 24564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1
transform -1 0 1840 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1
transform -1 0 1840 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1
transform -1 0 1840 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1
transform -1 0 1840 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1
transform -1 0 1840 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1
transform -1 0 1840 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1
transform -1 0 2116 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_X
timestamp 1
transform -1 0 1932 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1
transform -1 0 2116 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_X
timestamp 1
transform 1 0 2300 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1
transform -1 0 1840 0 -1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1
transform -1 0 1840 0 1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1
transform -1 0 1840 0 1 96832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1
transform -1 0 1840 0 -1 99008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1
transform -1 0 1840 0 -1 100096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1
transform -1 0 1840 0 1 101184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1
transform -1 0 1840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1
transform -1 0 1840 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1
transform -1 0 25852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1
transform -1 0 37444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1
transform -1 0 38732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1
transform -1 0 40020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1
transform -1 0 41308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1
transform -1 0 41952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1
transform -1 0 43240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1
transform -1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1
transform -1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1
transform -1 0 29072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1
transform -1 0 30360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1
transform -1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1
transform -1 0 32936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1
transform -1 0 34224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1
transform -1 0 35512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1
transform -1 0 36156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1
transform -1 0 2116 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_X
timestamp 1
transform 1 0 1748 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1
transform -1 0 2116 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_X
timestamp 1
transform 1 0 1748 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1
transform -1 0 2116 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_X
timestamp 1
transform 1 0 1748 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1
transform -1 0 2116 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_X
timestamp 1
transform 1 0 1748 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1
transform -1 0 2116 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_X
timestamp 1
transform -1 0 1932 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1
transform -1 0 2116 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_X
timestamp 1
transform 1 0 1748 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1
transform -1 0 2116 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_X
timestamp 1
transform 1 0 1748 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1
transform -1 0 2116 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_X
timestamp 1
transform -1 0 1932 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1
transform -1 0 2116 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_X
timestamp 1
transform 1 0 1748 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1
transform -1 0 2116 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_X
timestamp 1
transform -1 0 1932 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1
transform -1 0 2116 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_X
timestamp 1
transform 1 0 1748 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1
transform -1 0 2116 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_X
timestamp 1
transform 1 0 1748 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1
transform -1 0 2116 0 -1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_X
timestamp 1
transform 1 0 1748 0 -1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1
transform -1 0 2300 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_X
timestamp 1
transform -1 0 1932 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1
transform -1 0 2116 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_X
timestamp 1
transform -1 0 1932 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1
transform -1 0 2116 0 1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_X
timestamp 1
transform -1 0 1932 0 1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1
transform -1 0 108284 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew86_A
timestamp 1
transform -1 0 105340 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew86_X
timestamp 1
transform -1 0 105524 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew87_X
timestamp 1
transform -1 0 96048 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew88_X
timestamp 1
transform -1 0 105064 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew90_X
timestamp 1
transform -1 0 104880 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew91_A
timestamp 1
transform -1 0 104880 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew91_X
timestamp 1
transform -1 0 105064 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew92_X
timestamp 1
transform -1 0 99636 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew94_A
timestamp 1
transform -1 0 105340 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew94_X
timestamp 1
transform -1 0 105524 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew95_X
timestamp 1
transform 1 0 100648 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew98_X
timestamp 1
transform -1 0 102488 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew101_A
timestamp 1
transform -1 0 105064 0 -1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew102_X
timestamp 1
transform 1 0 97060 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew103_X
timestamp 1
transform -1 0 99820 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew104_X
timestamp 1
transform -1 0 104880 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew106_A
timestamp 1
transform -1 0 91632 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew107_X
timestamp 1
transform -1 0 104788 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew108_X
timestamp 1
transform -1 0 104880 0 1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew109_A
timestamp 1
transform -1 0 104880 0 -1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew110_X
timestamp 1
transform 1 0 96508 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[2]
timestamp 1
transform -1 0 104512 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[3]
timestamp 1
transform -1 0 104512 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[4]
timestamp 1
transform 1 0 104328 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[5]
timestamp 1
transform -1 0 90712 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[6]
timestamp 1
transform -1 0 90896 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[7]
timestamp 1
transform -1 0 91080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_clk0
timestamp 1
transform -1 0 16284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_clk1
timestamp 1
transform 1 0 96232 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[7]
timestamp 1
transform 1 0 53544 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr0[0]
timestamp 1
transform -1 0 23644 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr0[1]
timestamp 1
transform -1 0 24840 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[0]
timestamp 1
transform -1 0 87492 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[1]
timestamp 1
transform -1 0 86388 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[6]
timestamp 1
transform -1 0 90436 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_clk0
timestamp 1
transform 1 0 16100 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_clk1
timestamp 1
transform -1 0 96048 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[0]
timestamp 1
transform -1 0 26036 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[1]
timestamp 1
transform -1 0 27140 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[2]
timestamp 1
transform -1 0 28336 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[3]
timestamp 1
transform -1 0 29716 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[4]
timestamp 1
transform -1 0 30636 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[5]
timestamp 1
transform -1 0 31832 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[6]
timestamp 1
transform -1 0 33028 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[7]
timestamp 1
transform -1 0 34132 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[8]
timestamp 1
transform -1 0 35328 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[9]
timestamp 1
transform -1 0 36524 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[10]
timestamp 1
transform -1 0 37628 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[11]
timestamp 1
transform -1 0 38824 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[12]
timestamp 1
transform -1 0 40020 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[13]
timestamp 1
transform -1 0 41216 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[14]
timestamp 1
transform -1 0 42320 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[15]
timestamp 1
transform -1 0 43516 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output52_A
timestamp 1
transform -1 0 1840 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output53_A
timestamp 1
transform 1 0 108100 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1
transform -1 0 108284 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1
transform 1 0 108100 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output59_A
timestamp 1
transform 1 0 1656 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output60_A
timestamp 1
transform 1 0 1656 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output61_A
timestamp 1
transform -1 0 1840 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output62_A
timestamp 1
transform -1 0 1840 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output63_A
timestamp 1
transform 1 0 1656 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1
transform 1 0 1656 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output65_A
timestamp 1
transform -1 0 108284 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 1
transform 1 0 108100 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output67_A
timestamp 1
transform -1 0 108284 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire68_X
timestamp 1
transform -1 0 62284 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire69_X
timestamp 1
transform -1 0 59800 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire70_X
timestamp 1
transform -1 0 58880 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire71_X
timestamp 1
transform -1 0 50048 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire72_X
timestamp 1
transform -1 0 48852 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire73_X
timestamp 1
transform -1 0 45540 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire74_X
timestamp 1
transform -1 0 41952 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire75_X
timestamp 1
transform -1 0 41768 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire76_X
timestamp 1
transform -1 0 38088 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire77_X
timestamp 1
transform -1 0 77740 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire78_X
timestamp 1
transform -1 0 71852 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire79_X
timestamp 1
transform -1 0 70932 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire80_X
timestamp 1
transform -1 0 67160 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire81_X
timestamp 1
transform -1 0 66148 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire82_X
timestamp 1
transform -1 0 64400 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire83_X
timestamp 1
transform -1 0 36524 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform -1 0 62100 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1
transform -1 0 21252 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1
transform 1 0 55936 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1
transform 1 0 104328 0 -1 58752
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1
transform 1 0 104328 0 -1 78336
box -38 -48 1878 592
use sky130_fd_sc_hd__bufinv_8  clkload0
timestamp 1
transform 1 0 17848 0 -1 66368
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_8  clkload1
timestamp 1
transform 1 0 56120 0 1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__clkinvlp_4  clkload2
timestamp 1
transform 1 0 104328 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout84
timestamp 1
transform -1 0 70380 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout85
timestamp 1
transform -1 0 79396 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout112
timestamp 1
transform -1 0 89424 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout113
timestamp 1
transform 1 0 104328 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout114
timestamp 1
transform -1 0 105156 0 1 44608
box -38 -48 866 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_237
timestamp 1
transform 1 0 22908 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244
timestamp 1
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_258
timestamp 1
transform 1 0 24840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_266
timestamp 1
transform 1 0 25576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_286
timestamp 1
transform 1 0 27416 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_294
timestamp 1
transform 1 0 28152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_300
timestamp 1
transform 1 0 28704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309
timestamp 1
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_315
timestamp 1
transform 1 0 30084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_321
timestamp 1
transform 1 0 30636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_329
timestamp 1
transform 1 0 31372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_343
timestamp 1
transform 1 0 32660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_349
timestamp 1
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_357
timestamp 1
transform 1 0 33948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_365
timestamp 1
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_371
timestamp 1
transform 1 0 35236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_377
timestamp 1
transform 1 0 35788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_398
timestamp 1
transform 1 0 37720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_406
timestamp 1
transform 1 0 38456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_426
timestamp 1
transform 1 0 40296 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_434
timestamp 1
transform 1 0 41032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_440
timestamp 1
transform 1 0 41584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_449
timestamp 1
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_455
timestamp 1
transform 1 0 42964 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1636968456
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1636968456
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1636968456
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1636968456
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1636968456
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1636968456
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1636968456
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1636968456
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1636968456
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1636968456
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1636968456
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_617
timestamp 1636968456
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_629
timestamp 1636968456
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1636968456
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1636968456
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1636968456
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_685
timestamp 1636968456
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1636968456
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1636968456
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1636968456
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1636968456
transform 1 0 69276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1636968456
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1636968456
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1636968456
transform 1 0 73324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_797
timestamp 1636968456
transform 1 0 74428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 1
transform 1 0 75532 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1636968456
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1636968456
transform 1 0 77004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1
transform 1 0 78108 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1636968456
transform 1 0 78476 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1636968456
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1636968456
transform 1 0 81052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1636968456
transform 1 0 82156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 1
transform 1 0 83260 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1636968456
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1636968456
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1636968456
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1636968456
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1636968456
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1636968456
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1636968456
transform 1 0 91356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1636968456
transform 1 0 92460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1009
timestamp 1636968456
transform 1 0 93932 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1021
timestamp 1636968456
transform 1 0 95036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1037
timestamp 1636968456
transform 1 0 96508 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1049
timestamp 1636968456
transform 1 0 97612 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1061
timestamp 1
transform 1 0 98716 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1636968456
transform 1 0 99084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1636968456
transform 1 0 100188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1636968456
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1105
timestamp 1636968456
transform 1 0 102764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1121
timestamp 1636968456
transform 1 0 104236 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1133
timestamp 1636968456
transform 1 0 105340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1149
timestamp 1636968456
transform 1 0 106812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1161
timestamp 1
transform 1 0 107916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1167
timestamp 1
transform 1 0 108468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636968456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636968456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636968456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636968456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636968456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636968456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636968456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636968456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636968456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636968456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636968456
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636968456
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636968456
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636968456
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636968456
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636968456
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636968456
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636968456
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636968456
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636968456
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636968456
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636968456
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636968456
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636968456
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1636968456
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1636968456
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1636968456
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1636968456
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1636968456
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1636968456
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1636968456
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1636968456
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1636968456
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1636968456
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1636968456
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1636968456
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1636968456
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1636968456
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1636968456
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1636968456
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 1
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1636968456
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1636968456
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1636968456
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1636968456
transform 1 0 81788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 1
transform 1 0 82892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1636968456
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1636968456
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1636968456
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1636968456
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1636968456
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1636968456
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1636968456
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1636968456
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1636968456
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1636968456
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1636968456
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1045
timestamp 1636968456
transform 1 0 97244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1057
timestamp 1
transform 1 0 98348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1636968456
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1636968456
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1636968456
transform 1 0 101292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1636968456
transform 1 0 102396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1
transform 1 0 103500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1636968456
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1636968456
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1636968456
transform 1 0 106444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1157
timestamp 1
transform 1 0 107548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1165
timestamp 1
transform 1 0 108284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636968456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636968456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636968456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636968456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636968456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636968456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636968456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636968456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636968456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636968456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636968456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636968456
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636968456
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636968456
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636968456
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636968456
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636968456
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636968456
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636968456
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636968456
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636968456
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636968456
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636968456
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636968456
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1636968456
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1636968456
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1636968456
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1636968456
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1636968456
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1636968456
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1636968456
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1636968456
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1636968456
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1636968456
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1636968456
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1636968456
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1636968456
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1636968456
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1636968456
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1636968456
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1636968456
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1636968456
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1636968456
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1636968456
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1636968456
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1636968456
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1636968456
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1636968456
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1636968456
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1636968456
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1636968456
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1636968456
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1636968456
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1636968456
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1636968456
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1636968456
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1636968456
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1636968456
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1636968456
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1636968456
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1636968456
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1636968456
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1636968456
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1161
timestamp 1
transform 1 0 107916 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1167
timestamp 1
transform 1 0 108468 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636968456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636968456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636968456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636968456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636968456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636968456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636968456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636968456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636968456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636968456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636968456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636968456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636968456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636968456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636968456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636968456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636968456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636968456
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636968456
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636968456
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636968456
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636968456
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636968456
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636968456
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636968456
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636968456
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636968456
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636968456
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636968456
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636968456
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636968456
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636968456
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636968456
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636968456
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1636968456
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1636968456
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1636968456
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636968456
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636968456
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1636968456
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1636968456
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1636968456
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1636968456
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1636968456
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1636968456
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1636968456
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1636968456
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1636968456
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1636968456
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1636968456
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1636968456
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1636968456
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1636968456
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1636968456
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1636968456
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1636968456
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1636968456
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1636968456
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1636968456
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1636968456
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1636968456
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1636968456
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1636968456
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1636968456
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1636968456
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1636968456
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1636968456
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1636968456
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1157
timestamp 1
transform 1 0 107548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1165
timestamp 1
transform 1 0 108284 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636968456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636968456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636968456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636968456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636968456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636968456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636968456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636968456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636968456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636968456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636968456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636968456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636968456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636968456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636968456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636968456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636968456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636968456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636968456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636968456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1636968456
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1636968456
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636968456
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636968456
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1636968456
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1636968456
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636968456
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636968456
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1636968456
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1636968456
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636968456
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636968456
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1636968456
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1636968456
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636968456
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636968456
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1636968456
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1636968456
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636968456
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636968456
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1636968456
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1636968456
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636968456
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636968456
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1636968456
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1636968456
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1636968456
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1636968456
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1636968456
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1636968456
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1636968456
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1636968456
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1636968456
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1636968456
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1636968456
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1636968456
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1636968456
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1636968456
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1636968456
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1636968456
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1636968456
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1636968456
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1636968456
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1636968456
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1636968456
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1636968456
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1636968456
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1636968456
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1636968456
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1636968456
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1636968456
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1161
timestamp 1
transform 1 0 107916 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1167
timestamp 1
transform 1 0 108468 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636968456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636968456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636968456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636968456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636968456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636968456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636968456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636968456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636968456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636968456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636968456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636968456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636968456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636968456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636968456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636968456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636968456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636968456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636968456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636968456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636968456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636968456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636968456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636968456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636968456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636968456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1636968456
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1636968456
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1636968456
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1636968456
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1636968456
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1636968456
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1636968456
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1636968456
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1636968456
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1636968456
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1636968456
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1636968456
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1636968456
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1636968456
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1636968456
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1636968456
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1636968456
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1636968456
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1636968456
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1636968456
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1636968456
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1636968456
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1636968456
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1636968456
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1636968456
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1636968456
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1636968456
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1636968456
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1636968456
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1636968456
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1636968456
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1636968456
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1636968456
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1636968456
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1636968456
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1636968456
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1636968456
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1636968456
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1636968456
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1636968456
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1636968456
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1636968456
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1636968456
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1636968456
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1636968456
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1636968456
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1636968456
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1636968456
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1636968456
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1636968456
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1636968456
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1157
timestamp 1
transform 1 0 107548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1165
timestamp 1
transform 1 0 108284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636968456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636968456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636968456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636968456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636968456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636968456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636968456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636968456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636968456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636968456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636968456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636968456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636968456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636968456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636968456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636968456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636968456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636968456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636968456
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636968456
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636968456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636968456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636968456
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1636968456
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636968456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636968456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1636968456
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1636968456
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1636968456
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1636968456
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1636968456
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1636968456
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1636968456
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1636968456
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1636968456
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1636968456
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1636968456
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1636968456
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1636968456
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1636968456
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1636968456
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1636968456
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1636968456
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1636968456
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1636968456
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1636968456
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1636968456
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1636968456
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1636968456
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1636968456
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1636968456
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1636968456
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1636968456
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1636968456
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1636968456
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1636968456
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1636968456
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1636968456
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1636968456
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1636968456
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1636968456
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1636968456
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1636968456
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1636968456
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1636968456
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1636968456
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1636968456
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1636968456
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1636968456
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1636968456
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1636968456
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1636968456
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1636968456
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1636968456
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1636968456
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1636968456
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1636968456
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1161
timestamp 1
transform 1 0 107916 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1167
timestamp 1
transform 1 0 108468 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636968456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636968456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636968456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636968456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636968456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636968456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636968456
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636968456
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636968456
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636968456
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636968456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636968456
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636968456
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636968456
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636968456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636968456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636968456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636968456
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636968456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636968456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636968456
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636968456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636968456
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636968456
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636968456
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636968456
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636968456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636968456
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1636968456
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1636968456
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1636968456
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1636968456
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1636968456
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1636968456
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1636968456
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1636968456
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1636968456
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1636968456
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1636968456
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1636968456
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1636968456
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1636968456
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1636968456
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1636968456
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1636968456
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1636968456
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1636968456
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1636968456
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1636968456
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1636968456
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1636968456
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1636968456
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1636968456
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1636968456
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1636968456
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1636968456
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1636968456
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1636968456
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1636968456
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1636968456
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1636968456
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1636968456
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1636968456
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1636968456
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1636968456
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1636968456
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1636968456
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1636968456
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1636968456
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1636968456
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1636968456
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1636968456
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1636968456
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1636968456
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1636968456
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1636968456
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1636968456
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1636968456
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1636968456
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1636968456
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1636968456
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1157
timestamp 1
transform 1 0 107548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1165
timestamp 1
transform 1 0 108284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636968456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636968456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636968456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636968456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636968456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636968456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636968456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636968456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636968456
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636968456
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636968456
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636968456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636968456
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636968456
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636968456
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636968456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636968456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636968456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636968456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636968456
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636968456
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636968456
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636968456
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636968456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636968456
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1636968456
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1636968456
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636968456
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636968456
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1636968456
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1636968456
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1636968456
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1636968456
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1636968456
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1636968456
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1636968456
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1636968456
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1636968456
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1636968456
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1636968456
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1636968456
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1636968456
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1636968456
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1636968456
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1636968456
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1636968456
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1636968456
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1636968456
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1636968456
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1636968456
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1636968456
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1636968456
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1636968456
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1636968456
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1636968456
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1636968456
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1636968456
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1636968456
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1636968456
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1636968456
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1636968456
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1636968456
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1636968456
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1636968456
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1636968456
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1636968456
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1636968456
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1636968456
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1636968456
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1636968456
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1636968456
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1636968456
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1636968456
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1636968456
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1636968456
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1636968456
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1636968456
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1636968456
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1636968456
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1636968456
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1161
timestamp 1
transform 1 0 107916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1167
timestamp 1
transform 1 0 108468 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_29
timestamp 1636968456
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_41
timestamp 1636968456
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636968456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636968456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp 1
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_85
timestamp 1636968456
transform 1 0 8924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_97
timestamp 1636968456
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636968456
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636968456
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp 1
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_141
timestamp 1636968456
transform 1 0 14076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_153
timestamp 1
transform 1 0 15180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636968456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636968456
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1636968456
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_209
timestamp 1636968456
transform 1 0 20332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636968456
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636968456
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_249
timestamp 1
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1636968456
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1636968456
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636968456
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636968456
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_305
timestamp 1
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_309
timestamp 1636968456
transform 1 0 29532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_321
timestamp 1636968456
transform 1 0 30636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636968456
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1636968456
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp 1
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_365
timestamp 1636968456
transform 1 0 34684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_377
timestamp 1636968456
transform 1 0 35788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636968456
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1636968456
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_417
timestamp 1
transform 1 0 39468 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_421
timestamp 1636968456
transform 1 0 39836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_433
timestamp 1636968456
transform 1 0 40940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1636968456
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1636968456
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_473
timestamp 1
transform 1 0 44620 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_477
timestamp 1636968456
transform 1 0 44988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_489
timestamp 1636968456
transform 1 0 46092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1636968456
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1636968456
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_529
timestamp 1
transform 1 0 49772 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_533
timestamp 1636968456
transform 1 0 50140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_545
timestamp 1636968456
transform 1 0 51244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_557
timestamp 1
transform 1 0 52348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1636968456
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1636968456
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_585
timestamp 1
transform 1 0 54924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_589
timestamp 1636968456
transform 1 0 55292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_601
timestamp 1636968456
transform 1 0 56396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_613
timestamp 1
transform 1 0 57500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1636968456
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1636968456
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_641
timestamp 1
transform 1 0 60076 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_645
timestamp 1636968456
transform 1 0 60444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_657
timestamp 1636968456
transform 1 0 61548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_669
timestamp 1
transform 1 0 62652 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1636968456
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1636968456
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_697
timestamp 1
transform 1 0 65228 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_701
timestamp 1636968456
transform 1 0 65596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_713
timestamp 1636968456
transform 1 0 66700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_725
timestamp 1
transform 1 0 67804 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1636968456
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1636968456
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_753
timestamp 1
transform 1 0 70380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_757
timestamp 1636968456
transform 1 0 70748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_769
timestamp 1636968456
transform 1 0 71852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_781
timestamp 1
transform 1 0 72956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1636968456
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1636968456
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_809
timestamp 1
transform 1 0 75532 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_813
timestamp 1636968456
transform 1 0 75900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_825
timestamp 1636968456
transform 1 0 77004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_837
timestamp 1
transform 1 0 78108 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1636968456
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1636968456
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_865
timestamp 1
transform 1 0 80684 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_869
timestamp 1636968456
transform 1 0 81052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_881
timestamp 1636968456
transform 1 0 82156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_893
timestamp 1
transform 1 0 83260 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1636968456
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1636968456
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_921
timestamp 1
transform 1 0 85836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_925
timestamp 1636968456
transform 1 0 86204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_937
timestamp 1636968456
transform 1 0 87308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_949
timestamp 1
transform 1 0 88412 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1636968456
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_965
timestamp 1
transform 1 0 89884 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_971
timestamp 1
transform 1 0 90436 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_978
timestamp 1
transform 1 0 91080 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_981
timestamp 1636968456
transform 1 0 91356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_993
timestamp 1636968456
transform 1 0 92460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1005
timestamp 1
transform 1 0 93564 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1636968456
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1636968456
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1033
timestamp 1
transform 1 0 96140 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1037
timestamp 1636968456
transform 1 0 96508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1049
timestamp 1636968456
transform 1 0 97612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1061
timestamp 1
transform 1 0 98716 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1636968456
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1636968456
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1089
timestamp 1
transform 1 0 101292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1093
timestamp 1636968456
transform 1 0 101660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1105
timestamp 1636968456
transform 1 0 102764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1117
timestamp 1
transform 1 0 103868 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1636968456
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1636968456
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1145
timestamp 1
transform 1 0 106444 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1149
timestamp 1636968456
transform 1 0 106812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1161
timestamp 1
transform 1 0 107916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1167
timestamp 1
transform 1 0 108468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636968456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636968456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636968456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636968456
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 1
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1122
timestamp 1636968456
transform 1 0 104328 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1134
timestamp 1636968456
transform 1 0 105432 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1146
timestamp 1
transform 1 0 106536 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1148
timestamp 1636968456
transform 1 0 106720 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1160
timestamp 1
transform 1 0 107824 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636968456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636968456
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636968456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1122
timestamp 1636968456
transform 1 0 104328 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1134
timestamp 1636968456
transform 1 0 105432 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1146
timestamp 1636968456
transform 1 0 106536 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1158
timestamp 1
transform 1 0 107640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1166
timestamp 1
transform 1 0 108376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636968456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636968456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636968456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636968456
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_65
timestamp 1
transform 1 0 7084 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1122
timestamp 1636968456
transform 1 0 104328 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1134
timestamp 1636968456
transform 1 0 105432 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1146
timestamp 1
transform 1 0 106536 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1148
timestamp 1636968456
transform 1 0 106720 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1160
timestamp 1
transform 1 0 107824 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636968456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636968456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636968456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636968456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_69
timestamp 1
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1122
timestamp 1636968456
transform 1 0 104328 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1134
timestamp 1636968456
transform 1 0 105432 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1146
timestamp 1636968456
transform 1 0 106536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1158
timestamp 1
transform 1 0 107640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1166
timestamp 1
transform 1 0 108376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636968456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636968456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636968456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636968456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1
transform 1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1122
timestamp 1636968456
transform 1 0 104328 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1134
timestamp 1636968456
transform 1 0 105432 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1146
timestamp 1
transform 1 0 106536 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1148
timestamp 1636968456
transform 1 0 106720 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1160
timestamp 1
transform 1 0 107824 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636968456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636968456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636968456
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636968456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1122
timestamp 1636968456
transform 1 0 104328 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1134
timestamp 1636968456
transform 1 0 105432 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1146
timestamp 1636968456
transform 1 0 106536 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1158
timestamp 1
transform 1 0 107640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1166
timestamp 1
transform 1 0 108376 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636968456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636968456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636968456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636968456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_65
timestamp 1
transform 1 0 7084 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1122
timestamp 1636968456
transform 1 0 104328 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1134
timestamp 1636968456
transform 1 0 105432 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1146
timestamp 1
transform 1 0 106536 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1148
timestamp 1636968456
transform 1 0 106720 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1160
timestamp 1
transform 1 0 107824 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636968456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636968456
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1636968456
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1636968456
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636968456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1122
timestamp 1636968456
transform 1 0 104328 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1134
timestamp 1636968456
transform 1 0 105432 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1146
timestamp 1636968456
transform 1 0 106536 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1158
timestamp 1
transform 1 0 107640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1166
timestamp 1
transform 1 0 108376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636968456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636968456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636968456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636968456
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636968456
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_65
timestamp 1
transform 1 0 7084 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1122
timestamp 1636968456
transform 1 0 104328 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1134
timestamp 1636968456
transform 1 0 105432 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1146
timestamp 1
transform 1 0 106536 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1148
timestamp 1636968456
transform 1 0 106720 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1160
timestamp 1
transform 1 0 107824 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636968456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636968456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636968456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1636968456
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636968456
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1122
timestamp 1636968456
transform 1 0 104328 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1134
timestamp 1636968456
transform 1 0 105432 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1146
timestamp 1636968456
transform 1 0 106536 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1158
timestamp 1
transform 1 0 107640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1166
timestamp 1
transform 1 0 108376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636968456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636968456
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636968456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636968456
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636968456
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_65
timestamp 1
transform 1 0 7084 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1122
timestamp 1636968456
transform 1 0 104328 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1134
timestamp 1636968456
transform 1 0 105432 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1146
timestamp 1
transform 1 0 106536 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1148
timestamp 1636968456
transform 1 0 106720 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1160
timestamp 1
transform 1 0 107824 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636968456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636968456
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636968456
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1636968456
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636968456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1122
timestamp 1636968456
transform 1 0 104328 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1134
timestamp 1636968456
transform 1 0 105432 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1146
timestamp 1636968456
transform 1 0 106536 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_1158
timestamp 1
transform 1 0 107640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_1166
timestamp 1
transform 1 0 108376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636968456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636968456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636968456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636968456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636968456
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_65
timestamp 1
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1122
timestamp 1636968456
transform 1 0 104328 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1134
timestamp 1636968456
transform 1 0 105432 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1146
timestamp 1
transform 1 0 106536 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1148
timestamp 1636968456
transform 1 0 106720 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_1160
timestamp 1
transform 1 0 107824 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636968456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636968456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636968456
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636968456
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1122
timestamp 1636968456
transform 1 0 104328 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1134
timestamp 1636968456
transform 1 0 105432 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1146
timestamp 1636968456
transform 1 0 106536 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_1158
timestamp 1
transform 1 0 107640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_1166
timestamp 1
transform 1 0 108376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636968456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636968456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636968456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636968456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636968456
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_65
timestamp 1
transform 1 0 7084 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1122
timestamp 1636968456
transform 1 0 104328 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1134
timestamp 1636968456
transform 1 0 105432 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1146
timestamp 1
transform 1 0 106536 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1148
timestamp 1636968456
transform 1 0 106720 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_1160
timestamp 1
transform 1 0 107824 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1636968456
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1636968456
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_32
timestamp 1636968456
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1636968456
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636968456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1122
timestamp 1636968456
transform 1 0 104328 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1134
timestamp 1636968456
transform 1 0 105432 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1146
timestamp 1636968456
transform 1 0 106536 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_1158
timestamp 1
transform 1 0 107640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_1166
timestamp 1
transform 1 0 108376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636968456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636968456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636968456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636968456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636968456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_65
timestamp 1
transform 1 0 7084 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1122
timestamp 1636968456
transform 1 0 104328 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1134
timestamp 1636968456
transform 1 0 105432 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1146
timestamp 1
transform 1 0 106536 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1148
timestamp 1636968456
transform 1 0 106720 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_1160
timestamp 1
transform 1 0 107824 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636968456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636968456
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636968456
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636968456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1122
timestamp 1636968456
transform 1 0 104328 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1134
timestamp 1636968456
transform 1 0 105432 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1146
timestamp 1636968456
transform 1 0 106536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_1158
timestamp 1
transform 1 0 107640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_1166
timestamp 1
transform 1 0 108376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636968456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636968456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636968456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636968456
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_65
timestamp 1
transform 1 0 7084 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1122
timestamp 1636968456
transform 1 0 104328 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1134
timestamp 1636968456
transform 1 0 105432 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1146
timestamp 1
transform 1 0 106536 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1148
timestamp 1636968456
transform 1 0 106720 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_1160
timestamp 1
transform 1 0 107824 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636968456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636968456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636968456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636968456
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636968456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1122
timestamp 1636968456
transform 1 0 104328 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1134
timestamp 1636968456
transform 1 0 105432 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1146
timestamp 1636968456
transform 1 0 106536 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_1158
timestamp 1
transform 1 0 107640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_1166
timestamp 1
transform 1 0 108376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636968456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636968456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636968456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636968456
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636968456
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_65
timestamp 1
transform 1 0 7084 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1122
timestamp 1636968456
transform 1 0 104328 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1134
timestamp 1636968456
transform 1 0 105432 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1146
timestamp 1
transform 1 0 106536 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1148
timestamp 1636968456
transform 1 0 106720 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_1160
timestamp 1
transform 1 0 107824 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636968456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636968456
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636968456
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1636968456
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636968456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_69
timestamp 1
transform 1 0 7452 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1122
timestamp 1636968456
transform 1 0 104328 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1134
timestamp 1636968456
transform 1 0 105432 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1146
timestamp 1636968456
transform 1 0 106536 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_1158
timestamp 1
transform 1 0 107640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_1166
timestamp 1
transform 1 0 108376 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636968456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636968456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636968456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636968456
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636968456
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_65
timestamp 1
transform 1 0 7084 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1122
timestamp 1636968456
transform 1 0 104328 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1134
timestamp 1636968456
transform 1 0 105432 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1146
timestamp 1
transform 1 0 106536 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1148
timestamp 1636968456
transform 1 0 106720 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_1160
timestamp 1
transform 1 0 107824 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636968456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636968456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636968456
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1636968456
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636968456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1122
timestamp 1636968456
transform 1 0 104328 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1134
timestamp 1636968456
transform 1 0 105432 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1146
timestamp 1636968456
transform 1 0 106536 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_1158
timestamp 1
transform 1 0 107640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_1166
timestamp 1
transform 1 0 108376 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636968456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636968456
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636968456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1636968456
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1636968456
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_65
timestamp 1
transform 1 0 7084 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1122
timestamp 1636968456
transform 1 0 104328 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1134
timestamp 1636968456
transform 1 0 105432 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1146
timestamp 1
transform 1 0 106536 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1148
timestamp 1636968456
transform 1 0 106720 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_1160
timestamp 1
transform 1 0 107824 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636968456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636968456
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1636968456
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1636968456
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636968456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_69
timestamp 1
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1122
timestamp 1636968456
transform 1 0 104328 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1134
timestamp 1636968456
transform 1 0 105432 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1146
timestamp 1636968456
transform 1 0 106536 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_1158
timestamp 1
transform 1 0 107640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_1166
timestamp 1
transform 1 0 108376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636968456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636968456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636968456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1636968456
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1636968456
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_65
timestamp 1
transform 1 0 7084 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1122
timestamp 1636968456
transform 1 0 104328 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1134
timestamp 1636968456
transform 1 0 105432 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1146
timestamp 1
transform 1 0 106536 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1148
timestamp 1636968456
transform 1 0 106720 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_1160
timestamp 1
transform 1 0 107824 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1636968456
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1636968456
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1636968456
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1636968456
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636968456
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_69
timestamp 1
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1124
timestamp 1636968456
transform 1 0 104512 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1136
timestamp 1636968456
transform 1 0 105616 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1148
timestamp 1636968456
transform 1 0 106720 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_1160
timestamp 1
transform 1 0 107824 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636968456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636968456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636968456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636968456
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636968456
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_65
timestamp 1
transform 1 0 7084 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1122
timestamp 1636968456
transform 1 0 104328 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1134
timestamp 1636968456
transform 1 0 105432 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1146
timestamp 1
transform 1 0 106536 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1148
timestamp 1636968456
transform 1 0 106720 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_1160
timestamp 1
transform 1 0 107824 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636968456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636968456
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636968456
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1636968456
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636968456
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_69
timestamp 1
transform 1 0 7452 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1124
timestamp 1636968456
transform 1 0 104512 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1136
timestamp 1636968456
transform 1 0 105616 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1148
timestamp 1636968456
transform 1 0 106720 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_1160
timestamp 1
transform 1 0 107824 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636968456
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636968456
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636968456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636968456
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1636968456
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_65
timestamp 1
transform 1 0 7084 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1122
timestamp 1636968456
transform 1 0 104328 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1134
timestamp 1636968456
transform 1 0 105432 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1146
timestamp 1
transform 1 0 106536 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1148
timestamp 1636968456
transform 1 0 106720 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_1160
timestamp 1
transform 1 0 107824 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636968456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636968456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1636968456
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1636968456
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636968456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1122
timestamp 1636968456
transform 1 0 104328 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1134
timestamp 1636968456
transform 1 0 105432 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1146
timestamp 1636968456
transform 1 0 106536 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_1158
timestamp 1
transform 1 0 107640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_1166
timestamp 1
transform 1 0 108376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636968456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636968456
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636968456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636968456
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636968456
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_65
timestamp 1
transform 1 0 7084 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1124
timestamp 1636968456
transform 1 0 104512 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_1136
timestamp 1
transform 1 0 105616 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_1144
timestamp 1
transform 1 0 106352 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1148
timestamp 1636968456
transform 1 0 106720 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_1160
timestamp 1
transform 1 0 107824 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636968456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636968456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636968456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636968456
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636968456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_69
timestamp 1
transform 1 0 7452 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1122
timestamp 1636968456
transform 1 0 104328 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1134
timestamp 1636968456
transform 1 0 105432 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1146
timestamp 1636968456
transform 1 0 106536 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_1158
timestamp 1
transform 1 0 107640 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_1166
timestamp 1
transform 1 0 108376 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636968456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636968456
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636968456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636968456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636968456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_65
timestamp 1
transform 1 0 7084 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1122
timestamp 1636968456
transform 1 0 104328 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1134
timestamp 1636968456
transform 1 0 105432 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1146
timestamp 1
transform 1 0 106536 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1148
timestamp 1636968456
transform 1 0 106720 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_1160
timestamp 1
transform 1 0 107824 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636968456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636968456
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636968456
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636968456
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636968456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_69
timestamp 1
transform 1 0 7452 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1122
timestamp 1636968456
transform 1 0 104328 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1134
timestamp 1636968456
transform 1 0 105432 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1146
timestamp 1636968456
transform 1 0 106536 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_1158
timestamp 1
transform 1 0 107640 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_1166
timestamp 1
transform 1 0 108376 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636968456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636968456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636968456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636968456
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1636968456
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_65
timestamp 1
transform 1 0 7084 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1122
timestamp 1636968456
transform 1 0 104328 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1134
timestamp 1636968456
transform 1 0 105432 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1146
timestamp 1
transform 1 0 106536 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1148
timestamp 1636968456
transform 1 0 106720 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1160
timestamp 1
transform 1 0 107824 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636968456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636968456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1636968456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1636968456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636968456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_69
timestamp 1
transform 1 0 7452 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1122
timestamp 1636968456
transform 1 0 104328 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1134
timestamp 1636968456
transform 1 0 105432 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1146
timestamp 1636968456
transform 1 0 106536 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_1158
timestamp 1
transform 1 0 107640 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_1166
timestamp 1
transform 1 0 108376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636968456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636968456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636968456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636968456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1636968456
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_65
timestamp 1
transform 1 0 7084 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1122
timestamp 1636968456
transform 1 0 104328 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1134
timestamp 1636968456
transform 1 0 105432 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1146
timestamp 1
transform 1 0 106536 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1148
timestamp 1636968456
transform 1 0 106720 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_1160
timestamp 1
transform 1 0 107824 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636968456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1636968456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1636968456
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1636968456
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1636968456
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_69
timestamp 1
transform 1 0 7452 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1122
timestamp 1636968456
transform 1 0 104328 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1134
timestamp 1636968456
transform 1 0 105432 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1146
timestamp 1636968456
transform 1 0 106536 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_1158
timestamp 1
transform 1 0 107640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_1166
timestamp 1
transform 1 0 108376 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1636968456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1636968456
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636968456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1636968456
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1636968456
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_65
timestamp 1
transform 1 0 7084 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1122
timestamp 1636968456
transform 1 0 104328 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1134
timestamp 1636968456
transform 1 0 105432 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1146
timestamp 1
transform 1 0 106536 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1148
timestamp 1636968456
transform 1 0 106720 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_1160
timestamp 1
transform 1 0 107824 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636968456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636968456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1636968456
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1636968456
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1636968456
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_69
timestamp 1
transform 1 0 7452 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1122
timestamp 1636968456
transform 1 0 104328 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1134
timestamp 1636968456
transform 1 0 105432 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1146
timestamp 1636968456
transform 1 0 106536 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_1158
timestamp 1
transform 1 0 107640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_1166
timestamp 1
transform 1 0 108376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636968456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636968456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636968456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1636968456
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1636968456
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_65
timestamp 1
transform 1 0 7084 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1122
timestamp 1636968456
transform 1 0 104328 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1134
timestamp 1636968456
transform 1 0 105432 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1146
timestamp 1
transform 1 0 106536 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1148
timestamp 1636968456
transform 1 0 106720 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_1160
timestamp 1
transform 1 0 107824 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636968456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636968456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636968456
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1636968456
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1636968456
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_69
timestamp 1
transform 1 0 7452 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1122
timestamp 1636968456
transform 1 0 104328 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1134
timestamp 1636968456
transform 1 0 105432 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1146
timestamp 1636968456
transform 1 0 106536 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_1158
timestamp 1
transform 1 0 107640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_1166
timestamp 1
transform 1 0 108376 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636968456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636968456
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1636968456
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1636968456
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1636968456
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_65
timestamp 1
transform 1 0 7084 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1122
timestamp 1636968456
transform 1 0 104328 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1134
timestamp 1636968456
transform 1 0 105432 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1146
timestamp 1
transform 1 0 106536 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1148
timestamp 1636968456
transform 1 0 106720 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_1160
timestamp 1
transform 1 0 107824 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1636968456
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1636968456
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1636968456
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1636968456
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1636968456
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_69
timestamp 1
transform 1 0 7452 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1122
timestamp 1636968456
transform 1 0 104328 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1134
timestamp 1636968456
transform 1 0 105432 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1146
timestamp 1636968456
transform 1 0 106536 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_1158
timestamp 1
transform 1 0 107640 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_1166
timestamp 1
transform 1 0 108376 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636968456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636968456
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636968456
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1636968456
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1636968456
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_65
timestamp 1
transform 1 0 7084 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1122
timestamp 1636968456
transform 1 0 104328 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1134
timestamp 1636968456
transform 1 0 105432 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1146
timestamp 1
transform 1 0 106536 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1148
timestamp 1636968456
transform 1 0 106720 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_1160
timestamp 1
transform 1 0 107824 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1636968456
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1636968456
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1636968456
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1636968456
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1636968456
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_69
timestamp 1
transform 1 0 7452 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1122
timestamp 1636968456
transform 1 0 104328 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1134
timestamp 1636968456
transform 1 0 105432 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1146
timestamp 1636968456
transform 1 0 106536 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_1158
timestamp 1
transform 1 0 107640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_1166
timestamp 1
transform 1 0 108376 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636968456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636968456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636968456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1636968456
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1636968456
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_65
timestamp 1
transform 1 0 7084 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1122
timestamp 1636968456
transform 1 0 104328 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1134
timestamp 1636968456
transform 1 0 105432 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1146
timestamp 1
transform 1 0 106536 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1148
timestamp 1636968456
transform 1 0 106720 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_1160
timestamp 1
transform 1 0 107824 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_8
timestamp 1636968456
transform 1 0 1840 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_20
timestamp 1636968456
transform 1 0 2944 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_32
timestamp 1636968456
transform 1 0 4048 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_44
timestamp 1636968456
transform 1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1636968456
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_69
timestamp 1
transform 1 0 7452 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1122
timestamp 1636968456
transform 1 0 104328 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1134
timestamp 1636968456
transform 1 0 105432 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1146
timestamp 1636968456
transform 1 0 106536 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1158
timestamp 1
transform 1 0 107640 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_1166
timestamp 1
transform 1 0 108376 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1636968456
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1636968456
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636968456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1636968456
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1636968456
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_65
timestamp 1
transform 1 0 7084 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1122
timestamp 1636968456
transform 1 0 104328 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1134
timestamp 1636968456
transform 1 0 105432 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1146
timestamp 1
transform 1 0 106536 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1148
timestamp 1636968456
transform 1 0 106720 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_1160
timestamp 1
transform 1 0 107824 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_8
timestamp 1636968456
transform 1 0 1840 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_20
timestamp 1636968456
transform 1 0 2944 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_32
timestamp 1636968456
transform 1 0 4048 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_44
timestamp 1636968456
transform 1 0 5152 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1636968456
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_69
timestamp 1
transform 1 0 7452 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1122
timestamp 1636968456
transform 1 0 104328 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1134
timestamp 1636968456
transform 1 0 105432 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1146
timestamp 1636968456
transform 1 0 106536 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1158
timestamp 1
transform 1 0 107640 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1166
timestamp 1
transform 1 0 108376 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636968456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636968456
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1636968456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1636968456
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1636968456
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_65
timestamp 1
transform 1 0 7084 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1122
timestamp 1636968456
transform 1 0 104328 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1134
timestamp 1636968456
transform 1 0 105432 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1146
timestamp 1
transform 1 0 106536 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1148
timestamp 1636968456
transform 1 0 106720 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1160
timestamp 1
transform 1 0 107824 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636968456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636968456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1636968456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1636968456
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1636968456
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_69
timestamp 1
transform 1 0 7452 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1122
timestamp 1636968456
transform 1 0 104328 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1134
timestamp 1636968456
transform 1 0 105432 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1146
timestamp 1636968456
transform 1 0 106536 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1158
timestamp 1
transform 1 0 107640 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1166
timestamp 1
transform 1 0 108376 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_8
timestamp 1636968456
transform 1 0 1840 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_20
timestamp 1
transform 1 0 2944 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1636968456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1636968456
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1636968456
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_65
timestamp 1
transform 1 0 7084 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1128
timestamp 1636968456
transform 1 0 104880 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_1140
timestamp 1
transform 1 0 105984 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1146
timestamp 1
transform 1 0 106536 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1148
timestamp 1636968456
transform 1 0 106720 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_1160
timestamp 1
transform 1 0 107824 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1636968456
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1636968456
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1636968456
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1636968456
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1636968456
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_69
timestamp 1
transform 1 0 7452 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1144
timestamp 1636968456
transform 1 0 106352 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1156
timestamp 1636968456
transform 1 0 107456 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_8
timestamp 1636968456
transform 1 0 1840 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_20
timestamp 1
transform 1 0 2944 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1636968456
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1636968456
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1636968456
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_65
timestamp 1
transform 1 0 7084 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1122
timestamp 1636968456
transform 1 0 104328 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1134
timestamp 1636968456
transform 1 0 105432 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_1146
timestamp 1
transform 1 0 106536 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1148
timestamp 1636968456
transform 1 0 106720 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_1160
timestamp 1
transform 1 0 107824 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1636968456
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1636968456
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1636968456
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1636968456
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1636968456
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_69
timestamp 1
transform 1 0 7452 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1122
timestamp 1636968456
transform 1 0 104328 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1134
timestamp 1636968456
transform 1 0 105432 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1146
timestamp 1636968456
transform 1 0 106536 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_1158
timestamp 1
transform 1 0 107640 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_1166
timestamp 1
transform 1 0 108376 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636968456
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636968456
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636968456
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1636968456
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1636968456
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_65
timestamp 1
transform 1 0 7084 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1122
timestamp 1636968456
transform 1 0 104328 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1134
timestamp 1636968456
transform 1 0 105432 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_1146
timestamp 1
transform 1 0 106536 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1148
timestamp 1636968456
transform 1 0 106720 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_1160
timestamp 1
transform 1 0 107824 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_8
timestamp 1636968456
transform 1 0 1840 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_20
timestamp 1636968456
transform 1 0 2944 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_32
timestamp 1636968456
transform 1 0 4048 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_44
timestamp 1636968456
transform 1 0 5152 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1636968456
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_69
timestamp 1
transform 1 0 7452 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1122
timestamp 1636968456
transform 1 0 104328 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1134
timestamp 1636968456
transform 1 0 105432 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1146
timestamp 1636968456
transform 1 0 106536 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_1158
timestamp 1
transform 1 0 107640 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_1166
timestamp 1
transform 1 0 108376 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1636968456
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1636968456
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636968456
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1636968456
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1636968456
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_65
timestamp 1
transform 1 0 7084 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1122
timestamp 1636968456
transform 1 0 104328 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1134
timestamp 1636968456
transform 1 0 105432 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_1146
timestamp 1
transform 1 0 106536 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1148
timestamp 1636968456
transform 1 0 106720 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_1160
timestamp 1
transform 1 0 107824 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636968456
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636968456
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1636968456
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1636968456
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1636968456
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_69
timestamp 1
transform 1 0 7452 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1122
timestamp 1636968456
transform 1 0 104328 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1134
timestamp 1636968456
transform 1 0 105432 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1146
timestamp 1636968456
transform 1 0 106536 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_1158
timestamp 1
transform 1 0 107640 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_1166
timestamp 1
transform 1 0 108376 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_8
timestamp 1636968456
transform 1 0 1840 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_20
timestamp 1
transform 1 0 2944 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636968456
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1636968456
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1636968456
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_65
timestamp 1
transform 1 0 7084 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1122
timestamp 1636968456
transform 1 0 104328 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1134
timestamp 1636968456
transform 1 0 105432 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_1146
timestamp 1
transform 1 0 106536 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1148
timestamp 1636968456
transform 1 0 106720 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_1160
timestamp 1
transform 1 0 107824 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636968456
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636968456
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636968456
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1636968456
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1636968456
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_69
timestamp 1
transform 1 0 7452 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_1122
timestamp 1
transform 1 0 104328 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1131
timestamp 1636968456
transform 1 0 105156 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1143
timestamp 1636968456
transform 1 0 106260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1155
timestamp 1636968456
transform 1 0 107364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_1167
timestamp 1
transform 1 0 108468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636968456
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636968456
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636968456
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1636968456
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1636968456
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_65
timestamp 1
transform 1 0 7084 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1122
timestamp 1636968456
transform 1 0 104328 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1134
timestamp 1636968456
transform 1 0 105432 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1146
timestamp 1
transform 1 0 106536 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1148
timestamp 1636968456
transform 1 0 106720 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_1160
timestamp 1
transform 1 0 107824 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636968456
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1636968456
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1636968456
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1636968456
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1636968456
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_69
timestamp 1
transform 1 0 7452 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1122
timestamp 1636968456
transform 1 0 104328 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1134
timestamp 1636968456
transform 1 0 105432 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1146
timestamp 1636968456
transform 1 0 106536 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_1158
timestamp 1
transform 1 0 107640 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_1166
timestamp 1
transform 1 0 108376 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636968456
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636968456
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1636968456
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1636968456
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1636968456
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_65
timestamp 1
transform 1 0 7084 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1122
timestamp 1636968456
transform 1 0 104328 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1134
timestamp 1636968456
transform 1 0 105432 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_1146
timestamp 1
transform 1 0 106536 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1148
timestamp 1636968456
transform 1 0 106720 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_1160
timestamp 1
transform 1 0 107824 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1636968456
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1636968456
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1636968456
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1636968456
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1636968456
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_69
timestamp 1
transform 1 0 7452 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1137
timestamp 1636968456
transform 1 0 105708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1149
timestamp 1636968456
transform 1 0 106812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_1161
timestamp 1
transform 1 0 107916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_1167
timestamp 1
transform 1 0 108468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636968456
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636968456
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1636968456
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1636968456
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1636968456
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_65
timestamp 1
transform 1 0 7084 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1133
timestamp 1636968456
transform 1 0 105340 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_1145
timestamp 1
transform 1 0 106444 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1148
timestamp 1636968456
transform 1 0 106720 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_1160
timestamp 1
transform 1 0 107824 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636968456
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636968456
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1636968456
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1636968456
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1636968456
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_69
timestamp 1
transform 1 0 7452 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1129
timestamp 1636968456
transform 1 0 104972 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1141
timestamp 1636968456
transform 1 0 106076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1153
timestamp 1636968456
transform 1 0 107180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_1165
timestamp 1
transform 1 0 108284 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636968456
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636968456
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1636968456
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1636968456
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1636968456
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_65
timestamp 1
transform 1 0 7084 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1125
timestamp 1636968456
transform 1 0 104604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_1137
timestamp 1
transform 1 0 105708 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_1145
timestamp 1
transform 1 0 106444 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1148
timestamp 1636968456
transform 1 0 106720 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_1160
timestamp 1
transform 1 0 107824 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1636968456
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1636968456
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1636968456
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1636968456
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1636968456
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_69
timestamp 1
transform 1 0 7452 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1122
timestamp 1636968456
transform 1 0 104328 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1134
timestamp 1636968456
transform 1 0 105432 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1146
timestamp 1636968456
transform 1 0 106536 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_1158
timestamp 1
transform 1 0 107640 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_1166
timestamp 1
transform 1 0 108376 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1636968456
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1636968456
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1636968456
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1636968456
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1636968456
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_65
timestamp 1
transform 1 0 7084 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1122
timestamp 1636968456
transform 1 0 104328 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1134
timestamp 1636968456
transform 1 0 105432 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_1146
timestamp 1
transform 1 0 106536 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1148
timestamp 1636968456
transform 1 0 106720 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_1160
timestamp 1
transform 1 0 107824 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636968456
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636968456
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1636968456
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1636968456
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1636968456
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_69
timestamp 1
transform 1 0 7452 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1122
timestamp 1636968456
transform 1 0 104328 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1134
timestamp 1636968456
transform 1 0 105432 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1146
timestamp 1636968456
transform 1 0 106536 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_1158
timestamp 1
transform 1 0 107640 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_1166
timestamp 1
transform 1 0 108376 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636968456
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1636968456
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1636968456
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1636968456
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1636968456
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_65
timestamp 1
transform 1 0 7084 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1122
timestamp 1636968456
transform 1 0 104328 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1134
timestamp 1636968456
transform 1 0 105432 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_1146
timestamp 1
transform 1 0 106536 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1148
timestamp 1636968456
transform 1 0 106720 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_1160
timestamp 1
transform 1 0 107824 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1636968456
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1636968456
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1636968456
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1636968456
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1636968456
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_69
timestamp 1
transform 1 0 7452 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1122
timestamp 1636968456
transform 1 0 104328 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1134
timestamp 1636968456
transform 1 0 105432 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1146
timestamp 1636968456
transform 1 0 106536 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_1158
timestamp 1
transform 1 0 107640 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_1166
timestamp 1
transform 1 0 108376 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1636968456
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1636968456
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1636968456
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1636968456
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1636968456
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_65
timestamp 1
transform 1 0 7084 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1124
timestamp 1636968456
transform 1 0 104512 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_1136
timestamp 1
transform 1 0 105616 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_1144
timestamp 1
transform 1 0 106352 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1148
timestamp 1636968456
transform 1 0 106720 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_1160
timestamp 1
transform 1 0 107824 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1636968456
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1636968456
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1636968456
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1636968456
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1636968456
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_69
timestamp 1
transform 1 0 7452 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1135
timestamp 1636968456
transform 1 0 105524 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1147
timestamp 1636968456
transform 1 0 106628 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_1159
timestamp 1
transform 1 0 107732 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_1167
timestamp 1
transform 1 0 108468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1636968456
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1636968456
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1636968456
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1636968456
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1636968456
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_65
timestamp 1
transform 1 0 7084 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1122
timestamp 1636968456
transform 1 0 104328 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1134
timestamp 1636968456
transform 1 0 105432 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_1146
timestamp 1
transform 1 0 106536 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1148
timestamp 1636968456
transform 1 0 106720 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_1160
timestamp 1
transform 1 0 107824 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1636968456
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1636968456
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1636968456
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1636968456
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1636968456
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_69
timestamp 1
transform 1 0 7452 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1126
timestamp 1636968456
transform 1 0 104696 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1138
timestamp 1636968456
transform 1 0 105800 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1150
timestamp 1636968456
transform 1 0 106904 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_1162
timestamp 1
transform 1 0 108008 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1636968456
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1636968456
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1636968456
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1636968456
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1636968456
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_65
timestamp 1
transform 1 0 7084 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1135
timestamp 1636968456
transform 1 0 105524 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1148
timestamp 1636968456
transform 1 0 106720 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_1160
timestamp 1
transform 1 0 107824 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1636968456
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1636968456
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1636968456
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1636968456
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1636968456
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_69
timestamp 1
transform 1 0 7452 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1124
timestamp 1636968456
transform 1 0 104512 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1136
timestamp 1636968456
transform 1 0 105616 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1148
timestamp 1636968456
transform 1 0 106720 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_1160
timestamp 1
transform 1 0 107824 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1636968456
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1636968456
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1636968456
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1636968456
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1636968456
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_65
timestamp 1
transform 1 0 7084 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1122
timestamp 1636968456
transform 1 0 104328 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1134
timestamp 1636968456
transform 1 0 105432 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_1146
timestamp 1
transform 1 0 106536 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1148
timestamp 1636968456
transform 1 0 106720 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_1160
timestamp 1
transform 1 0 107824 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1636968456
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1636968456
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1636968456
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1636968456
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1636968456
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_69
timestamp 1
transform 1 0 7452 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1122
timestamp 1636968456
transform 1 0 104328 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1134
timestamp 1636968456
transform 1 0 105432 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1146
timestamp 1636968456
transform 1 0 106536 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_1158
timestamp 1
transform 1 0 107640 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_1166
timestamp 1
transform 1 0 108376 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1636968456
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1636968456
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1636968456
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1636968456
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1636968456
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_65
timestamp 1
transform 1 0 7084 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1122
timestamp 1636968456
transform 1 0 104328 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1134
timestamp 1636968456
transform 1 0 105432 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_1146
timestamp 1
transform 1 0 106536 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1148
timestamp 1636968456
transform 1 0 106720 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_1160
timestamp 1
transform 1 0 107824 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1636968456
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1636968456
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1636968456
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1636968456
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1636968456
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_69
timestamp 1
transform 1 0 7452 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1126
timestamp 1636968456
transform 1 0 104696 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1138
timestamp 1636968456
transform 1 0 105800 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1150
timestamp 1636968456
transform 1 0 106904 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_1162
timestamp 1
transform 1 0 108008 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1636968456
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1636968456
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1636968456
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1636968456
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1636968456
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_65
timestamp 1
transform 1 0 7084 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1134
timestamp 1636968456
transform 1 0 105432 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_1146
timestamp 1
transform 1 0 106536 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1148
timestamp 1636968456
transform 1 0 106720 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_1160
timestamp 1
transform 1 0 107824 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1636968456
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1636968456
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1636968456
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1636968456
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1636968456
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_69
timestamp 1
transform 1 0 7452 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1130
timestamp 1636968456
transform 1 0 105064 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1142
timestamp 1636968456
transform 1 0 106168 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1154
timestamp 1636968456
transform 1 0 107272 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_1166
timestamp 1
transform 1 0 108376 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1636968456
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1636968456
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1636968456
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1636968456
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1636968456
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_65
timestamp 1
transform 1 0 7084 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1122
timestamp 1636968456
transform 1 0 104328 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1134
timestamp 1636968456
transform 1 0 105432 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_1146
timestamp 1
transform 1 0 106536 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1148
timestamp 1636968456
transform 1 0 106720 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_1160
timestamp 1
transform 1 0 107824 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1636968456
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1636968456
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1636968456
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1636968456
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1636968456
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_69
timestamp 1
transform 1 0 7452 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1130
timestamp 1636968456
transform 1 0 105064 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1142
timestamp 1636968456
transform 1 0 106168 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1154
timestamp 1636968456
transform 1 0 107272 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_1166
timestamp 1
transform 1 0 108376 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1636968456
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1636968456
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1636968456
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1636968456
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1636968456
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_65
timestamp 1
transform 1 0 7084 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1134
timestamp 1636968456
transform 1 0 105432 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_1146
timestamp 1
transform 1 0 106536 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1148
timestamp 1636968456
transform 1 0 106720 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_1160
timestamp 1
transform 1 0 107824 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1636968456
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1636968456
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_27
timestamp 1636968456
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_39
timestamp 1636968456
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1636968456
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_69
timestamp 1
transform 1 0 7452 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1126
timestamp 1636968456
transform 1 0 104696 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1138
timestamp 1636968456
transform 1 0 105800 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1150
timestamp 1636968456
transform 1 0 106904 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_1162
timestamp 1
transform 1 0 108008 0 -1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_102_3
timestamp 1636968456
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_15
timestamp 1636968456
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1636968456
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1636968456
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1636968456
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_65
timestamp 1
transform 1 0 7084 0 1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1124
timestamp 1636968456
transform 1 0 104512 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_1136
timestamp 1
transform 1 0 105616 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_102_1144
timestamp 1
transform 1 0 106352 0 1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1148
timestamp 1636968456
transform 1 0 106720 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_1160
timestamp 1
transform 1 0 107824 0 1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1636968456
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1636968456
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_27
timestamp 1636968456
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_39
timestamp 1636968456
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_51
timestamp 1
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1636968456
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_69
timestamp 1
transform 1 0 7452 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1144
timestamp 1636968456
transform 1 0 106352 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1156
timestamp 1636968456
transform 1 0 107456 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_3
timestamp 1636968456
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_15
timestamp 1636968456
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1636968456
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1636968456
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1636968456
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_65
timestamp 1
transform 1 0 7084 0 1 58752
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1122
timestamp 1636968456
transform 1 0 104328 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1134
timestamp 1636968456
transform 1 0 105432 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_1146
timestamp 1
transform 1 0 106536 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1148
timestamp 1636968456
transform 1 0 106720 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_1160
timestamp 1
transform 1 0 107824 0 1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_105_3
timestamp 1636968456
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_15
timestamp 1636968456
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_27
timestamp 1636968456
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_39
timestamp 1636968456
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_57
timestamp 1636968456
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_69
timestamp 1
transform 1 0 7452 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1125
timestamp 1636968456
transform 1 0 104604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1137
timestamp 1636968456
transform 1 0 105708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1149
timestamp 1636968456
transform 1 0 106812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_1161
timestamp 1
transform 1 0 107916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_1167
timestamp 1
transform 1 0 108468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1636968456
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1636968456
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1636968456
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1636968456
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_53
timestamp 1636968456
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_65
timestamp 1
transform 1 0 7084 0 1 59840
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1125
timestamp 1636968456
transform 1 0 104604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_1137
timestamp 1
transform 1 0 105708 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_1145
timestamp 1
transform 1 0 106444 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1148
timestamp 1636968456
transform 1 0 106720 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_1160
timestamp 1
transform 1 0 107824 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_107_3
timestamp 1636968456
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_15
timestamp 1636968456
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_27
timestamp 1636968456
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_39
timestamp 1636968456
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_51
timestamp 1
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1636968456
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_69
timestamp 1
transform 1 0 7452 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1122
timestamp 1636968456
transform 1 0 104328 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1134
timestamp 1636968456
transform 1 0 105432 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1146
timestamp 1636968456
transform 1 0 106536 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_1158
timestamp 1
transform 1 0 107640 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_1166
timestamp 1
transform 1 0 108376 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1636968456
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1636968456
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1636968456
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_41
timestamp 1636968456
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_53
timestamp 1636968456
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_65
timestamp 1
transform 1 0 7084 0 1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1122
timestamp 1636968456
transform 1 0 104328 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1134
timestamp 1636968456
transform 1 0 105432 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_1146
timestamp 1
transform 1 0 106536 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1148
timestamp 1636968456
transform 1 0 106720 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_1160
timestamp 1
transform 1 0 107824 0 1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_109_11
timestamp 1636968456
transform 1 0 2116 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_23
timestamp 1636968456
transform 1 0 3220 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_35
timestamp 1636968456
transform 1 0 4324 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_47
timestamp 1
transform 1 0 5428 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_57
timestamp 1636968456
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_69
timestamp 1
transform 1 0 7452 0 -1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1122
timestamp 1636968456
transform 1 0 104328 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1134
timestamp 1636968456
transform 1 0 105432 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1146
timestamp 1636968456
transform 1 0 106536 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_1158
timestamp 1
transform 1 0 107640 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_1166
timestamp 1
transform 1 0 108376 0 -1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_110_11
timestamp 1636968456
transform 1 0 2116 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_23
timestamp 1
transform 1 0 3220 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_29
timestamp 1636968456
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_41
timestamp 1636968456
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_53
timestamp 1636968456
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_65
timestamp 1
transform 1 0 7084 0 1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1122
timestamp 1636968456
transform 1 0 104328 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1134
timestamp 1636968456
transform 1 0 105432 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_1146
timestamp 1
transform 1 0 106536 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1148
timestamp 1636968456
transform 1 0 106720 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_1160
timestamp 1
transform 1 0 107824 0 1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_111_8
timestamp 1636968456
transform 1 0 1840 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_20
timestamp 1636968456
transform 1 0 2944 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_32
timestamp 1636968456
transform 1 0 4048 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_44
timestamp 1636968456
transform 1 0 5152 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_57
timestamp 1636968456
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_69
timestamp 1
transform 1 0 7452 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1122
timestamp 1636968456
transform 1 0 104328 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1134
timestamp 1636968456
transform 1 0 105432 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1146
timestamp 1636968456
transform 1 0 106536 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_1158
timestamp 1
transform 1 0 107640 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_111_1166
timestamp 1
transform 1 0 108376 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_112_8
timestamp 1636968456
transform 1 0 1840 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_20
timestamp 1
transform 1 0 2944 0 1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1636968456
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_41
timestamp 1636968456
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_53
timestamp 1636968456
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_65
timestamp 1
transform 1 0 7084 0 1 63104
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1122
timestamp 1636968456
transform 1 0 104328 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1134
timestamp 1636968456
transform 1 0 105432 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_1146
timestamp 1
transform 1 0 106536 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1148
timestamp 1636968456
transform 1 0 106720 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_1160
timestamp 1
transform 1 0 107824 0 1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1636968456
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1636968456
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_27
timestamp 1636968456
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_39
timestamp 1636968456
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_57
timestamp 1636968456
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_113_69
timestamp 1
transform 1 0 7452 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1122
timestamp 1636968456
transform 1 0 104328 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1134
timestamp 1636968456
transform 1 0 105432 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1146
timestamp 1636968456
transform 1 0 106536 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_1158
timestamp 1
transform 1 0 107640 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_113_1166
timestamp 1
transform 1 0 108376 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_114_8
timestamp 1636968456
transform 1 0 1840 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_20
timestamp 1
transform 1 0 2944 0 1 64192
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1636968456
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_41
timestamp 1636968456
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_53
timestamp 1636968456
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_65
timestamp 1
transform 1 0 7084 0 1 64192
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1122
timestamp 1636968456
transform 1 0 104328 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1134
timestamp 1636968456
transform 1 0 105432 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_1146
timestamp 1
transform 1 0 106536 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1148
timestamp 1636968456
transform 1 0 106720 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_114_1160
timestamp 1
transform 1 0 107824 0 1 64192
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_115_8
timestamp 1636968456
transform 1 0 1840 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_20
timestamp 1636968456
transform 1 0 2944 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_32
timestamp 1636968456
transform 1 0 4048 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_44
timestamp 1636968456
transform 1 0 5152 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_57
timestamp 1636968456
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_115_69
timestamp 1
transform 1 0 7452 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1122
timestamp 1636968456
transform 1 0 104328 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1134
timestamp 1636968456
transform 1 0 105432 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1146
timestamp 1636968456
transform 1 0 106536 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_1158
timestamp 1
transform 1 0 107640 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_1162
timestamp 1
transform 1 0 108008 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_8
timestamp 1636968456
transform 1 0 1840 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_20
timestamp 1
transform 1 0 2944 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_116_29
timestamp 1636968456
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_41
timestamp 1636968456
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_53
timestamp 1636968456
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_65
timestamp 1
transform 1 0 7084 0 1 65280
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1122
timestamp 1636968456
transform 1 0 104328 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1134
timestamp 1636968456
transform 1 0 105432 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_1146
timestamp 1
transform 1 0 106536 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1148
timestamp 1636968456
transform 1 0 106720 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_116_1160
timestamp 1
transform 1 0 107824 0 1 65280
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_8
timestamp 1636968456
transform 1 0 1840 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_20
timestamp 1
transform 1 0 2944 0 -1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_117_29
timestamp 1636968456
transform 1 0 3772 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_41
timestamp 1636968456
transform 1 0 4876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_53
timestamp 1
transform 1 0 5980 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_57
timestamp 1636968456
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_69
timestamp 1636968456
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_81
timestamp 1
transform 1 0 8556 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_85
timestamp 1636968456
transform 1 0 8924 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_97
timestamp 1636968456
transform 1 0 10028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_109
timestamp 1
transform 1 0 11132 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_113
timestamp 1636968456
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_125
timestamp 1636968456
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_137
timestamp 1
transform 1 0 13708 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_141
timestamp 1636968456
transform 1 0 14076 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_153
timestamp 1636968456
transform 1 0 15180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_165
timestamp 1
transform 1 0 16284 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_169
timestamp 1636968456
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_181
timestamp 1
transform 1 0 17756 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_117_219
timestamp 1
transform 1 0 21252 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_117_249
timestamp 1
transform 1 0 24012 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_253
timestamp 1636968456
transform 1 0 24380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_265
timestamp 1636968456
transform 1 0 25484 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_277
timestamp 1
transform 1 0 26588 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_281
timestamp 1636968456
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_293
timestamp 1
transform 1 0 28060 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_117_301
timestamp 1
transform 1 0 28796 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_304
timestamp 1
transform 1 0 29072 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_117_309
timestamp 1636968456
transform 1 0 29532 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_321
timestamp 1
transform 1 0 30636 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_117_329
timestamp 1
transform 1 0 31372 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_335
timestamp 1
transform 1 0 31924 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_337
timestamp 1636968456
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_349
timestamp 1636968456
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_361
timestamp 1
transform 1 0 34316 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_365
timestamp 1636968456
transform 1 0 34684 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_377
timestamp 1636968456
transform 1 0 35788 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_389
timestamp 1
transform 1 0 36892 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_393
timestamp 1636968456
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_405
timestamp 1636968456
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_417
timestamp 1
transform 1 0 39468 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_421
timestamp 1636968456
transform 1 0 39836 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_433
timestamp 1636968456
transform 1 0 40940 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_445
timestamp 1
transform 1 0 42044 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_449
timestamp 1636968456
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_461
timestamp 1636968456
transform 1 0 43516 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_473
timestamp 1
transform 1 0 44620 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_477
timestamp 1636968456
transform 1 0 44988 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_489
timestamp 1636968456
transform 1 0 46092 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_501
timestamp 1
transform 1 0 47196 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_505
timestamp 1636968456
transform 1 0 47564 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_517
timestamp 1636968456
transform 1 0 48668 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_529
timestamp 1
transform 1 0 49772 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_533
timestamp 1636968456
transform 1 0 50140 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_545
timestamp 1636968456
transform 1 0 51244 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_557
timestamp 1
transform 1 0 52348 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_117_561
timestamp 1
transform 1 0 52716 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_117_569
timestamp 1
transform 1 0 53452 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_572
timestamp 1636968456
transform 1 0 53728 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_584
timestamp 1
transform 1 0 54832 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_117_589
timestamp 1
transform 1 0 55292 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_595
timestamp 1
transform 1 0 55844 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_621
timestamp 1636968456
transform 1 0 58236 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_633
timestamp 1
transform 1 0 59340 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_117_641
timestamp 1
transform 1 0 60076 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_645
timestamp 1636968456
transform 1 0 60444 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_657
timestamp 1636968456
transform 1 0 61548 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_669
timestamp 1
transform 1 0 62652 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_673
timestamp 1636968456
transform 1 0 63020 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_685
timestamp 1636968456
transform 1 0 64124 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_697
timestamp 1
transform 1 0 65228 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_701
timestamp 1636968456
transform 1 0 65596 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_713
timestamp 1636968456
transform 1 0 66700 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_725
timestamp 1
transform 1 0 67804 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_729
timestamp 1636968456
transform 1 0 68172 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_741
timestamp 1636968456
transform 1 0 69276 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_753
timestamp 1
transform 1 0 70380 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_757
timestamp 1636968456
transform 1 0 70748 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_769
timestamp 1636968456
transform 1 0 71852 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_781
timestamp 1
transform 1 0 72956 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_785
timestamp 1636968456
transform 1 0 73324 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_797
timestamp 1636968456
transform 1 0 74428 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_809
timestamp 1
transform 1 0 75532 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_813
timestamp 1636968456
transform 1 0 75900 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_825
timestamp 1636968456
transform 1 0 77004 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_837
timestamp 1
transform 1 0 78108 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_841
timestamp 1636968456
transform 1 0 78476 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_853
timestamp 1636968456
transform 1 0 79580 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_865
timestamp 1
transform 1 0 80684 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_869
timestamp 1636968456
transform 1 0 81052 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_881
timestamp 1636968456
transform 1 0 82156 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_893
timestamp 1
transform 1 0 83260 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_919
timestamp 1
transform 1 0 85652 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_923
timestamp 1
transform 1 0 86020 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_117_953
timestamp 1
transform 1 0 88780 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1000
timestamp 1
transform 1 0 93104 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1005
timestamp 1
transform 1 0 93564 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1063
timestamp 1
transform 1 0 98900 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_1084
timestamp 1
transform 1 0 100832 0 -1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1093
timestamp 1636968456
transform 1 0 101660 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1105
timestamp 1636968456
transform 1 0 102764 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1117
timestamp 1
transform 1 0 103868 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1121
timestamp 1636968456
transform 1 0 104236 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1133
timestamp 1636968456
transform 1 0 105340 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1145
timestamp 1
transform 1 0 106444 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1149
timestamp 1636968456
transform 1 0 106812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_1161
timestamp 1
transform 1 0 107916 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1636968456
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1636968456
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1636968456
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_41
timestamp 1636968456
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_53
timestamp 1636968456
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_65
timestamp 1636968456
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_85
timestamp 1636968456
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_97
timestamp 1636968456
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_109
timestamp 1636968456
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_121
timestamp 1636968456
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_141
timestamp 1636968456
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_153
timestamp 1636968456
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_165
timestamp 1
transform 1 0 16284 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_118_173
timestamp 1
transform 1 0 17020 0 1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_118_180
timestamp 1636968456
transform 1 0 17664 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_192
timestamp 1
transform 1 0 18768 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_118_197
timestamp 1
transform 1 0 19228 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_205
timestamp 1
transform 1 0 19964 0 1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_118_234
timestamp 1636968456
transform 1 0 22632 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_246
timestamp 1
transform 1 0 23736 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_118_275
timestamp 1
transform 1 0 26404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_281
timestamp 1
transform 1 0 26956 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_118_305
timestamp 1
transform 1 0 29164 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_118_313
timestamp 1
transform 1 0 29900 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_118_339
timestamp 1
transform 1 0 32292 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_118_361
timestamp 1
transform 1 0 34316 0 1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_118_365
timestamp 1636968456
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_377
timestamp 1636968456
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_389
timestamp 1636968456
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_401
timestamp 1636968456
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_413
timestamp 1
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_419
timestamp 1
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_421
timestamp 1636968456
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_433
timestamp 1636968456
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_445
timestamp 1636968456
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_457
timestamp 1636968456
transform 1 0 43148 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_469
timestamp 1
transform 1 0 44252 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_475
timestamp 1
transform 1 0 44804 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_477
timestamp 1636968456
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_489
timestamp 1636968456
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_501
timestamp 1636968456
transform 1 0 47196 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_513
timestamp 1636968456
transform 1 0 48300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_525
timestamp 1
transform 1 0 49404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_531
timestamp 1
transform 1 0 49956 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_533
timestamp 1636968456
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_545
timestamp 1636968456
transform 1 0 51244 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_557
timestamp 1636968456
transform 1 0 52348 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_569
timestamp 1636968456
transform 1 0 53452 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_581
timestamp 1
transform 1 0 54556 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_587
timestamp 1
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_589
timestamp 1
transform 1 0 55292 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_597
timestamp 1
transform 1 0 56028 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_609
timestamp 1636968456
transform 1 0 57132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_621
timestamp 1636968456
transform 1 0 58236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_633
timestamp 1
transform 1 0 59340 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_641
timestamp 1
transform 1 0 60076 0 1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_118_645
timestamp 1636968456
transform 1 0 60444 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_657
timestamp 1636968456
transform 1 0 61548 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_669
timestamp 1636968456
transform 1 0 62652 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_681
timestamp 1636968456
transform 1 0 63756 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_693
timestamp 1
transform 1 0 64860 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_699
timestamp 1
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_701
timestamp 1636968456
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_713
timestamp 1636968456
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_118_725
timestamp 1
transform 1 0 67804 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_118_729
timestamp 1
transform 1 0 68172 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_733
timestamp 1
transform 1 0 68540 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_118_755
timestamp 1
transform 1 0 70564 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_118_759
timestamp 1
transform 1 0 70932 0 1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_118_765
timestamp 1636968456
transform 1 0 71484 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_777
timestamp 1636968456
transform 1 0 72588 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_789
timestamp 1636968456
transform 1 0 73692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_801
timestamp 1
transform 1 0 74796 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_809
timestamp 1
transform 1 0 75532 0 1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_118_813
timestamp 1636968456
transform 1 0 75900 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_825
timestamp 1
transform 1 0 77004 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_118_860
timestamp 1
transform 1 0 80224 0 1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_118_869
timestamp 1636968456
transform 1 0 81052 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_881
timestamp 1
transform 1 0 82156 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_118_922
timestamp 1
transform 1 0 85928 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_118_977
timestamp 1
transform 1 0 90988 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1037
timestamp 1
transform 1 0 96508 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1043
timestamp 1636968456
transform 1 0 97060 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1073
timestamp 1636968456
transform 1 0 99820 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1085
timestamp 1
transform 1 0 100924 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1091
timestamp 1
transform 1 0 101476 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1102
timestamp 1636968456
transform 1 0 102488 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1114
timestamp 1636968456
transform 1 0 103592 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1126
timestamp 1636968456
transform 1 0 104696 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_1138
timestamp 1
transform 1 0 105800 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_118_1146
timestamp 1
transform 1 0 106536 0 1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1149
timestamp 1636968456
transform 1 0 106812 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1161
timestamp 1
transform 1 0 107916 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1167
timestamp 1
transform 1 0 108468 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_8
timestamp 1636968456
transform 1 0 1840 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_20
timestamp 1636968456
transform 1 0 2944 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_32
timestamp 1636968456
transform 1 0 4048 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_44
timestamp 1636968456
transform 1 0 5152 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_57
timestamp 1636968456
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_69
timestamp 1636968456
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_81
timestamp 1636968456
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_93
timestamp 1636968456
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_113
timestamp 1636968456
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_125
timestamp 1636968456
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_137
timestamp 1636968456
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_149
timestamp 1636968456
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_169
timestamp 1636968456
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_181
timestamp 1636968456
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_119_217
timestamp 1
transform 1 0 21068 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_119_221
timestamp 1
transform 1 0 21436 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_119_225
timestamp 1636968456
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_119_237
timestamp 1
transform 1 0 22908 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_119_263
timestamp 1636968456
transform 1 0 25300 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_275
timestamp 1
transform 1 0 26404 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_279
timestamp 1
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_281
timestamp 1636968456
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_293
timestamp 1636968456
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_305
timestamp 1
transform 1 0 29164 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_313
timestamp 1
transform 1 0 29900 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_119_326
timestamp 1
transform 1 0 31096 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_119_334
timestamp 1
transform 1 0 31832 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_119_337
timestamp 1
transform 1 0 32108 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_119_345
timestamp 1
transform 1 0 32844 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_119_362
timestamp 1
transform 1 0 34408 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_119_381
timestamp 1
transform 1 0 36156 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_389
timestamp 1
transform 1 0 36892 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_119_393
timestamp 1636968456
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_405
timestamp 1
transform 1 0 38364 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_119_421
timestamp 1
transform 1 0 39836 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_119_437
timestamp 1
transform 1 0 41308 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_445
timestamp 1
transform 1 0 42044 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_119_449
timestamp 1636968456
transform 1 0 42412 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_461
timestamp 1
transform 1 0 43516 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_465
timestamp 1
transform 1 0 43884 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_119_479
timestamp 1
transform 1 0 45172 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_487
timestamp 1
transform 1 0 45908 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_119_503
timestamp 1
transform 1 0 47380 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_507
timestamp 1636968456
transform 1 0 47748 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_519
timestamp 1636968456
transform 1 0 48852 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_531
timestamp 1636968456
transform 1 0 49956 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_543
timestamp 1636968456
transform 1 0 51060 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_555
timestamp 1
transform 1 0 52164 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_559
timestamp 1
transform 1 0 52532 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_561
timestamp 1636968456
transform 1 0 52716 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_573
timestamp 1636968456
transform 1 0 53820 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_585
timestamp 1636968456
transform 1 0 54924 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_597
timestamp 1636968456
transform 1 0 56028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_609
timestamp 1
transform 1 0 57132 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_615
timestamp 1
transform 1 0 57684 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_617
timestamp 1636968456
transform 1 0 57868 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_629
timestamp 1636968456
transform 1 0 58972 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_119_641
timestamp 1
transform 1 0 60076 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_119_667
timestamp 1
transform 1 0 62468 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_671
timestamp 1
transform 1 0 62836 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_673
timestamp 1636968456
transform 1 0 63020 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_685
timestamp 1636968456
transform 1 0 64124 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_697
timestamp 1636968456
transform 1 0 65228 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_119_724
timestamp 1
transform 1 0 67712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_119_727
timestamp 1
transform 1 0 67988 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_738
timestamp 1
transform 1 0 69000 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_742
timestamp 1
transform 1 0 69368 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_119_776
timestamp 1
transform 1 0 72496 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_119_796
timestamp 1
transform 1 0 74336 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_119_813
timestamp 1
transform 1 0 75900 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_119_821
timestamp 1
transform 1 0 76636 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_119_829
timestamp 1
transform 1 0 77372 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_837
timestamp 1
transform 1 0 78108 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_119_841
timestamp 1
transform 1 0 78476 0 -1 67456
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_119_851
timestamp 1636968456
transform 1 0 79396 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_863
timestamp 1636968456
transform 1 0 80500 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_875
timestamp 1636968456
transform 1 0 81604 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_887
timestamp 1
transform 1 0 82708 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_119_895
timestamp 1
transform 1 0 83444 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_897
timestamp 1636968456
transform 1 0 83628 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_909
timestamp 1
transform 1 0 84732 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_940
timestamp 1
transform 1 0 87584 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_119_944
timestamp 1
transform 1 0 87952 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_119_955
timestamp 1
transform 1 0 88964 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_984
timestamp 1
transform 1 0 91632 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1038
timestamp 1
transform 1 0 96600 0 -1 67456
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1074
timestamp 1636968456
transform 1 0 99912 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1086
timestamp 1
transform 1 0 101016 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1092
timestamp 1
transform 1 0 101568 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1097
timestamp 1636968456
transform 1 0 102028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_1109
timestamp 1
transform 1 0 103132 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_1117
timestamp 1
transform 1 0 103868 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1121
timestamp 1636968456
transform 1 0 104236 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1133
timestamp 1636968456
transform 1 0 105340 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1145
timestamp 1636968456
transform 1 0 106444 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1157
timestamp 1
transform 1 0 107548 0 -1 67456
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_120_11
timestamp 1636968456
transform 1 0 2116 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_120_23
timestamp 1
transform 1 0 3220 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1636968456
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_41
timestamp 1636968456
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_53
timestamp 1
transform 1 0 5980 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_57
timestamp 1636968456
transform 1 0 6348 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_69
timestamp 1636968456
transform 1 0 7452 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_81
timestamp 1
transform 1 0 8556 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_85
timestamp 1636968456
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_97
timestamp 1636968456
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_109
timestamp 1
transform 1 0 11132 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_113
timestamp 1636968456
transform 1 0 11500 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_125
timestamp 1636968456
transform 1 0 12604 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_137
timestamp 1
transform 1 0 13708 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_141
timestamp 1636968456
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_153
timestamp 1
transform 1 0 15180 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_120_161
timestamp 1
transform 1 0 15916 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_120_165
timestamp 1
transform 1 0 16284 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_169
timestamp 1636968456
transform 1 0 16652 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_181
timestamp 1636968456
transform 1 0 17756 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_193
timestamp 1
transform 1 0 18860 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_197
timestamp 1636968456
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_209
timestamp 1636968456
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_221
timestamp 1
transform 1 0 21436 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_225
timestamp 1636968456
transform 1 0 21804 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_237
timestamp 1
transform 1 0 22908 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_120_245
timestamp 1
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_251
timestamp 1
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_120_253
timestamp 1
transform 1 0 24380 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_120_258
timestamp 1
transform 1 0 24840 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_266
timestamp 1
transform 1 0 25576 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_120_271
timestamp 1
transform 1 0 26036 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_120_279
timestamp 1
transform 1 0 26772 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_283
timestamp 1
transform 1 0 27140 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_291
timestamp 1
transform 1 0 27876 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_120_296
timestamp 1
transform 1 0 28336 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_300
timestamp 1
transform 1 0 28704 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_120_306
timestamp 1
transform 1 0 29256 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_120_311
timestamp 1
transform 1 0 29716 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_120_321
timestamp 1
transform 1 0 30636 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_329
timestamp 1
transform 1 0 31372 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_120_334
timestamp 1
transform 1 0 31832 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_120_337
timestamp 1
transform 1 0 32108 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_120_347
timestamp 1
transform 1 0 33028 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_120_355
timestamp 1
transform 1 0 33764 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_120_359
timestamp 1
transform 1 0 34132 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_363
timestamp 1
transform 1 0 34500 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_120_365
timestamp 1
transform 1 0 34684 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_369
timestamp 1
transform 1 0 35052 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_372
timestamp 1
transform 1 0 35328 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_380
timestamp 1
transform 1 0 36064 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_120_385
timestamp 1
transform 1 0 36524 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_391
timestamp 1
transform 1 0 37076 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_120_393
timestamp 1
transform 1 0 37260 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_120_397
timestamp 1
transform 1 0 37628 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_405
timestamp 1
transform 1 0 38364 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_120_410
timestamp 1
transform 1 0 38824 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_120_418
timestamp 1
transform 1 0 39560 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_120_423
timestamp 1
transform 1 0 40020 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_431
timestamp 1
transform 1 0 40756 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_120_436
timestamp 1
transform 1 0 41216 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_120_444
timestamp 1
transform 1 0 41952 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_120_449
timestamp 1
transform 1 0 42412 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_120_457
timestamp 1
transform 1 0 43148 0 1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_120_461
timestamp 1636968456
transform 1 0 43516 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_473
timestamp 1
transform 1 0 44620 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_477
timestamp 1636968456
transform 1 0 44988 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_489
timestamp 1636968456
transform 1 0 46092 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_501
timestamp 1
transform 1 0 47196 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_505
timestamp 1636968456
transform 1 0 47564 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_517
timestamp 1636968456
transform 1 0 48668 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_529
timestamp 1
transform 1 0 49772 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_533
timestamp 1636968456
transform 1 0 50140 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_545
timestamp 1636968456
transform 1 0 51244 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_557
timestamp 1
transform 1 0 52348 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_561
timestamp 1636968456
transform 1 0 52716 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_573
timestamp 1636968456
transform 1 0 53820 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_585
timestamp 1
transform 1 0 54924 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_589
timestamp 1636968456
transform 1 0 55292 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_601
timestamp 1636968456
transform 1 0 56396 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_613
timestamp 1
transform 1 0 57500 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_617
timestamp 1636968456
transform 1 0 57868 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_629
timestamp 1636968456
transform 1 0 58972 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_641
timestamp 1
transform 1 0 60076 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_645
timestamp 1636968456
transform 1 0 60444 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_657
timestamp 1636968456
transform 1 0 61548 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_669
timestamp 1
transform 1 0 62652 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_673
timestamp 1636968456
transform 1 0 63020 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_685
timestamp 1636968456
transform 1 0 64124 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_697
timestamp 1
transform 1 0 65228 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_701
timestamp 1636968456
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_713
timestamp 1636968456
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_725
timestamp 1
transform 1 0 67804 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_729
timestamp 1636968456
transform 1 0 68172 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_120_741
timestamp 1
transform 1 0 69276 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_120_749
timestamp 1
transform 1 0 70012 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_755
timestamp 1
transform 1 0 70564 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_757
timestamp 1636968456
transform 1 0 70748 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_769
timestamp 1636968456
transform 1 0 71852 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_781
timestamp 1
transform 1 0 72956 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_785
timestamp 1636968456
transform 1 0 73324 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_797
timestamp 1636968456
transform 1 0 74428 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_809
timestamp 1
transform 1 0 75532 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_813
timestamp 1636968456
transform 1 0 75900 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_825
timestamp 1636968456
transform 1 0 77004 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_837
timestamp 1
transform 1 0 78108 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_841
timestamp 1636968456
transform 1 0 78476 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_853
timestamp 1636968456
transform 1 0 79580 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_865
timestamp 1
transform 1 0 80684 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_869
timestamp 1636968456
transform 1 0 81052 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_881
timestamp 1636968456
transform 1 0 82156 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_893
timestamp 1
transform 1 0 83260 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_897
timestamp 1636968456
transform 1 0 83628 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_909
timestamp 1636968456
transform 1 0 84732 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_921
timestamp 1
transform 1 0 85836 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_925
timestamp 1636968456
transform 1 0 86204 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_120_942
timestamp 1
transform 1 0 87768 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_946
timestamp 1
transform 1 0 88136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_120_950
timestamp 1
transform 1 0 88504 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_120_959
timestamp 1
transform 1 0 89332 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_120_979
timestamp 1
transform 1 0 91172 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1009
timestamp 1
transform 1 0 93932 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1045
timestamp 1636968456
transform 1 0 97244 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_1057
timestamp 1
transform 1 0 98348 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1063
timestamp 1
transform 1 0 98900 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1065
timestamp 1636968456
transform 1 0 99084 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1077
timestamp 1636968456
transform 1 0 100188 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_1089
timestamp 1
transform 1 0 101292 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1093
timestamp 1636968456
transform 1 0 101660 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1105
timestamp 1636968456
transform 1 0 102764 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_1117
timestamp 1
transform 1 0 103868 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1121
timestamp 1636968456
transform 1 0 104236 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1133
timestamp 1636968456
transform 1 0 105340 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_1145
timestamp 1
transform 1 0 106444 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1149
timestamp 1636968456
transform 1 0 106812 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_120_1161
timestamp 1
transform 1 0 107916 0 1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_121_11
timestamp 1636968456
transform 1 0 2116 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_23
timestamp 1636968456
transform 1 0 3220 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_35
timestamp 1636968456
transform 1 0 4324 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_47
timestamp 1
transform 1 0 5428 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_57
timestamp 1636968456
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_121_69
timestamp 1
transform 1 0 7452 0 -1 68544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1122
timestamp 1636968456
transform 1 0 104328 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1134
timestamp 1
transform 1 0 105432 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1140
timestamp 1636968456
transform 1 0 105984 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1152
timestamp 1636968456
transform 1 0 107088 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1164
timestamp 1
transform 1 0 108192 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_11
timestamp 1636968456
transform 1 0 2116 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_23
timestamp 1
transform 1 0 3220 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1636968456
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_41
timestamp 1636968456
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_53
timestamp 1636968456
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_65
timestamp 1
transform 1 0 7084 0 1 68544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1122
timestamp 1636968456
transform 1 0 104328 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1134
timestamp 1636968456
transform 1 0 105432 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1146
timestamp 1
transform 1 0 106536 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1148
timestamp 1636968456
transform 1 0 106720 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_122_1160
timestamp 1
transform 1 0 107824 0 1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1636968456
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1636968456
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_27
timestamp 1636968456
transform 1 0 3588 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_39
timestamp 1636968456
transform 1 0 4692 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_51
timestamp 1
transform 1 0 5796 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_57
timestamp 1636968456
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_69
timestamp 1
transform 1 0 7452 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1122
timestamp 1636968456
transform 1 0 104328 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1134
timestamp 1636968456
transform 1 0 105432 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1146
timestamp 1636968456
transform 1 0 106536 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_1158
timestamp 1
transform 1 0 107640 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_123_1166
timestamp 1
transform 1 0 108376 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_124_11
timestamp 1636968456
transform 1 0 2116 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_23
timestamp 1
transform 1 0 3220 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 1
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_29
timestamp 1636968456
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_41
timestamp 1636968456
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_53
timestamp 1636968456
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_65
timestamp 1
transform 1 0 7084 0 1 69632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1122
timestamp 1636968456
transform 1 0 104328 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1134
timestamp 1636968456
transform 1 0 105432 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1146
timestamp 1
transform 1 0 106536 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1148
timestamp 1636968456
transform 1 0 106720 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_124_1160
timestamp 1
transform 1 0 107824 0 1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_125_15
timestamp 1636968456
transform 1 0 2484 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_27
timestamp 1636968456
transform 1 0 3588 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_39
timestamp 1636968456
transform 1 0 4692 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_51
timestamp 1
transform 1 0 5796 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_57
timestamp 1636968456
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_125_69
timestamp 1
transform 1 0 7452 0 -1 70720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1122
timestamp 1636968456
transform 1 0 104328 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1134
timestamp 1636968456
transform 1 0 105432 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1146
timestamp 1636968456
transform 1 0 106536 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_1158
timestamp 1
transform 1 0 107640 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_125_1166
timestamp 1
transform 1 0 108376 0 -1 70720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_126_13
timestamp 1636968456
transform 1 0 2300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_126_25
timestamp 1
transform 1 0 3404 0 1 70720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_126_29
timestamp 1636968456
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_41
timestamp 1636968456
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_53
timestamp 1636968456
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_65
timestamp 1
transform 1 0 7084 0 1 70720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1122
timestamp 1636968456
transform 1 0 104328 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1134
timestamp 1636968456
transform 1 0 105432 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1146
timestamp 1
transform 1 0 106536 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1148
timestamp 1636968456
transform 1 0 106720 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_1160
timestamp 1
transform 1 0 107824 0 1 70720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_127_11
timestamp 1636968456
transform 1 0 2116 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_23
timestamp 1636968456
transform 1 0 3220 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_35
timestamp 1636968456
transform 1 0 4324 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_47
timestamp 1
transform 1 0 5428 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_57
timestamp 1636968456
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_127_69
timestamp 1
transform 1 0 7452 0 -1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1122
timestamp 1636968456
transform 1 0 104328 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1134
timestamp 1636968456
transform 1 0 105432 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1146
timestamp 1636968456
transform 1 0 106536 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_1158
timestamp 1
transform 1 0 107640 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_127_1166
timestamp 1
transform 1 0 108376 0 -1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_128_3
timestamp 1636968456
transform 1 0 1380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_15
timestamp 1636968456
transform 1 0 2484 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 1
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_29
timestamp 1636968456
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_41
timestamp 1636968456
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_53
timestamp 1636968456
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_65
timestamp 1
transform 1 0 7084 0 1 71808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1122
timestamp 1636968456
transform 1 0 104328 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1134
timestamp 1636968456
transform 1 0 105432 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1146
timestamp 1
transform 1 0 106536 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1148
timestamp 1636968456
transform 1 0 106720 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_1160
timestamp 1
transform 1 0 107824 0 1 71808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_129_11
timestamp 1636968456
transform 1 0 2116 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_23
timestamp 1636968456
transform 1 0 3220 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_35
timestamp 1636968456
transform 1 0 4324 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_47
timestamp 1
transform 1 0 5428 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_129_55
timestamp 1
transform 1 0 6164 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_57
timestamp 1636968456
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_129_69
timestamp 1
transform 1 0 7452 0 -1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1122
timestamp 1636968456
transform 1 0 104328 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1134
timestamp 1636968456
transform 1 0 105432 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1146
timestamp 1636968456
transform 1 0 106536 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_1158
timestamp 1
transform 1 0 107640 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_129_1166
timestamp 1
transform 1 0 108376 0 -1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_130_11
timestamp 1636968456
transform 1 0 2116 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_130_23
timestamp 1
transform 1 0 3220 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 1
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_29
timestamp 1636968456
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_41
timestamp 1636968456
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_53
timestamp 1636968456
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_65
timestamp 1
transform 1 0 7084 0 1 72896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1122
timestamp 1636968456
transform 1 0 104328 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1134
timestamp 1636968456
transform 1 0 105432 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1146
timestamp 1
transform 1 0 106536 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1148
timestamp 1636968456
transform 1 0 106720 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_1160
timestamp 1
transform 1 0 107824 0 1 72896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_131_11
timestamp 1636968456
transform 1 0 2116 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_23
timestamp 1636968456
transform 1 0 3220 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_35
timestamp 1636968456
transform 1 0 4324 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_47
timestamp 1
transform 1 0 5428 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_131_55
timestamp 1
transform 1 0 6164 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_57
timestamp 1636968456
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_131_69
timestamp 1
transform 1 0 7452 0 -1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1122
timestamp 1636968456
transform 1 0 104328 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1134
timestamp 1636968456
transform 1 0 105432 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1146
timestamp 1636968456
transform 1 0 106536 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_1158
timestamp 1
transform 1 0 107640 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_131_1166
timestamp 1
transform 1 0 108376 0 -1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_132_11
timestamp 1636968456
transform 1 0 2116 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_132_23
timestamp 1
transform 1 0 3220 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 1
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_29
timestamp 1636968456
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_41
timestamp 1636968456
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_53
timestamp 1636968456
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_65
timestamp 1
transform 1 0 7084 0 1 73984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1122
timestamp 1636968456
transform 1 0 104328 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1134
timestamp 1636968456
transform 1 0 105432 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1146
timestamp 1
transform 1 0 106536 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1148
timestamp 1636968456
transform 1 0 106720 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_1160
timestamp 1
transform 1 0 107824 0 1 73984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_133_3
timestamp 1636968456
transform 1 0 1380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_15
timestamp 1636968456
transform 1 0 2484 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_27
timestamp 1636968456
transform 1 0 3588 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_39
timestamp 1636968456
transform 1 0 4692 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_51
timestamp 1
transform 1 0 5796 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_133_55
timestamp 1
transform 1 0 6164 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_57
timestamp 1636968456
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_133_69
timestamp 1
transform 1 0 7452 0 -1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1122
timestamp 1636968456
transform 1 0 104328 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1134
timestamp 1636968456
transform 1 0 105432 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1146
timestamp 1636968456
transform 1 0 106536 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_1158
timestamp 1
transform 1 0 107640 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_133_1166
timestamp 1
transform 1 0 108376 0 -1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_134_11
timestamp 1636968456
transform 1 0 2116 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_134_23
timestamp 1
transform 1 0 3220 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 1
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_29
timestamp 1636968456
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_41
timestamp 1636968456
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_53
timestamp 1636968456
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_65
timestamp 1
transform 1 0 7084 0 1 75072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1127
timestamp 1636968456
transform 1 0 104788 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_1139
timestamp 1
transform 1 0 105892 0 1 75072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1148
timestamp 1636968456
transform 1 0 106720 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_1160
timestamp 1
transform 1 0 107824 0 1 75072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_135_8
timestamp 1636968456
transform 1 0 1840 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_20
timestamp 1636968456
transform 1 0 2944 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_32
timestamp 1636968456
transform 1 0 4048 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_44
timestamp 1636968456
transform 1 0 5152 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_57
timestamp 1636968456
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_135_69
timestamp 1
transform 1 0 7452 0 -1 76160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1144
timestamp 1636968456
transform 1 0 106352 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1156
timestamp 1636968456
transform 1 0 107456 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_11
timestamp 1636968456
transform 1 0 2116 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_23
timestamp 1
transform 1 0 3220 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 1
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_29
timestamp 1636968456
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_41
timestamp 1636968456
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_53
timestamp 1636968456
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_65
timestamp 1
transform 1 0 7084 0 1 76160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1122
timestamp 1636968456
transform 1 0 104328 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1134
timestamp 1636968456
transform 1 0 105432 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1146
timestamp 1
transform 1 0 106536 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1148
timestamp 1636968456
transform 1 0 106720 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_1160
timestamp 1
transform 1 0 107824 0 1 76160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_137_11
timestamp 1636968456
transform 1 0 2116 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_23
timestamp 1636968456
transform 1 0 3220 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_35
timestamp 1636968456
transform 1 0 4324 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_47
timestamp 1
transform 1 0 5428 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_57
timestamp 1636968456
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_137_69
timestamp 1
transform 1 0 7452 0 -1 77248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1122
timestamp 1636968456
transform 1 0 104328 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1134
timestamp 1636968456
transform 1 0 105432 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1146
timestamp 1636968456
transform 1 0 106536 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_1158
timestamp 1
transform 1 0 107640 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_137_1166
timestamp 1
transform 1 0 108376 0 -1 77248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_138_3
timestamp 1636968456
transform 1 0 1380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_15
timestamp 1636968456
transform 1 0 2484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 1
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_29
timestamp 1636968456
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_41
timestamp 1636968456
transform 1 0 4876 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_53
timestamp 1636968456
transform 1 0 5980 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_65
timestamp 1
transform 1 0 7084 0 1 77248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1132
timestamp 1636968456
transform 1 0 105248 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_1144
timestamp 1
transform 1 0 106352 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1148
timestamp 1636968456
transform 1 0 106720 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_1160
timestamp 1
transform 1 0 107824 0 1 77248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_139_11
timestamp 1636968456
transform 1 0 2116 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_23
timestamp 1636968456
transform 1 0 3220 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_35
timestamp 1636968456
transform 1 0 4324 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_47
timestamp 1
transform 1 0 5428 0 -1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_139_55
timestamp 1
transform 1 0 6164 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_57
timestamp 1636968456
transform 1 0 6348 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_139_69
timestamp 1
transform 1 0 7452 0 -1 78336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1144
timestamp 1636968456
transform 1 0 106352 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1156
timestamp 1636968456
transform 1 0 107456 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_11
timestamp 1636968456
transform 1 0 2116 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_140_23
timestamp 1
transform 1 0 3220 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_140_27
timestamp 1
transform 1 0 3588 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_29
timestamp 1636968456
transform 1 0 3772 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_41
timestamp 1636968456
transform 1 0 4876 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_53
timestamp 1636968456
transform 1 0 5980 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_65
timestamp 1
transform 1 0 7084 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_140_1137
timestamp 1
transform 1 0 105708 0 1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_140_1145
timestamp 1
transform 1 0 106444 0 1 78336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1148
timestamp 1636968456
transform 1 0 106720 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_1160
timestamp 1
transform 1 0 107824 0 1 78336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_141_3
timestamp 1636968456
transform 1 0 1380 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_15
timestamp 1636968456
transform 1 0 2484 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_27
timestamp 1636968456
transform 1 0 3588 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_39
timestamp 1636968456
transform 1 0 4692 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_141_51
timestamp 1
transform 1 0 5796 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_141_55
timestamp 1
transform 1 0 6164 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_57
timestamp 1636968456
transform 1 0 6348 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_141_69
timestamp 1
transform 1 0 7452 0 -1 79424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1130
timestamp 1636968456
transform 1 0 105064 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1142
timestamp 1636968456
transform 1 0 106168 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1154
timestamp 1636968456
transform 1 0 107272 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_141_1166
timestamp 1
transform 1 0 108376 0 -1 79424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_142_3
timestamp 1636968456
transform 1 0 1380 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_15
timestamp 1636968456
transform 1 0 2484 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_27
timestamp 1
transform 1 0 3588 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_29
timestamp 1636968456
transform 1 0 3772 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_41
timestamp 1636968456
transform 1 0 4876 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_53
timestamp 1636968456
transform 1 0 5980 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_65
timestamp 1
transform 1 0 7084 0 1 79424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1122
timestamp 1636968456
transform 1 0 104328 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1134
timestamp 1636968456
transform 1 0 105432 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_1146
timestamp 1
transform 1 0 106536 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1148
timestamp 1636968456
transform 1 0 106720 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_142_1160
timestamp 1
transform 1 0 107824 0 1 79424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_143_3
timestamp 1636968456
transform 1 0 1380 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_15
timestamp 1636968456
transform 1 0 2484 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_27
timestamp 1636968456
transform 1 0 3588 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_39
timestamp 1636968456
transform 1 0 4692 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_143_51
timestamp 1
transform 1 0 5796 0 -1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_143_55
timestamp 1
transform 1 0 6164 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_57
timestamp 1636968456
transform 1 0 6348 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_143_69
timestamp 1
transform 1 0 7452 0 -1 80512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1127
timestamp 1636968456
transform 1 0 104788 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1139
timestamp 1636968456
transform 1 0 105892 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1151
timestamp 1636968456
transform 1 0 106996 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_143_1163
timestamp 1
transform 1 0 108100 0 -1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_143_1167
timestamp 1
transform 1 0 108468 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_3
timestamp 1636968456
transform 1 0 1380 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_15
timestamp 1636968456
transform 1 0 2484 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_27
timestamp 1
transform 1 0 3588 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_29
timestamp 1636968456
transform 1 0 3772 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_41
timestamp 1636968456
transform 1 0 4876 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_53
timestamp 1636968456
transform 1 0 5980 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_65
timestamp 1
transform 1 0 7084 0 1 80512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1122
timestamp 1636968456
transform 1 0 104328 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1134
timestamp 1636968456
transform 1 0 105432 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_1146
timestamp 1
transform 1 0 106536 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1148
timestamp 1636968456
transform 1 0 106720 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_144_1160
timestamp 1
transform 1 0 107824 0 1 80512
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_145_3
timestamp 1636968456
transform 1 0 1380 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_15
timestamp 1636968456
transform 1 0 2484 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_27
timestamp 1636968456
transform 1 0 3588 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_39
timestamp 1636968456
transform 1 0 4692 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_145_51
timestamp 1
transform 1 0 5796 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_145_55
timestamp 1
transform 1 0 6164 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_57
timestamp 1636968456
transform 1 0 6348 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_145_69
timestamp 1
transform 1 0 7452 0 -1 81600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1122
timestamp 1636968456
transform 1 0 104328 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1134
timestamp 1636968456
transform 1 0 105432 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1146
timestamp 1636968456
transform 1 0 106536 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_145_1158
timestamp 1
transform 1 0 107640 0 -1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_145_1166
timestamp 1
transform 1 0 108376 0 -1 81600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_146_3
timestamp 1636968456
transform 1 0 1380 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_15
timestamp 1636968456
transform 1 0 2484 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_27
timestamp 1
transform 1 0 3588 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_29
timestamp 1636968456
transform 1 0 3772 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_41
timestamp 1636968456
transform 1 0 4876 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_53
timestamp 1636968456
transform 1 0 5980 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_65
timestamp 1
transform 1 0 7084 0 1 81600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1122
timestamp 1636968456
transform 1 0 104328 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1134
timestamp 1636968456
transform 1 0 105432 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_1146
timestamp 1
transform 1 0 106536 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1148
timestamp 1636968456
transform 1 0 106720 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_1160
timestamp 1
transform 1 0 107824 0 1 81600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_147_3
timestamp 1636968456
transform 1 0 1380 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_15
timestamp 1636968456
transform 1 0 2484 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_27
timestamp 1636968456
transform 1 0 3588 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_39
timestamp 1636968456
transform 1 0 4692 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_147_51
timestamp 1
transform 1 0 5796 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_147_55
timestamp 1
transform 1 0 6164 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_57
timestamp 1636968456
transform 1 0 6348 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_147_69
timestamp 1
transform 1 0 7452 0 -1 82688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1122
timestamp 1636968456
transform 1 0 104328 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1134
timestamp 1636968456
transform 1 0 105432 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1146
timestamp 1636968456
transform 1 0 106536 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_1158
timestamp 1
transform 1 0 107640 0 -1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_147_1166
timestamp 1
transform 1 0 108376 0 -1 82688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_148_3
timestamp 1636968456
transform 1 0 1380 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_15
timestamp 1636968456
transform 1 0 2484 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_27
timestamp 1
transform 1 0 3588 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_29
timestamp 1636968456
transform 1 0 3772 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_41
timestamp 1636968456
transform 1 0 4876 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_53
timestamp 1636968456
transform 1 0 5980 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_65
timestamp 1
transform 1 0 7084 0 1 82688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1122
timestamp 1636968456
transform 1 0 104328 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1134
timestamp 1636968456
transform 1 0 105432 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_1146
timestamp 1
transform 1 0 106536 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1148
timestamp 1636968456
transform 1 0 106720 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_148_1160
timestamp 1
transform 1 0 107824 0 1 82688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_149_3
timestamp 1636968456
transform 1 0 1380 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_15
timestamp 1636968456
transform 1 0 2484 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_27
timestamp 1636968456
transform 1 0 3588 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_39
timestamp 1636968456
transform 1 0 4692 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_149_51
timestamp 1
transform 1 0 5796 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_149_55
timestamp 1
transform 1 0 6164 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_57
timestamp 1636968456
transform 1 0 6348 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_149_69
timestamp 1
transform 1 0 7452 0 -1 83776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1122
timestamp 1636968456
transform 1 0 104328 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1134
timestamp 1636968456
transform 1 0 105432 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1146
timestamp 1636968456
transform 1 0 106536 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_1158
timestamp 1
transform 1 0 107640 0 -1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_149_1166
timestamp 1
transform 1 0 108376 0 -1 83776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_150_3
timestamp 1636968456
transform 1 0 1380 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_15
timestamp 1636968456
transform 1 0 2484 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_27
timestamp 1
transform 1 0 3588 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_29
timestamp 1636968456
transform 1 0 3772 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_41
timestamp 1636968456
transform 1 0 4876 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_53
timestamp 1636968456
transform 1 0 5980 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_65
timestamp 1
transform 1 0 7084 0 1 83776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1122
timestamp 1636968456
transform 1 0 104328 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1134
timestamp 1636968456
transform 1 0 105432 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_1146
timestamp 1
transform 1 0 106536 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1148
timestamp 1636968456
transform 1 0 106720 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_1160
timestamp 1
transform 1 0 107824 0 1 83776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_151_3
timestamp 1636968456
transform 1 0 1380 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_15
timestamp 1636968456
transform 1 0 2484 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_27
timestamp 1636968456
transform 1 0 3588 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_39
timestamp 1636968456
transform 1 0 4692 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_151_51
timestamp 1
transform 1 0 5796 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_151_55
timestamp 1
transform 1 0 6164 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_57
timestamp 1636968456
transform 1 0 6348 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_151_69
timestamp 1
transform 1 0 7452 0 -1 84864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1122
timestamp 1636968456
transform 1 0 104328 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1134
timestamp 1636968456
transform 1 0 105432 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1146
timestamp 1636968456
transform 1 0 106536 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_1158
timestamp 1
transform 1 0 107640 0 -1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_1166
timestamp 1
transform 1 0 108376 0 -1 84864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_152_3
timestamp 1636968456
transform 1 0 1380 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_15
timestamp 1636968456
transform 1 0 2484 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_152_27
timestamp 1
transform 1 0 3588 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_29
timestamp 1636968456
transform 1 0 3772 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_41
timestamp 1636968456
transform 1 0 4876 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_53
timestamp 1636968456
transform 1 0 5980 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_65
timestamp 1
transform 1 0 7084 0 1 84864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1128
timestamp 1636968456
transform 1 0 104880 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_1140
timestamp 1
transform 1 0 105984 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_1146
timestamp 1
transform 1 0 106536 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1148
timestamp 1636968456
transform 1 0 106720 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_1160
timestamp 1
transform 1 0 107824 0 1 84864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_153_3
timestamp 1636968456
transform 1 0 1380 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_15
timestamp 1636968456
transform 1 0 2484 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_27
timestamp 1636968456
transform 1 0 3588 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_39
timestamp 1636968456
transform 1 0 4692 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_153_51
timestamp 1
transform 1 0 5796 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_153_55
timestamp 1
transform 1 0 6164 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_57
timestamp 1636968456
transform 1 0 6348 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_153_69
timestamp 1
transform 1 0 7452 0 -1 85952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1129
timestamp 1636968456
transform 1 0 104972 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1141
timestamp 1636968456
transform 1 0 106076 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1153
timestamp 1636968456
transform 1 0 107180 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_153_1165
timestamp 1
transform 1 0 108284 0 -1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_154_3
timestamp 1636968456
transform 1 0 1380 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_15
timestamp 1636968456
transform 1 0 2484 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_27
timestamp 1
transform 1 0 3588 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_29
timestamp 1636968456
transform 1 0 3772 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_41
timestamp 1636968456
transform 1 0 4876 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_53
timestamp 1636968456
transform 1 0 5980 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_65
timestamp 1
transform 1 0 7084 0 1 85952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1128
timestamp 1636968456
transform 1 0 104880 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_1140
timestamp 1
transform 1 0 105984 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_1146
timestamp 1
transform 1 0 106536 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1148
timestamp 1636968456
transform 1 0 106720 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_1160
timestamp 1
transform 1 0 107824 0 1 85952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_155_3
timestamp 1636968456
transform 1 0 1380 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_15
timestamp 1636968456
transform 1 0 2484 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_27
timestamp 1636968456
transform 1 0 3588 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_39
timestamp 1636968456
transform 1 0 4692 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_155_51
timestamp 1
transform 1 0 5796 0 -1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_155_55
timestamp 1
transform 1 0 6164 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_57
timestamp 1636968456
transform 1 0 6348 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_155_69
timestamp 1
transform 1 0 7452 0 -1 87040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1122
timestamp 1636968456
transform 1 0 104328 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1134
timestamp 1636968456
transform 1 0 105432 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1146
timestamp 1636968456
transform 1 0 106536 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_155_1158
timestamp 1
transform 1 0 107640 0 -1 87040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_155_1166
timestamp 1
transform 1 0 108376 0 -1 87040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_156_3
timestamp 1636968456
transform 1 0 1380 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_15
timestamp 1636968456
transform 1 0 2484 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_156_27
timestamp 1
transform 1 0 3588 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_29
timestamp 1636968456
transform 1 0 3772 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_41
timestamp 1636968456
transform 1 0 4876 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_53
timestamp 1636968456
transform 1 0 5980 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_65
timestamp 1
transform 1 0 7084 0 1 87040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1122
timestamp 1636968456
transform 1 0 104328 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1134
timestamp 1636968456
transform 1 0 105432 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_156_1146
timestamp 1
transform 1 0 106536 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1148
timestamp 1636968456
transform 1 0 106720 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_156_1160
timestamp 1
transform 1 0 107824 0 1 87040
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_157_3
timestamp 1636968456
transform 1 0 1380 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_15
timestamp 1636968456
transform 1 0 2484 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_27
timestamp 1636968456
transform 1 0 3588 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_39
timestamp 1636968456
transform 1 0 4692 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_157_51
timestamp 1
transform 1 0 5796 0 -1 88128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_157_55
timestamp 1
transform 1 0 6164 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_57
timestamp 1636968456
transform 1 0 6348 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_157_69
timestamp 1
transform 1 0 7452 0 -1 88128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1122
timestamp 1636968456
transform 1 0 104328 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1134
timestamp 1636968456
transform 1 0 105432 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1146
timestamp 1636968456
transform 1 0 106536 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_1158
timestamp 1
transform 1 0 107640 0 -1 88128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_157_1166
timestamp 1
transform 1 0 108376 0 -1 88128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_158_3
timestamp 1636968456
transform 1 0 1380 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_15
timestamp 1636968456
transform 1 0 2484 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_27
timestamp 1
transform 1 0 3588 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_29
timestamp 1636968456
transform 1 0 3772 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_41
timestamp 1636968456
transform 1 0 4876 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_53
timestamp 1636968456
transform 1 0 5980 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_65
timestamp 1
transform 1 0 7084 0 1 88128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1122
timestamp 1636968456
transform 1 0 104328 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1134
timestamp 1636968456
transform 1 0 105432 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_1146
timestamp 1
transform 1 0 106536 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1148
timestamp 1636968456
transform 1 0 106720 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_158_1160
timestamp 1
transform 1 0 107824 0 1 88128
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_159_3
timestamp 1636968456
transform 1 0 1380 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_15
timestamp 1636968456
transform 1 0 2484 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_27
timestamp 1636968456
transform 1 0 3588 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_39
timestamp 1636968456
transform 1 0 4692 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_159_51
timestamp 1
transform 1 0 5796 0 -1 89216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_159_55
timestamp 1
transform 1 0 6164 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_57
timestamp 1636968456
transform 1 0 6348 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_159_69
timestamp 1
transform 1 0 7452 0 -1 89216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1122
timestamp 1636968456
transform 1 0 104328 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1134
timestamp 1636968456
transform 1 0 105432 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1146
timestamp 1636968456
transform 1 0 106536 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_1158
timestamp 1
transform 1 0 107640 0 -1 89216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_159_1166
timestamp 1
transform 1 0 108376 0 -1 89216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_160_3
timestamp 1636968456
transform 1 0 1380 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_15
timestamp 1636968456
transform 1 0 2484 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_27
timestamp 1
transform 1 0 3588 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_29
timestamp 1636968456
transform 1 0 3772 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_41
timestamp 1636968456
transform 1 0 4876 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_53
timestamp 1636968456
transform 1 0 5980 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_65
timestamp 1
transform 1 0 7084 0 1 89216
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1122
timestamp 1636968456
transform 1 0 104328 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1134
timestamp 1636968456
transform 1 0 105432 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_1146
timestamp 1
transform 1 0 106536 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1148
timestamp 1636968456
transform 1 0 106720 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_160_1160
timestamp 1
transform 1 0 107824 0 1 89216
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_161_3
timestamp 1636968456
transform 1 0 1380 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_15
timestamp 1636968456
transform 1 0 2484 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_27
timestamp 1636968456
transform 1 0 3588 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_39
timestamp 1636968456
transform 1 0 4692 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_161_51
timestamp 1
transform 1 0 5796 0 -1 90304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_161_55
timestamp 1
transform 1 0 6164 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_57
timestamp 1636968456
transform 1 0 6348 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_161_69
timestamp 1
transform 1 0 7452 0 -1 90304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1122
timestamp 1636968456
transform 1 0 104328 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1134
timestamp 1636968456
transform 1 0 105432 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1146
timestamp 1636968456
transform 1 0 106536 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_1158
timestamp 1
transform 1 0 107640 0 -1 90304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_161_1166
timestamp 1
transform 1 0 108376 0 -1 90304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_162_3
timestamp 1636968456
transform 1 0 1380 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_15
timestamp 1636968456
transform 1 0 2484 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_27
timestamp 1
transform 1 0 3588 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_29
timestamp 1636968456
transform 1 0 3772 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_41
timestamp 1636968456
transform 1 0 4876 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_53
timestamp 1636968456
transform 1 0 5980 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_65
timestamp 1
transform 1 0 7084 0 1 90304
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1122
timestamp 1636968456
transform 1 0 104328 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1134
timestamp 1636968456
transform 1 0 105432 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_1146
timestamp 1
transform 1 0 106536 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1148
timestamp 1636968456
transform 1 0 106720 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_162_1160
timestamp 1
transform 1 0 107824 0 1 90304
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_163_3
timestamp 1636968456
transform 1 0 1380 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_15
timestamp 1636968456
transform 1 0 2484 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_27
timestamp 1636968456
transform 1 0 3588 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_39
timestamp 1636968456
transform 1 0 4692 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_163_51
timestamp 1
transform 1 0 5796 0 -1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_163_55
timestamp 1
transform 1 0 6164 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_57
timestamp 1636968456
transform 1 0 6348 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_163_69
timestamp 1
transform 1 0 7452 0 -1 91392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1122
timestamp 1636968456
transform 1 0 104328 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1134
timestamp 1636968456
transform 1 0 105432 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1146
timestamp 1636968456
transform 1 0 106536 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_163_1158
timestamp 1
transform 1 0 107640 0 -1 91392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_163_1166
timestamp 1
transform 1 0 108376 0 -1 91392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_164_3
timestamp 1636968456
transform 1 0 1380 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_15
timestamp 1636968456
transform 1 0 2484 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_27
timestamp 1
transform 1 0 3588 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_29
timestamp 1636968456
transform 1 0 3772 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_41
timestamp 1636968456
transform 1 0 4876 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_53
timestamp 1636968456
transform 1 0 5980 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_65
timestamp 1
transform 1 0 7084 0 1 91392
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1122
timestamp 1636968456
transform 1 0 104328 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1134
timestamp 1636968456
transform 1 0 105432 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_1146
timestamp 1
transform 1 0 106536 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1148
timestamp 1636968456
transform 1 0 106720 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_164_1160
timestamp 1
transform 1 0 107824 0 1 91392
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_165_3
timestamp 1636968456
transform 1 0 1380 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_15
timestamp 1636968456
transform 1 0 2484 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_27
timestamp 1636968456
transform 1 0 3588 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_39
timestamp 1636968456
transform 1 0 4692 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_165_51
timestamp 1
transform 1 0 5796 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_165_55
timestamp 1
transform 1 0 6164 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_57
timestamp 1636968456
transform 1 0 6348 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_165_69
timestamp 1
transform 1 0 7452 0 -1 92480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1122
timestamp 1636968456
transform 1 0 104328 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1134
timestamp 1636968456
transform 1 0 105432 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1146
timestamp 1636968456
transform 1 0 106536 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_1158
timestamp 1
transform 1 0 107640 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_165_1166
timestamp 1
transform 1 0 108376 0 -1 92480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_166_3
timestamp 1636968456
transform 1 0 1380 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_15
timestamp 1636968456
transform 1 0 2484 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_27
timestamp 1
transform 1 0 3588 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_29
timestamp 1636968456
transform 1 0 3772 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_41
timestamp 1636968456
transform 1 0 4876 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_53
timestamp 1636968456
transform 1 0 5980 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_65
timestamp 1
transform 1 0 7084 0 1 92480
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1122
timestamp 1636968456
transform 1 0 104328 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1134
timestamp 1636968456
transform 1 0 105432 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_1146
timestamp 1
transform 1 0 106536 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1148
timestamp 1636968456
transform 1 0 106720 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_1160
timestamp 1
transform 1 0 107824 0 1 92480
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_167_3
timestamp 1636968456
transform 1 0 1380 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_15
timestamp 1636968456
transform 1 0 2484 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_27
timestamp 1636968456
transform 1 0 3588 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_39
timestamp 1636968456
transform 1 0 4692 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_167_51
timestamp 1
transform 1 0 5796 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_55
timestamp 1
transform 1 0 6164 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_57
timestamp 1636968456
transform 1 0 6348 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_167_69
timestamp 1
transform 1 0 7452 0 -1 93568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1122
timestamp 1636968456
transform 1 0 104328 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1134
timestamp 1636968456
transform 1 0 105432 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1146
timestamp 1636968456
transform 1 0 106536 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_1158
timestamp 1
transform 1 0 107640 0 -1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_167_1166
timestamp 1
transform 1 0 108376 0 -1 93568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_168_3
timestamp 1636968456
transform 1 0 1380 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_15
timestamp 1636968456
transform 1 0 2484 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_27
timestamp 1
transform 1 0 3588 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_29
timestamp 1636968456
transform 1 0 3772 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_41
timestamp 1636968456
transform 1 0 4876 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_53
timestamp 1636968456
transform 1 0 5980 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_65
timestamp 1
transform 1 0 7084 0 1 93568
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1122
timestamp 1636968456
transform 1 0 104328 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1134
timestamp 1636968456
transform 1 0 105432 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_1146
timestamp 1
transform 1 0 106536 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1148
timestamp 1636968456
transform 1 0 106720 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_168_1160
timestamp 1
transform 1 0 107824 0 1 93568
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_169_8
timestamp 1636968456
transform 1 0 1840 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_20
timestamp 1636968456
transform 1 0 2944 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_32
timestamp 1636968456
transform 1 0 4048 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_44
timestamp 1636968456
transform 1 0 5152 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_57
timestamp 1636968456
transform 1 0 6348 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_169_69
timestamp 1
transform 1 0 7452 0 -1 94656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1122
timestamp 1636968456
transform 1 0 104328 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1134
timestamp 1636968456
transform 1 0 105432 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1146
timestamp 1636968456
transform 1 0 106536 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_169_1158
timestamp 1
transform 1 0 107640 0 -1 94656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_169_1166
timestamp 1
transform 1 0 108376 0 -1 94656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_170_3
timestamp 1636968456
transform 1 0 1380 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_15
timestamp 1636968456
transform 1 0 2484 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_27
timestamp 1
transform 1 0 3588 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_29
timestamp 1636968456
transform 1 0 3772 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_41
timestamp 1636968456
transform 1 0 4876 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_53
timestamp 1636968456
transform 1 0 5980 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_65
timestamp 1
transform 1 0 7084 0 1 94656
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1122
timestamp 1636968456
transform 1 0 104328 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1134
timestamp 1636968456
transform 1 0 105432 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_1146
timestamp 1
transform 1 0 106536 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1148
timestamp 1636968456
transform 1 0 106720 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_170_1160
timestamp 1
transform 1 0 107824 0 1 94656
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_171_3
timestamp 1636968456
transform 1 0 1380 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_15
timestamp 1636968456
transform 1 0 2484 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_27
timestamp 1636968456
transform 1 0 3588 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_39
timestamp 1636968456
transform 1 0 4692 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_171_51
timestamp 1
transform 1 0 5796 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_171_55
timestamp 1
transform 1 0 6164 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_57
timestamp 1636968456
transform 1 0 6348 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_171_69
timestamp 1
transform 1 0 7452 0 -1 95744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1122
timestamp 1636968456
transform 1 0 104328 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1134
timestamp 1636968456
transform 1 0 105432 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1146
timestamp 1636968456
transform 1 0 106536 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_1158
timestamp 1
transform 1 0 107640 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_171_1166
timestamp 1
transform 1 0 108376 0 -1 95744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_172_8
timestamp 1636968456
transform 1 0 1840 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_20
timestamp 1
transform 1 0 2944 0 1 95744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_172_29
timestamp 1636968456
transform 1 0 3772 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_41
timestamp 1636968456
transform 1 0 4876 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_53
timestamp 1636968456
transform 1 0 5980 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_65
timestamp 1
transform 1 0 7084 0 1 95744
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1122
timestamp 1636968456
transform 1 0 104328 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1134
timestamp 1636968456
transform 1 0 105432 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_172_1146
timestamp 1
transform 1 0 106536 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1148
timestamp 1636968456
transform 1 0 106720 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_1160
timestamp 1
transform 1 0 107824 0 1 95744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_173_3
timestamp 1636968456
transform 1 0 1380 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_15
timestamp 1636968456
transform 1 0 2484 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_27
timestamp 1636968456
transform 1 0 3588 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_39
timestamp 1636968456
transform 1 0 4692 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_173_51
timestamp 1
transform 1 0 5796 0 -1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_173_55
timestamp 1
transform 1 0 6164 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_57
timestamp 1636968456
transform 1 0 6348 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_173_69
timestamp 1
transform 1 0 7452 0 -1 96832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1122
timestamp 1636968456
transform 1 0 104328 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1134
timestamp 1636968456
transform 1 0 105432 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1146
timestamp 1636968456
transform 1 0 106536 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_1158
timestamp 1
transform 1 0 107640 0 -1 96832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_173_1166
timestamp 1
transform 1 0 108376 0 -1 96832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_174_8
timestamp 1636968456
transform 1 0 1840 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_174_20
timestamp 1
transform 1 0 2944 0 1 96832
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_174_29
timestamp 1636968456
transform 1 0 3772 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_41
timestamp 1636968456
transform 1 0 4876 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_53
timestamp 1636968456
transform 1 0 5980 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_65
timestamp 1
transform 1 0 7084 0 1 96832
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1122
timestamp 1636968456
transform 1 0 104328 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1134
timestamp 1636968456
transform 1 0 105432 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_174_1146
timestamp 1
transform 1 0 106536 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1148
timestamp 1636968456
transform 1 0 106720 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_174_1160
timestamp 1
transform 1 0 107824 0 1 96832
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_175_3
timestamp 1636968456
transform 1 0 1380 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_15
timestamp 1636968456
transform 1 0 2484 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_27
timestamp 1636968456
transform 1 0 3588 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_39
timestamp 1636968456
transform 1 0 4692 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_175_51
timestamp 1
transform 1 0 5796 0 -1 97920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_175_55
timestamp 1
transform 1 0 6164 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_57
timestamp 1636968456
transform 1 0 6348 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_175_69
timestamp 1
transform 1 0 7452 0 -1 97920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1122
timestamp 1636968456
transform 1 0 104328 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1134
timestamp 1636968456
transform 1 0 105432 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1146
timestamp 1636968456
transform 1 0 106536 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_175_1158
timestamp 1
transform 1 0 107640 0 -1 97920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_175_1166
timestamp 1
transform 1 0 108376 0 -1 97920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_176_3
timestamp 1636968456
transform 1 0 1380 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_15
timestamp 1636968456
transform 1 0 2484 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_176_27
timestamp 1
transform 1 0 3588 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_29
timestamp 1636968456
transform 1 0 3772 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_41
timestamp 1636968456
transform 1 0 4876 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_53
timestamp 1636968456
transform 1 0 5980 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_65
timestamp 1
transform 1 0 7084 0 1 97920
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1122
timestamp 1636968456
transform 1 0 104328 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1134
timestamp 1636968456
transform 1 0 105432 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_176_1146
timestamp 1
transform 1 0 106536 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1148
timestamp 1636968456
transform 1 0 106720 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_176_1160
timestamp 1
transform 1 0 107824 0 1 97920
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_177_8
timestamp 1636968456
transform 1 0 1840 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_20
timestamp 1636968456
transform 1 0 2944 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_32
timestamp 1636968456
transform 1 0 4048 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_44
timestamp 1636968456
transform 1 0 5152 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_57
timestamp 1636968456
transform 1 0 6348 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_177_69
timestamp 1
transform 1 0 7452 0 -1 99008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1122
timestamp 1636968456
transform 1 0 104328 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1134
timestamp 1636968456
transform 1 0 105432 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1146
timestamp 1636968456
transform 1 0 106536 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_177_1158
timestamp 1
transform 1 0 107640 0 -1 99008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_177_1166
timestamp 1
transform 1 0 108376 0 -1 99008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_178_3
timestamp 1636968456
transform 1 0 1380 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_15
timestamp 1636968456
transform 1 0 2484 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_178_27
timestamp 1
transform 1 0 3588 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_29
timestamp 1636968456
transform 1 0 3772 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_41
timestamp 1636968456
transform 1 0 4876 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_53
timestamp 1636968456
transform 1 0 5980 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_65
timestamp 1
transform 1 0 7084 0 1 99008
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1122
timestamp 1636968456
transform 1 0 104328 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1134
timestamp 1636968456
transform 1 0 105432 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_178_1146
timestamp 1
transform 1 0 106536 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1148
timestamp 1636968456
transform 1 0 106720 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_178_1160
timestamp 1
transform 1 0 107824 0 1 99008
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_179_8
timestamp 1636968456
transform 1 0 1840 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_20
timestamp 1636968456
transform 1 0 2944 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_32
timestamp 1636968456
transform 1 0 4048 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_44
timestamp 1636968456
transform 1 0 5152 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_57
timestamp 1636968456
transform 1 0 6348 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_179_69
timestamp 1
transform 1 0 7452 0 -1 100096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1122
timestamp 1636968456
transform 1 0 104328 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1134
timestamp 1636968456
transform 1 0 105432 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1146
timestamp 1636968456
transform 1 0 106536 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_1158
timestamp 1
transform 1 0 107640 0 -1 100096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_179_1166
timestamp 1
transform 1 0 108376 0 -1 100096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_180_3
timestamp 1636968456
transform 1 0 1380 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_15
timestamp 1636968456
transform 1 0 2484 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_180_27
timestamp 1
transform 1 0 3588 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_29
timestamp 1636968456
transform 1 0 3772 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_41
timestamp 1636968456
transform 1 0 4876 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_53
timestamp 1636968456
transform 1 0 5980 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_65
timestamp 1
transform 1 0 7084 0 1 100096
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1122
timestamp 1636968456
transform 1 0 104328 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1134
timestamp 1636968456
transform 1 0 105432 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_180_1146
timestamp 1
transform 1 0 106536 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1148
timestamp 1636968456
transform 1 0 106720 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_180_1160
timestamp 1
transform 1 0 107824 0 1 100096
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_181_3
timestamp 1636968456
transform 1 0 1380 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_15
timestamp 1636968456
transform 1 0 2484 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_27
timestamp 1636968456
transform 1 0 3588 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_39
timestamp 1636968456
transform 1 0 4692 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_181_51
timestamp 1
transform 1 0 5796 0 -1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_181_55
timestamp 1
transform 1 0 6164 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_57
timestamp 1636968456
transform 1 0 6348 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_181_69
timestamp 1
transform 1 0 7452 0 -1 101184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1122
timestamp 1636968456
transform 1 0 104328 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1134
timestamp 1636968456
transform 1 0 105432 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1146
timestamp 1636968456
transform 1 0 106536 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_181_1158
timestamp 1
transform 1 0 107640 0 -1 101184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_181_1166
timestamp 1
transform 1 0 108376 0 -1 101184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_182_8
timestamp 1636968456
transform 1 0 1840 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_182_20
timestamp 1
transform 1 0 2944 0 1 101184
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_182_29
timestamp 1636968456
transform 1 0 3772 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_41
timestamp 1636968456
transform 1 0 4876 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_53
timestamp 1636968456
transform 1 0 5980 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_65
timestamp 1
transform 1 0 7084 0 1 101184
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1122
timestamp 1636968456
transform 1 0 104328 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1134
timestamp 1636968456
transform 1 0 105432 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_182_1146
timestamp 1
transform 1 0 106536 0 1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1148
timestamp 1636968456
transform 1 0 106720 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_182_1160
timestamp 1
transform 1 0 107824 0 1 101184
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_183_3
timestamp 1636968456
transform 1 0 1380 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_15
timestamp 1636968456
transform 1 0 2484 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_27
timestamp 1636968456
transform 1 0 3588 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_39
timestamp 1636968456
transform 1 0 4692 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_183_51
timestamp 1
transform 1 0 5796 0 -1 102272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_183_55
timestamp 1
transform 1 0 6164 0 -1 102272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_183_57
timestamp 1636968456
transform 1 0 6348 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_183_69
timestamp 1
transform 1 0 7452 0 -1 102272
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_183_1122
timestamp 1636968456
transform 1 0 104328 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_1134
timestamp 1636968456
transform 1 0 105432 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_1146
timestamp 1636968456
transform 1 0 106536 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_183_1158
timestamp 1
transform 1 0 107640 0 -1 102272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_183_1166
timestamp 1
transform 1 0 108376 0 -1 102272
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_184_3
timestamp 1636968456
transform 1 0 1380 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_15
timestamp 1636968456
transform 1 0 2484 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_184_27
timestamp 1
transform 1 0 3588 0 1 102272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_184_29
timestamp 1636968456
transform 1 0 3772 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_41
timestamp 1636968456
transform 1 0 4876 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_53
timestamp 1636968456
transform 1 0 5980 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_65
timestamp 1
transform 1 0 7084 0 1 102272
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_184_1122
timestamp 1636968456
transform 1 0 104328 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_1134
timestamp 1636968456
transform 1 0 105432 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_184_1146
timestamp 1
transform 1 0 106536 0 1 102272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_184_1148
timestamp 1636968456
transform 1 0 106720 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_184_1160
timestamp 1
transform 1 0 107824 0 1 102272
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_185_3
timestamp 1636968456
transform 1 0 1380 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_15
timestamp 1636968456
transform 1 0 2484 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_27
timestamp 1636968456
transform 1 0 3588 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_39
timestamp 1636968456
transform 1 0 4692 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_185_51
timestamp 1
transform 1 0 5796 0 -1 103360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_185_55
timestamp 1
transform 1 0 6164 0 -1 103360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_185_57
timestamp 1636968456
transform 1 0 6348 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_185_69
timestamp 1
transform 1 0 7452 0 -1 103360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_185_1122
timestamp 1636968456
transform 1 0 104328 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_1134
timestamp 1636968456
transform 1 0 105432 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_1146
timestamp 1636968456
transform 1 0 106536 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_185_1158
timestamp 1
transform 1 0 107640 0 -1 103360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_185_1166
timestamp 1
transform 1 0 108376 0 -1 103360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_186_3
timestamp 1636968456
transform 1 0 1380 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_15
timestamp 1636968456
transform 1 0 2484 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_186_27
timestamp 1
transform 1 0 3588 0 1 103360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_186_29
timestamp 1636968456
transform 1 0 3772 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_41
timestamp 1636968456
transform 1 0 4876 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_53
timestamp 1636968456
transform 1 0 5980 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_65
timestamp 1
transform 1 0 7084 0 1 103360
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_186_1122
timestamp 1636968456
transform 1 0 104328 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_1134
timestamp 1636968456
transform 1 0 105432 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_186_1146
timestamp 1
transform 1 0 106536 0 1 103360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_186_1148
timestamp 1636968456
transform 1 0 106720 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_1160
timestamp 1
transform 1 0 107824 0 1 103360
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_187_3
timestamp 1636968456
transform 1 0 1380 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_15
timestamp 1636968456
transform 1 0 2484 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_27
timestamp 1636968456
transform 1 0 3588 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_39
timestamp 1636968456
transform 1 0 4692 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_187_51
timestamp 1
transform 1 0 5796 0 -1 104448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_187_55
timestamp 1
transform 1 0 6164 0 -1 104448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_187_57
timestamp 1636968456
transform 1 0 6348 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_187_69
timestamp 1
transform 1 0 7452 0 -1 104448
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_187_1122
timestamp 1636968456
transform 1 0 104328 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_1134
timestamp 1636968456
transform 1 0 105432 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_1146
timestamp 1636968456
transform 1 0 106536 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_187_1158
timestamp 1
transform 1 0 107640 0 -1 104448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_187_1166
timestamp 1
transform 1 0 108376 0 -1 104448
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_188_3
timestamp 1636968456
transform 1 0 1380 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_15
timestamp 1636968456
transform 1 0 2484 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_188_27
timestamp 1
transform 1 0 3588 0 1 104448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_188_29
timestamp 1636968456
transform 1 0 3772 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_41
timestamp 1636968456
transform 1 0 4876 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_53
timestamp 1636968456
transform 1 0 5980 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_65
timestamp 1
transform 1 0 7084 0 1 104448
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_188_1122
timestamp 1636968456
transform 1 0 104328 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_1134
timestamp 1636968456
transform 1 0 105432 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_188_1146
timestamp 1
transform 1 0 106536 0 1 104448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_188_1148
timestamp 1636968456
transform 1 0 106720 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_188_1160
timestamp 1
transform 1 0 107824 0 1 104448
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_189_3
timestamp 1636968456
transform 1 0 1380 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_15
timestamp 1636968456
transform 1 0 2484 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_27
timestamp 1636968456
transform 1 0 3588 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_39
timestamp 1636968456
transform 1 0 4692 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_189_51
timestamp 1
transform 1 0 5796 0 -1 105536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_189_55
timestamp 1
transform 1 0 6164 0 -1 105536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_189_57
timestamp 1636968456
transform 1 0 6348 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_189_69
timestamp 1
transform 1 0 7452 0 -1 105536
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_189_1122
timestamp 1636968456
transform 1 0 104328 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_1134
timestamp 1636968456
transform 1 0 105432 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_1146
timestamp 1636968456
transform 1 0 106536 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_189_1158
timestamp 1
transform 1 0 107640 0 -1 105536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_189_1166
timestamp 1
transform 1 0 108376 0 -1 105536
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_190_3
timestamp 1636968456
transform 1 0 1380 0 1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_190_15
timestamp 1636968456
transform 1 0 2484 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_190_27
timestamp 1
transform 1 0 3588 0 1 105536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_190_29
timestamp 1636968456
transform 1 0 3772 0 1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_190_41
timestamp 1636968456
transform 1 0 4876 0 1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_190_53
timestamp 1636968456
transform 1 0 5980 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_65
timestamp 1
transform 1 0 7084 0 1 105536
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_190_1122
timestamp 1636968456
transform 1 0 104328 0 1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_190_1134
timestamp 1636968456
transform 1 0 105432 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_190_1146
timestamp 1
transform 1 0 106536 0 1 105536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_190_1148
timestamp 1636968456
transform 1 0 106720 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_190_1160
timestamp 1
transform 1 0 107824 0 1 105536
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_191_3
timestamp 1636968456
transform 1 0 1380 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_15
timestamp 1636968456
transform 1 0 2484 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_27
timestamp 1636968456
transform 1 0 3588 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_39
timestamp 1636968456
transform 1 0 4692 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_191_51
timestamp 1
transform 1 0 5796 0 -1 106624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_191_55
timestamp 1
transform 1 0 6164 0 -1 106624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_191_57
timestamp 1636968456
transform 1 0 6348 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_191_69
timestamp 1
transform 1 0 7452 0 -1 106624
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_191_1122
timestamp 1636968456
transform 1 0 104328 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_1134
timestamp 1636968456
transform 1 0 105432 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_1146
timestamp 1636968456
transform 1 0 106536 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_191_1158
timestamp 1
transform 1 0 107640 0 -1 106624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_191_1166
timestamp 1
transform 1 0 108376 0 -1 106624
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_192_3
timestamp 1636968456
transform 1 0 1380 0 1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_192_15
timestamp 1636968456
transform 1 0 2484 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_192_27
timestamp 1
transform 1 0 3588 0 1 106624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_192_29
timestamp 1636968456
transform 1 0 3772 0 1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_192_41
timestamp 1636968456
transform 1 0 4876 0 1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_192_53
timestamp 1636968456
transform 1 0 5980 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_65
timestamp 1
transform 1 0 7084 0 1 106624
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_192_1122
timestamp 1636968456
transform 1 0 104328 0 1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_192_1134
timestamp 1636968456
transform 1 0 105432 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_192_1146
timestamp 1
transform 1 0 106536 0 1 106624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_192_1148
timestamp 1636968456
transform 1 0 106720 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_1160
timestamp 1
transform 1 0 107824 0 1 106624
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_193_3
timestamp 1636968456
transform 1 0 1380 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_15
timestamp 1636968456
transform 1 0 2484 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_27
timestamp 1636968456
transform 1 0 3588 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_39
timestamp 1636968456
transform 1 0 4692 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_193_51
timestamp 1
transform 1 0 5796 0 -1 107712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_193_55
timestamp 1
transform 1 0 6164 0 -1 107712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_193_57
timestamp 1636968456
transform 1 0 6348 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_193_69
timestamp 1
transform 1 0 7452 0 -1 107712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_193_1122
timestamp 1636968456
transform 1 0 104328 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_1134
timestamp 1636968456
transform 1 0 105432 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_1146
timestamp 1636968456
transform 1 0 106536 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_193_1158
timestamp 1
transform 1 0 107640 0 -1 107712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_193_1166
timestamp 1
transform 1 0 108376 0 -1 107712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_194_3
timestamp 1636968456
transform 1 0 1380 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_15
timestamp 1636968456
transform 1 0 2484 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_194_27
timestamp 1
transform 1 0 3588 0 1 107712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_194_29
timestamp 1636968456
transform 1 0 3772 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_41
timestamp 1636968456
transform 1 0 4876 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_53
timestamp 1636968456
transform 1 0 5980 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_65
timestamp 1
transform 1 0 7084 0 1 107712
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_194_1122
timestamp 1636968456
transform 1 0 104328 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_1134
timestamp 1636968456
transform 1 0 105432 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_194_1146
timestamp 1
transform 1 0 106536 0 1 107712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_194_1148
timestamp 1636968456
transform 1 0 106720 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_194_1160
timestamp 1
transform 1 0 107824 0 1 107712
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_195_3
timestamp 1636968456
transform 1 0 1380 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_15
timestamp 1636968456
transform 1 0 2484 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_27
timestamp 1636968456
transform 1 0 3588 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_39
timestamp 1636968456
transform 1 0 4692 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_195_51
timestamp 1
transform 1 0 5796 0 -1 108800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_195_55
timestamp 1
transform 1 0 6164 0 -1 108800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_195_57
timestamp 1636968456
transform 1 0 6348 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_195_69
timestamp 1
transform 1 0 7452 0 -1 108800
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_195_1122
timestamp 1636968456
transform 1 0 104328 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_1134
timestamp 1636968456
transform 1 0 105432 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_1146
timestamp 1636968456
transform 1 0 106536 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_195_1158
timestamp 1
transform 1 0 107640 0 -1 108800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_195_1166
timestamp 1
transform 1 0 108376 0 -1 108800
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_196_3
timestamp 1636968456
transform 1 0 1380 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_15
timestamp 1636968456
transform 1 0 2484 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_196_27
timestamp 1
transform 1 0 3588 0 1 108800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_196_29
timestamp 1636968456
transform 1 0 3772 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_41
timestamp 1636968456
transform 1 0 4876 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_53
timestamp 1636968456
transform 1 0 5980 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_65
timestamp 1
transform 1 0 7084 0 1 108800
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_196_1122
timestamp 1636968456
transform 1 0 104328 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_1134
timestamp 1636968456
transform 1 0 105432 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_196_1146
timestamp 1
transform 1 0 106536 0 1 108800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_196_1148
timestamp 1636968456
transform 1 0 106720 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_196_1160
timestamp 1
transform 1 0 107824 0 1 108800
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_197_3
timestamp 1636968456
transform 1 0 1380 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_15
timestamp 1636968456
transform 1 0 2484 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_27
timestamp 1636968456
transform 1 0 3588 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_39
timestamp 1636968456
transform 1 0 4692 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_197_51
timestamp 1
transform 1 0 5796 0 -1 109888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_197_55
timestamp 1
transform 1 0 6164 0 -1 109888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_197_57
timestamp 1636968456
transform 1 0 6348 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_197_69
timestamp 1
transform 1 0 7452 0 -1 109888
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_197_1122
timestamp 1636968456
transform 1 0 104328 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_1134
timestamp 1636968456
transform 1 0 105432 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_1146
timestamp 1636968456
transform 1 0 106536 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_197_1158
timestamp 1
transform 1 0 107640 0 -1 109888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_197_1166
timestamp 1
transform 1 0 108376 0 -1 109888
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_198_3
timestamp 1636968456
transform 1 0 1380 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_15
timestamp 1636968456
transform 1 0 2484 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_198_27
timestamp 1
transform 1 0 3588 0 1 109888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_198_29
timestamp 1636968456
transform 1 0 3772 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_41
timestamp 1636968456
transform 1 0 4876 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_53
timestamp 1636968456
transform 1 0 5980 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_65
timestamp 1
transform 1 0 7084 0 1 109888
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_198_1122
timestamp 1636968456
transform 1 0 104328 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_1134
timestamp 1636968456
transform 1 0 105432 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_198_1146
timestamp 1
transform 1 0 106536 0 1 109888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_198_1148
timestamp 1636968456
transform 1 0 106720 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_198_1160
timestamp 1
transform 1 0 107824 0 1 109888
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_199_3
timestamp 1636968456
transform 1 0 1380 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_15
timestamp 1636968456
transform 1 0 2484 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_27
timestamp 1636968456
transform 1 0 3588 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_39
timestamp 1636968456
transform 1 0 4692 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_199_51
timestamp 1
transform 1 0 5796 0 -1 110976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_199_55
timestamp 1
transform 1 0 6164 0 -1 110976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_199_57
timestamp 1636968456
transform 1 0 6348 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_199_69
timestamp 1
transform 1 0 7452 0 -1 110976
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_199_1122
timestamp 1636968456
transform 1 0 104328 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_1134
timestamp 1636968456
transform 1 0 105432 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_1146
timestamp 1636968456
transform 1 0 106536 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_1158
timestamp 1
transform 1 0 107640 0 -1 110976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_199_1166
timestamp 1
transform 1 0 108376 0 -1 110976
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_200_3
timestamp 1636968456
transform 1 0 1380 0 1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_200_15
timestamp 1636968456
transform 1 0 2484 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_200_27
timestamp 1
transform 1 0 3588 0 1 110976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_200_29
timestamp 1636968456
transform 1 0 3772 0 1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_200_41
timestamp 1636968456
transform 1 0 4876 0 1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_200_53
timestamp 1636968456
transform 1 0 5980 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_65
timestamp 1
transform 1 0 7084 0 1 110976
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_200_1122
timestamp 1636968456
transform 1 0 104328 0 1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_200_1134
timestamp 1636968456
transform 1 0 105432 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_200_1146
timestamp 1
transform 1 0 106536 0 1 110976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_200_1148
timestamp 1636968456
transform 1 0 106720 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_200_1160
timestamp 1
transform 1 0 107824 0 1 110976
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_201_3
timestamp 1636968456
transform 1 0 1380 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_15
timestamp 1636968456
transform 1 0 2484 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_27
timestamp 1636968456
transform 1 0 3588 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_39
timestamp 1636968456
transform 1 0 4692 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_201_51
timestamp 1
transform 1 0 5796 0 -1 112064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_201_55
timestamp 1
transform 1 0 6164 0 -1 112064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_201_57
timestamp 1636968456
transform 1 0 6348 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_201_69
timestamp 1
transform 1 0 7452 0 -1 112064
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_201_1122
timestamp 1636968456
transform 1 0 104328 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_1134
timestamp 1636968456
transform 1 0 105432 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_1146
timestamp 1636968456
transform 1 0 106536 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_201_1158
timestamp 1
transform 1 0 107640 0 -1 112064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_201_1166
timestamp 1
transform 1 0 108376 0 -1 112064
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_202_3
timestamp 1636968456
transform 1 0 1380 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_15
timestamp 1636968456
transform 1 0 2484 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_202_27
timestamp 1
transform 1 0 3588 0 1 112064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_202_29
timestamp 1636968456
transform 1 0 3772 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_41
timestamp 1636968456
transform 1 0 4876 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_53
timestamp 1636968456
transform 1 0 5980 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_65
timestamp 1
transform 1 0 7084 0 1 112064
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_202_1122
timestamp 1636968456
transform 1 0 104328 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_1134
timestamp 1636968456
transform 1 0 105432 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_202_1146
timestamp 1
transform 1 0 106536 0 1 112064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_202_1148
timestamp 1636968456
transform 1 0 106720 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_202_1160
timestamp 1
transform 1 0 107824 0 1 112064
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_203_3
timestamp 1636968456
transform 1 0 1380 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_15
timestamp 1636968456
transform 1 0 2484 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_27
timestamp 1636968456
transform 1 0 3588 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_39
timestamp 1636968456
transform 1 0 4692 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_203_51
timestamp 1
transform 1 0 5796 0 -1 113152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_203_55
timestamp 1
transform 1 0 6164 0 -1 113152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_203_57
timestamp 1636968456
transform 1 0 6348 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_203_69
timestamp 1
transform 1 0 7452 0 -1 113152
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_203_1122
timestamp 1636968456
transform 1 0 104328 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_1134
timestamp 1636968456
transform 1 0 105432 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_1146
timestamp 1636968456
transform 1 0 106536 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_203_1158
timestamp 1
transform 1 0 107640 0 -1 113152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_203_1166
timestamp 1
transform 1 0 108376 0 -1 113152
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_204_3
timestamp 1636968456
transform 1 0 1380 0 1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_204_15
timestamp 1636968456
transform 1 0 2484 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_204_27
timestamp 1
transform 1 0 3588 0 1 113152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_204_29
timestamp 1636968456
transform 1 0 3772 0 1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_204_41
timestamp 1636968456
transform 1 0 4876 0 1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_204_53
timestamp 1636968456
transform 1 0 5980 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_65
timestamp 1
transform 1 0 7084 0 1 113152
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_204_1122
timestamp 1636968456
transform 1 0 104328 0 1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_204_1134
timestamp 1636968456
transform 1 0 105432 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_204_1146
timestamp 1
transform 1 0 106536 0 1 113152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_204_1148
timestamp 1636968456
transform 1 0 106720 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_204_1160
timestamp 1
transform 1 0 107824 0 1 113152
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_205_3
timestamp 1636968456
transform 1 0 1380 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_15
timestamp 1636968456
transform 1 0 2484 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_27
timestamp 1636968456
transform 1 0 3588 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_39
timestamp 1636968456
transform 1 0 4692 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_205_51
timestamp 1
transform 1 0 5796 0 -1 114240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_205_55
timestamp 1
transform 1 0 6164 0 -1 114240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_205_57
timestamp 1636968456
transform 1 0 6348 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_205_69
timestamp 1
transform 1 0 7452 0 -1 114240
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_205_1122
timestamp 1636968456
transform 1 0 104328 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_1134
timestamp 1636968456
transform 1 0 105432 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_1146
timestamp 1636968456
transform 1 0 106536 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_205_1158
timestamp 1
transform 1 0 107640 0 -1 114240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_205_1166
timestamp 1
transform 1 0 108376 0 -1 114240
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_206_3
timestamp 1636968456
transform 1 0 1380 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_15
timestamp 1636968456
transform 1 0 2484 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_206_27
timestamp 1
transform 1 0 3588 0 1 114240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_206_29
timestamp 1636968456
transform 1 0 3772 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_41
timestamp 1636968456
transform 1 0 4876 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_53
timestamp 1636968456
transform 1 0 5980 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_65
timestamp 1
transform 1 0 7084 0 1 114240
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_206_1122
timestamp 1636968456
transform 1 0 104328 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_1134
timestamp 1636968456
transform 1 0 105432 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_206_1146
timestamp 1
transform 1 0 106536 0 1 114240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_206_1148
timestamp 1636968456
transform 1 0 106720 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_206_1160
timestamp 1
transform 1 0 107824 0 1 114240
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_207_3
timestamp 1636968456
transform 1 0 1380 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_15
timestamp 1636968456
transform 1 0 2484 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_27
timestamp 1636968456
transform 1 0 3588 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_39
timestamp 1636968456
transform 1 0 4692 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_207_51
timestamp 1
transform 1 0 5796 0 -1 115328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_55
timestamp 1
transform 1 0 6164 0 -1 115328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_207_57
timestamp 1636968456
transform 1 0 6348 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_207_69
timestamp 1
transform 1 0 7452 0 -1 115328
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_207_1122
timestamp 1636968456
transform 1 0 104328 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_1134
timestamp 1636968456
transform 1 0 105432 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_1146
timestamp 1636968456
transform 1 0 106536 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_207_1158
timestamp 1
transform 1 0 107640 0 -1 115328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_207_1166
timestamp 1
transform 1 0 108376 0 -1 115328
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_208_3
timestamp 1636968456
transform 1 0 1380 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_15
timestamp 1636968456
transform 1 0 2484 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_208_27
timestamp 1
transform 1 0 3588 0 1 115328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_208_29
timestamp 1636968456
transform 1 0 3772 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_41
timestamp 1636968456
transform 1 0 4876 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_53
timestamp 1636968456
transform 1 0 5980 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_65
timestamp 1
transform 1 0 7084 0 1 115328
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_208_1122
timestamp 1636968456
transform 1 0 104328 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_1134
timestamp 1636968456
transform 1 0 105432 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_208_1146
timestamp 1
transform 1 0 106536 0 1 115328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_208_1148
timestamp 1636968456
transform 1 0 106720 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_208_1160
timestamp 1
transform 1 0 107824 0 1 115328
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_209_3
timestamp 1636968456
transform 1 0 1380 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_15
timestamp 1636968456
transform 1 0 2484 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_27
timestamp 1636968456
transform 1 0 3588 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_39
timestamp 1636968456
transform 1 0 4692 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_209_51
timestamp 1
transform 1 0 5796 0 -1 116416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_55
timestamp 1
transform 1 0 6164 0 -1 116416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_209_57
timestamp 1636968456
transform 1 0 6348 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_209_69
timestamp 1
transform 1 0 7452 0 -1 116416
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_209_1122
timestamp 1636968456
transform 1 0 104328 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_1134
timestamp 1636968456
transform 1 0 105432 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_1146
timestamp 1636968456
transform 1 0 106536 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_209_1158
timestamp 1
transform 1 0 107640 0 -1 116416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_209_1166
timestamp 1
transform 1 0 108376 0 -1 116416
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_210_3
timestamp 1636968456
transform 1 0 1380 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_15
timestamp 1636968456
transform 1 0 2484 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_210_27
timestamp 1
transform 1 0 3588 0 1 116416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_210_29
timestamp 1636968456
transform 1 0 3772 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_41
timestamp 1636968456
transform 1 0 4876 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_53
timestamp 1636968456
transform 1 0 5980 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_65
timestamp 1
transform 1 0 7084 0 1 116416
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_210_1122
timestamp 1636968456
transform 1 0 104328 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_1134
timestamp 1636968456
transform 1 0 105432 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_210_1146
timestamp 1
transform 1 0 106536 0 1 116416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_210_1148
timestamp 1636968456
transform 1 0 106720 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_210_1160
timestamp 1
transform 1 0 107824 0 1 116416
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_211_3
timestamp 1636968456
transform 1 0 1380 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_15
timestamp 1636968456
transform 1 0 2484 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_27
timestamp 1636968456
transform 1 0 3588 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_39
timestamp 1636968456
transform 1 0 4692 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_211_51
timestamp 1
transform 1 0 5796 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_211_55
timestamp 1
transform 1 0 6164 0 -1 117504
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_211_57
timestamp 1636968456
transform 1 0 6348 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_211_69
timestamp 1
transform 1 0 7452 0 -1 117504
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_211_1122
timestamp 1636968456
transform 1 0 104328 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_1134
timestamp 1636968456
transform 1 0 105432 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_1146
timestamp 1636968456
transform 1 0 106536 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_211_1158
timestamp 1
transform 1 0 107640 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_211_1166
timestamp 1
transform 1 0 108376 0 -1 117504
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_212_3
timestamp 1636968456
transform 1 0 1380 0 1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_212_15
timestamp 1636968456
transform 1 0 2484 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_212_27
timestamp 1
transform 1 0 3588 0 1 117504
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_212_29
timestamp 1636968456
transform 1 0 3772 0 1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_212_41
timestamp 1636968456
transform 1 0 4876 0 1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_212_53
timestamp 1636968456
transform 1 0 5980 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_212_65
timestamp 1
transform 1 0 7084 0 1 117504
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_212_1122
timestamp 1636968456
transform 1 0 104328 0 1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_212_1134
timestamp 1636968456
transform 1 0 105432 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_212_1146
timestamp 1
transform 1 0 106536 0 1 117504
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_212_1148
timestamp 1636968456
transform 1 0 106720 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_212_1160
timestamp 1
transform 1 0 107824 0 1 117504
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_213_3
timestamp 1636968456
transform 1 0 1380 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_15
timestamp 1636968456
transform 1 0 2484 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_27
timestamp 1636968456
transform 1 0 3588 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_39
timestamp 1636968456
transform 1 0 4692 0 -1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_213_51
timestamp 1
transform 1 0 5796 0 -1 118592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_213_55
timestamp 1
transform 1 0 6164 0 -1 118592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_213_57
timestamp 1636968456
transform 1 0 6348 0 -1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_213_69
timestamp 1
transform 1 0 7452 0 -1 118592
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_213_1122
timestamp 1636968456
transform 1 0 104328 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_1134
timestamp 1636968456
transform 1 0 105432 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_1146
timestamp 1636968456
transform 1 0 106536 0 -1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_213_1158
timestamp 1
transform 1 0 107640 0 -1 118592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_213_1166
timestamp 1
transform 1 0 108376 0 -1 118592
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_214_3
timestamp 1636968456
transform 1 0 1380 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_15
timestamp 1636968456
transform 1 0 2484 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_214_27
timestamp 1
transform 1 0 3588 0 1 118592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_214_29
timestamp 1636968456
transform 1 0 3772 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_41
timestamp 1636968456
transform 1 0 4876 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_53
timestamp 1636968456
transform 1 0 5980 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_214_65
timestamp 1
transform 1 0 7084 0 1 118592
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_214_1122
timestamp 1636968456
transform 1 0 104328 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_1134
timestamp 1636968456
transform 1 0 105432 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_214_1146
timestamp 1
transform 1 0 106536 0 1 118592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_214_1148
timestamp 1636968456
transform 1 0 106720 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_214_1160
timestamp 1
transform 1 0 107824 0 1 118592
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_215_3
timestamp 1636968456
transform 1 0 1380 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_15
timestamp 1636968456
transform 1 0 2484 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_27
timestamp 1636968456
transform 1 0 3588 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_39
timestamp 1636968456
transform 1 0 4692 0 -1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_215_51
timestamp 1
transform 1 0 5796 0 -1 119680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_215_55
timestamp 1
transform 1 0 6164 0 -1 119680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_215_57
timestamp 1636968456
transform 1 0 6348 0 -1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_215_69
timestamp 1
transform 1 0 7452 0 -1 119680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_215_1122
timestamp 1636968456
transform 1 0 104328 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_1134
timestamp 1636968456
transform 1 0 105432 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_1146
timestamp 1636968456
transform 1 0 106536 0 -1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_215_1158
timestamp 1
transform 1 0 107640 0 -1 119680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_215_1166
timestamp 1
transform 1 0 108376 0 -1 119680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_216_3
timestamp 1636968456
transform 1 0 1380 0 1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_216_15
timestamp 1636968456
transform 1 0 2484 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_216_27
timestamp 1
transform 1 0 3588 0 1 119680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_216_29
timestamp 1636968456
transform 1 0 3772 0 1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_216_41
timestamp 1636968456
transform 1 0 4876 0 1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_216_53
timestamp 1636968456
transform 1 0 5980 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_216_65
timestamp 1
transform 1 0 7084 0 1 119680
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_216_1125
timestamp 1636968456
transform 1 0 104604 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_216_1137
timestamp 1
transform 1 0 105708 0 1 119680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_216_1145
timestamp 1
transform 1 0 106444 0 1 119680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_216_1148
timestamp 1636968456
transform 1 0 106720 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_216_1160
timestamp 1
transform 1 0 107824 0 1 119680
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_217_3
timestamp 1636968456
transform 1 0 1380 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_15
timestamp 1636968456
transform 1 0 2484 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_27
timestamp 1636968456
transform 1 0 3588 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_39
timestamp 1636968456
transform 1 0 4692 0 -1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_217_51
timestamp 1
transform 1 0 5796 0 -1 120768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_217_55
timestamp 1
transform 1 0 6164 0 -1 120768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_217_57
timestamp 1636968456
transform 1 0 6348 0 -1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_217_69
timestamp 1
transform 1 0 7452 0 -1 120768
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_217_1122
timestamp 1636968456
transform 1 0 104328 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_1134
timestamp 1636968456
transform 1 0 105432 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_1146
timestamp 1636968456
transform 1 0 106536 0 -1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_217_1158
timestamp 1
transform 1 0 107640 0 -1 120768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_217_1166
timestamp 1
transform 1 0 108376 0 -1 120768
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_218_3
timestamp 1636968456
transform 1 0 1380 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_15
timestamp 1636968456
transform 1 0 2484 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_218_27
timestamp 1
transform 1 0 3588 0 1 120768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_218_29
timestamp 1636968456
transform 1 0 3772 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_41
timestamp 1636968456
transform 1 0 4876 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_53
timestamp 1636968456
transform 1 0 5980 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_218_65
timestamp 1
transform 1 0 7084 0 1 120768
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_218_1122
timestamp 1636968456
transform 1 0 104328 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_1134
timestamp 1636968456
transform 1 0 105432 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_218_1146
timestamp 1
transform 1 0 106536 0 1 120768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_218_1148
timestamp 1636968456
transform 1 0 106720 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_218_1160
timestamp 1
transform 1 0 107824 0 1 120768
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_219_3
timestamp 1636968456
transform 1 0 1380 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_15
timestamp 1636968456
transform 1 0 2484 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_27
timestamp 1636968456
transform 1 0 3588 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_39
timestamp 1636968456
transform 1 0 4692 0 -1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_219_51
timestamp 1
transform 1 0 5796 0 -1 121856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_219_55
timestamp 1
transform 1 0 6164 0 -1 121856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_219_57
timestamp 1636968456
transform 1 0 6348 0 -1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_219_69
timestamp 1
transform 1 0 7452 0 -1 121856
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_219_1122
timestamp 1636968456
transform 1 0 104328 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_1134
timestamp 1636968456
transform 1 0 105432 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_1146
timestamp 1636968456
transform 1 0 106536 0 -1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_219_1158
timestamp 1
transform 1 0 107640 0 -1 121856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_219_1166
timestamp 1
transform 1 0 108376 0 -1 121856
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_220_3
timestamp 1636968456
transform 1 0 1380 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_15
timestamp 1636968456
transform 1 0 2484 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_220_27
timestamp 1
transform 1 0 3588 0 1 121856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_220_29
timestamp 1636968456
transform 1 0 3772 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_41
timestamp 1636968456
transform 1 0 4876 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_53
timestamp 1636968456
transform 1 0 5980 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_220_65
timestamp 1
transform 1 0 7084 0 1 121856
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_220_1122
timestamp 1636968456
transform 1 0 104328 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_1134
timestamp 1636968456
transform 1 0 105432 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_220_1146
timestamp 1
transform 1 0 106536 0 1 121856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_220_1148
timestamp 1636968456
transform 1 0 106720 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_220_1160
timestamp 1
transform 1 0 107824 0 1 121856
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_221_3
timestamp 1636968456
transform 1 0 1380 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_15
timestamp 1636968456
transform 1 0 2484 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_27
timestamp 1636968456
transform 1 0 3588 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_39
timestamp 1636968456
transform 1 0 4692 0 -1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_221_51
timestamp 1
transform 1 0 5796 0 -1 122944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_221_55
timestamp 1
transform 1 0 6164 0 -1 122944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_221_57
timestamp 1636968456
transform 1 0 6348 0 -1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_221_69
timestamp 1
transform 1 0 7452 0 -1 122944
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_221_1122
timestamp 1636968456
transform 1 0 104328 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_1134
timestamp 1636968456
transform 1 0 105432 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_1146
timestamp 1636968456
transform 1 0 106536 0 -1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_221_1158
timestamp 1
transform 1 0 107640 0 -1 122944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_221_1166
timestamp 1
transform 1 0 108376 0 -1 122944
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_222_3
timestamp 1636968456
transform 1 0 1380 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_15
timestamp 1636968456
transform 1 0 2484 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_222_27
timestamp 1
transform 1 0 3588 0 1 122944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_222_29
timestamp 1636968456
transform 1 0 3772 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_41
timestamp 1636968456
transform 1 0 4876 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_53
timestamp 1636968456
transform 1 0 5980 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_222_65
timestamp 1
transform 1 0 7084 0 1 122944
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_222_1122
timestamp 1636968456
transform 1 0 104328 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_1134
timestamp 1636968456
transform 1 0 105432 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_222_1146
timestamp 1
transform 1 0 106536 0 1 122944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_222_1148
timestamp 1636968456
transform 1 0 106720 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_222_1160
timestamp 1
transform 1 0 107824 0 1 122944
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_223_3
timestamp 1636968456
transform 1 0 1380 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_15
timestamp 1636968456
transform 1 0 2484 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_27
timestamp 1636968456
transform 1 0 3588 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_39
timestamp 1636968456
transform 1 0 4692 0 -1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_223_51
timestamp 1
transform 1 0 5796 0 -1 124032
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_223_55
timestamp 1
transform 1 0 6164 0 -1 124032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_223_57
timestamp 1636968456
transform 1 0 6348 0 -1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_223_69
timestamp 1
transform 1 0 7452 0 -1 124032
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_223_1122
timestamp 1636968456
transform 1 0 104328 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_1134
timestamp 1636968456
transform 1 0 105432 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_1146
timestamp 1636968456
transform 1 0 106536 0 -1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_223_1158
timestamp 1
transform 1 0 107640 0 -1 124032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_223_1166
timestamp 1
transform 1 0 108376 0 -1 124032
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_224_3
timestamp 1636968456
transform 1 0 1380 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_15
timestamp 1636968456
transform 1 0 2484 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_224_27
timestamp 1
transform 1 0 3588 0 1 124032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_224_29
timestamp 1636968456
transform 1 0 3772 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_41
timestamp 1636968456
transform 1 0 4876 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_53
timestamp 1636968456
transform 1 0 5980 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_224_65
timestamp 1
transform 1 0 7084 0 1 124032
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_224_1122
timestamp 1636968456
transform 1 0 104328 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_1134
timestamp 1636968456
transform 1 0 105432 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_224_1146
timestamp 1
transform 1 0 106536 0 1 124032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_224_1148
timestamp 1636968456
transform 1 0 106720 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_224_1160
timestamp 1
transform 1 0 107824 0 1 124032
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_225_3
timestamp 1636968456
transform 1 0 1380 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_15
timestamp 1636968456
transform 1 0 2484 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_27
timestamp 1636968456
transform 1 0 3588 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_39
timestamp 1636968456
transform 1 0 4692 0 -1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_225_51
timestamp 1
transform 1 0 5796 0 -1 125120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_225_55
timestamp 1
transform 1 0 6164 0 -1 125120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_225_57
timestamp 1636968456
transform 1 0 6348 0 -1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_225_69
timestamp 1
transform 1 0 7452 0 -1 125120
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_225_1122
timestamp 1636968456
transform 1 0 104328 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_1134
timestamp 1636968456
transform 1 0 105432 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_1146
timestamp 1636968456
transform 1 0 106536 0 -1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_225_1158
timestamp 1
transform 1 0 107640 0 -1 125120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_225_1166
timestamp 1
transform 1 0 108376 0 -1 125120
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_226_3
timestamp 1636968456
transform 1 0 1380 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_15
timestamp 1636968456
transform 1 0 2484 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_226_27
timestamp 1
transform 1 0 3588 0 1 125120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_226_29
timestamp 1636968456
transform 1 0 3772 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_41
timestamp 1636968456
transform 1 0 4876 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_53
timestamp 1636968456
transform 1 0 5980 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_226_65
timestamp 1
transform 1 0 7084 0 1 125120
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_226_1122
timestamp 1636968456
transform 1 0 104328 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_1134
timestamp 1636968456
transform 1 0 105432 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_226_1146
timestamp 1
transform 1 0 106536 0 1 125120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_226_1148
timestamp 1636968456
transform 1 0 106720 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_226_1160
timestamp 1
transform 1 0 107824 0 1 125120
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_227_3
timestamp 1636968456
transform 1 0 1380 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_15
timestamp 1636968456
transform 1 0 2484 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_27
timestamp 1636968456
transform 1 0 3588 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_39
timestamp 1636968456
transform 1 0 4692 0 -1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_227_51
timestamp 1
transform 1 0 5796 0 -1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_227_55
timestamp 1
transform 1 0 6164 0 -1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_227_57
timestamp 1636968456
transform 1 0 6348 0 -1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_227_69
timestamp 1
transform 1 0 7452 0 -1 126208
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_227_1122
timestamp 1636968456
transform 1 0 104328 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_1134
timestamp 1636968456
transform 1 0 105432 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_1146
timestamp 1636968456
transform 1 0 106536 0 -1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_227_1158
timestamp 1
transform 1 0 107640 0 -1 126208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_227_1166
timestamp 1
transform 1 0 108376 0 -1 126208
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_228_3
timestamp 1636968456
transform 1 0 1380 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_15
timestamp 1636968456
transform 1 0 2484 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_228_27
timestamp 1
transform 1 0 3588 0 1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_228_29
timestamp 1636968456
transform 1 0 3772 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_41
timestamp 1636968456
transform 1 0 4876 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_53
timestamp 1
transform 1 0 5980 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_57
timestamp 1636968456
transform 1 0 6348 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_69
timestamp 1636968456
transform 1 0 7452 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_81
timestamp 1
transform 1 0 8556 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_85
timestamp 1636968456
transform 1 0 8924 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_97
timestamp 1636968456
transform 1 0 10028 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_109
timestamp 1
transform 1 0 11132 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_113
timestamp 1636968456
transform 1 0 11500 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_125
timestamp 1636968456
transform 1 0 12604 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_137
timestamp 1
transform 1 0 13708 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_141
timestamp 1636968456
transform 1 0 14076 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_153
timestamp 1636968456
transform 1 0 15180 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_165
timestamp 1
transform 1 0 16284 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_169
timestamp 1636968456
transform 1 0 16652 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_181
timestamp 1636968456
transform 1 0 17756 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_193
timestamp 1
transform 1 0 18860 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_197
timestamp 1636968456
transform 1 0 19228 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_209
timestamp 1636968456
transform 1 0 20332 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_221
timestamp 1
transform 1 0 21436 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_225
timestamp 1636968456
transform 1 0 21804 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_237
timestamp 1636968456
transform 1 0 22908 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_249
timestamp 1
transform 1 0 24012 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_253
timestamp 1636968456
transform 1 0 24380 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_265
timestamp 1636968456
transform 1 0 25484 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_277
timestamp 1
transform 1 0 26588 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_281
timestamp 1636968456
transform 1 0 26956 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_293
timestamp 1636968456
transform 1 0 28060 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_305
timestamp 1
transform 1 0 29164 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_309
timestamp 1636968456
transform 1 0 29532 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_321
timestamp 1636968456
transform 1 0 30636 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_333
timestamp 1
transform 1 0 31740 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_337
timestamp 1636968456
transform 1 0 32108 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_349
timestamp 1636968456
transform 1 0 33212 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_361
timestamp 1
transform 1 0 34316 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_365
timestamp 1636968456
transform 1 0 34684 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_228_377
timestamp 1
transform 1 0 35788 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_228_385
timestamp 1
transform 1 0 36524 0 1 126208
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_228_391
timestamp 1
transform 1 0 37076 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_228_393
timestamp 1
transform 1 0 37260 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_402
timestamp 1636968456
transform 1 0 38088 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_228_414
timestamp 1
transform 1 0 39192 0 1 126208
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_228_421
timestamp 1
transform 1 0 39836 0 1 126208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_228_429
timestamp 1
transform 1 0 40572 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_228_444
timestamp 1
transform 1 0 41952 0 1 126208
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_228_449
timestamp 1636968456
transform 1 0 42412 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_461
timestamp 1636968456
transform 1 0 43516 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_473
timestamp 1
transform 1 0 44620 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_483
timestamp 1636968456
transform 1 0 45540 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_228_495
timestamp 1
transform 1 0 46644 0 1 126208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_228_503
timestamp 1
transform 1 0 47380 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_228_505
timestamp 1
transform 1 0 47564 0 1 126208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_228_519
timestamp 1
transform 1 0 48852 0 1 126208
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_228_525
timestamp 1
transform 1 0 49404 0 1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_228_533
timestamp 1636968456
transform 1 0 50140 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_545
timestamp 1636968456
transform 1 0 51244 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_557
timestamp 1
transform 1 0 52348 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_561
timestamp 1636968456
transform 1 0 52716 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_573
timestamp 1636968456
transform 1 0 53820 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_585
timestamp 1
transform 1 0 54924 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_589
timestamp 1636968456
transform 1 0 55292 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_601
timestamp 1636968456
transform 1 0 56396 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_613
timestamp 1
transform 1 0 57500 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_228_617
timestamp 1
transform 1 0 57868 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_228_621
timestamp 1
transform 1 0 58236 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_228_628
timestamp 1
transform 1 0 58880 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_228_638
timestamp 1
transform 1 0 59800 0 1 126208
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_228_645
timestamp 1636968456
transform 1 0 60444 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_228_657
timestamp 1
transform 1 0 61548 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_228_665
timestamp 1
transform 1 0 62284 0 1 126208
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_228_671
timestamp 1
transform 1 0 62836 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_228_673
timestamp 1
transform 1 0 63020 0 1 126208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_228_681
timestamp 1
transform 1 0 63756 0 1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_228_688
timestamp 1636968456
transform 1 0 64400 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_228_707
timestamp 1
transform 1 0 66148 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_228_711
timestamp 1
transform 1 0 66516 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_228_718
timestamp 1
transform 1 0 67160 0 1 126208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_228_726
timestamp 1
transform 1 0 67896 0 1 126208
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_228_729
timestamp 1636968456
transform 1 0 68172 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_228_741
timestamp 1
transform 1 0 69276 0 1 126208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_228_749
timestamp 1
transform 1 0 70012 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_228_755
timestamp 1
transform 1 0 70564 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_228_759
timestamp 1
transform 1 0 70932 0 1 126208
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_228_769
timestamp 1636968456
transform 1 0 71852 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_781
timestamp 1
transform 1 0 72956 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_785
timestamp 1636968456
transform 1 0 73324 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_797
timestamp 1636968456
transform 1 0 74428 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_809
timestamp 1
transform 1 0 75532 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_813
timestamp 1636968456
transform 1 0 75900 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_228_825
timestamp 1
transform 1 0 77004 0 1 126208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_228_833
timestamp 1
transform 1 0 77740 0 1 126208
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_228_839
timestamp 1
transform 1 0 78292 0 1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_228_841
timestamp 1636968456
transform 1 0 78476 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_853
timestamp 1636968456
transform 1 0 79580 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_865
timestamp 1
transform 1 0 80684 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_869
timestamp 1636968456
transform 1 0 81052 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_881
timestamp 1636968456
transform 1 0 82156 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_893
timestamp 1
transform 1 0 83260 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_897
timestamp 1636968456
transform 1 0 83628 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_909
timestamp 1636968456
transform 1 0 84732 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_921
timestamp 1
transform 1 0 85836 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_228_927
timestamp 1
transform 1 0 86388 0 1 126208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_228_935
timestamp 1
transform 1 0 87124 0 1 126208
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_228_939
timestamp 1636968456
transform 1 0 87492 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_228_951
timestamp 1
transform 1 0 88596 0 1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_228_953
timestamp 1636968456
transform 1 0 88780 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_965
timestamp 1636968456
transform 1 0 89884 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_977
timestamp 1
transform 1 0 90988 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_981
timestamp 1636968456
transform 1 0 91356 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_993
timestamp 1636968456
transform 1 0 92460 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_1005
timestamp 1
transform 1 0 93564 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1009
timestamp 1636968456
transform 1 0 93932 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_228_1021
timestamp 1
transform 1 0 95036 0 1 126208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_228_1029
timestamp 1
transform 1 0 95772 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_228_1032
timestamp 1
transform 1 0 96048 0 1 126208
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1037
timestamp 1636968456
transform 1 0 96508 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1049
timestamp 1636968456
transform 1 0 97612 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_1061
timestamp 1
transform 1 0 98716 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1065
timestamp 1636968456
transform 1 0 99084 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1077
timestamp 1636968456
transform 1 0 100188 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_1089
timestamp 1
transform 1 0 101292 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1093
timestamp 1636968456
transform 1 0 101660 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1105
timestamp 1636968456
transform 1 0 102764 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_1117
timestamp 1
transform 1 0 103868 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1121
timestamp 1636968456
transform 1 0 104236 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1133
timestamp 1636968456
transform 1 0 105340 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_228_1145
timestamp 1
transform 1 0 106444 0 1 126208
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1149
timestamp 1636968456
transform 1 0 106812 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_228_1161
timestamp 1
transform 1 0 107916 0 1 126208
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_228_1167
timestamp 1
transform 1 0 108468 0 1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_229_3
timestamp 1636968456
transform 1 0 1380 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_15
timestamp 1636968456
transform 1 0 2484 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_229_27
timestamp 1
transform 1 0 3588 0 -1 127296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_229_29
timestamp 1636968456
transform 1 0 3772 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_41
timestamp 1636968456
transform 1 0 4876 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_53
timestamp 1
transform 1 0 5980 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_57
timestamp 1636968456
transform 1 0 6348 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_69
timestamp 1636968456
transform 1 0 7452 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_81
timestamp 1
transform 1 0 8556 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_85
timestamp 1636968456
transform 1 0 8924 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_97
timestamp 1636968456
transform 1 0 10028 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_109
timestamp 1
transform 1 0 11132 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_113
timestamp 1636968456
transform 1 0 11500 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_125
timestamp 1636968456
transform 1 0 12604 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_137
timestamp 1
transform 1 0 13708 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_141
timestamp 1636968456
transform 1 0 14076 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_153
timestamp 1636968456
transform 1 0 15180 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_165
timestamp 1
transform 1 0 16284 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_169
timestamp 1636968456
transform 1 0 16652 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_181
timestamp 1636968456
transform 1 0 17756 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_193
timestamp 1
transform 1 0 18860 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_197
timestamp 1636968456
transform 1 0 19228 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_209
timestamp 1636968456
transform 1 0 20332 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_221
timestamp 1
transform 1 0 21436 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_225
timestamp 1636968456
transform 1 0 21804 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_237
timestamp 1636968456
transform 1 0 22908 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_249
timestamp 1
transform 1 0 24012 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_253
timestamp 1636968456
transform 1 0 24380 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_265
timestamp 1636968456
transform 1 0 25484 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_277
timestamp 1
transform 1 0 26588 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_281
timestamp 1636968456
transform 1 0 26956 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_293
timestamp 1636968456
transform 1 0 28060 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_305
timestamp 1
transform 1 0 29164 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_309
timestamp 1636968456
transform 1 0 29532 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_321
timestamp 1636968456
transform 1 0 30636 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_333
timestamp 1
transform 1 0 31740 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_337
timestamp 1636968456
transform 1 0 32108 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_349
timestamp 1636968456
transform 1 0 33212 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_361
timestamp 1
transform 1 0 34316 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_365
timestamp 1636968456
transform 1 0 34684 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_377
timestamp 1636968456
transform 1 0 35788 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_389
timestamp 1
transform 1 0 36892 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_393
timestamp 1636968456
transform 1 0 37260 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_405
timestamp 1636968456
transform 1 0 38364 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_417
timestamp 1
transform 1 0 39468 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_421
timestamp 1636968456
transform 1 0 39836 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_433
timestamp 1636968456
transform 1 0 40940 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_445
timestamp 1
transform 1 0 42044 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_449
timestamp 1636968456
transform 1 0 42412 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_461
timestamp 1636968456
transform 1 0 43516 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_473
timestamp 1
transform 1 0 44620 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_477
timestamp 1636968456
transform 1 0 44988 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_489
timestamp 1636968456
transform 1 0 46092 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_501
timestamp 1
transform 1 0 47196 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_505
timestamp 1636968456
transform 1 0 47564 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_517
timestamp 1636968456
transform 1 0 48668 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_529
timestamp 1
transform 1 0 49772 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_533
timestamp 1636968456
transform 1 0 50140 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_545
timestamp 1636968456
transform 1 0 51244 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_557
timestamp 1
transform 1 0 52348 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_561
timestamp 1636968456
transform 1 0 52716 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_573
timestamp 1636968456
transform 1 0 53820 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_585
timestamp 1
transform 1 0 54924 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_589
timestamp 1636968456
transform 1 0 55292 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_601
timestamp 1636968456
transform 1 0 56396 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_613
timestamp 1
transform 1 0 57500 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_617
timestamp 1636968456
transform 1 0 57868 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_629
timestamp 1636968456
transform 1 0 58972 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_641
timestamp 1
transform 1 0 60076 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_645
timestamp 1636968456
transform 1 0 60444 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_657
timestamp 1636968456
transform 1 0 61548 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_669
timestamp 1
transform 1 0 62652 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_673
timestamp 1636968456
transform 1 0 63020 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_685
timestamp 1636968456
transform 1 0 64124 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_697
timestamp 1
transform 1 0 65228 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_701
timestamp 1636968456
transform 1 0 65596 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_713
timestamp 1636968456
transform 1 0 66700 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_725
timestamp 1
transform 1 0 67804 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_729
timestamp 1636968456
transform 1 0 68172 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_741
timestamp 1636968456
transform 1 0 69276 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_753
timestamp 1
transform 1 0 70380 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_757
timestamp 1636968456
transform 1 0 70748 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_769
timestamp 1636968456
transform 1 0 71852 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_781
timestamp 1
transform 1 0 72956 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_785
timestamp 1636968456
transform 1 0 73324 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_797
timestamp 1636968456
transform 1 0 74428 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_809
timestamp 1
transform 1 0 75532 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_813
timestamp 1636968456
transform 1 0 75900 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_825
timestamp 1636968456
transform 1 0 77004 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_837
timestamp 1
transform 1 0 78108 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_841
timestamp 1636968456
transform 1 0 78476 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_853
timestamp 1636968456
transform 1 0 79580 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_865
timestamp 1
transform 1 0 80684 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_869
timestamp 1636968456
transform 1 0 81052 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_881
timestamp 1636968456
transform 1 0 82156 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_893
timestamp 1
transform 1 0 83260 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_897
timestamp 1636968456
transform 1 0 83628 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_909
timestamp 1636968456
transform 1 0 84732 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_921
timestamp 1
transform 1 0 85836 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_925
timestamp 1636968456
transform 1 0 86204 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_937
timestamp 1636968456
transform 1 0 87308 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_949
timestamp 1
transform 1 0 88412 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_953
timestamp 1636968456
transform 1 0 88780 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_965
timestamp 1636968456
transform 1 0 89884 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_977
timestamp 1
transform 1 0 90988 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_981
timestamp 1636968456
transform 1 0 91356 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_993
timestamp 1636968456
transform 1 0 92460 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_1005
timestamp 1
transform 1 0 93564 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1009
timestamp 1636968456
transform 1 0 93932 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1021
timestamp 1636968456
transform 1 0 95036 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_1033
timestamp 1
transform 1 0 96140 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1037
timestamp 1636968456
transform 1 0 96508 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1049
timestamp 1636968456
transform 1 0 97612 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_1061
timestamp 1
transform 1 0 98716 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1065
timestamp 1636968456
transform 1 0 99084 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1077
timestamp 1636968456
transform 1 0 100188 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_1089
timestamp 1
transform 1 0 101292 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1093
timestamp 1636968456
transform 1 0 101660 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1105
timestamp 1636968456
transform 1 0 102764 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_1117
timestamp 1
transform 1 0 103868 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1121
timestamp 1636968456
transform 1 0 104236 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1133
timestamp 1636968456
transform 1 0 105340 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_229_1145
timestamp 1
transform 1 0 106444 0 -1 127296
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1149
timestamp 1636968456
transform 1 0 106812 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_229_1161
timestamp 1
transform 1 0 107916 0 -1 127296
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_229_1167
timestamp 1
transform 1 0 108468 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 92644 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 93380 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform 1 0 104420 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1
transform 1 0 1380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1
transform 1 0 1380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1
transform 1 0 1380 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1
transform 1 0 1380 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1
transform 1 0 1380 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1
transform -1 0 2300 0 -1 70720
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1
transform 1 0 1380 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1
transform 1 0 1380 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1
transform 1 0 1380 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1
transform 1 0 1380 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1
transform 1 0 1380 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1
transform 1 0 1380 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1
transform 1 0 1380 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1
transform -1 0 26128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1
transform -1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1
transform -1 0 39008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1
transform -1 0 40296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1
transform -1 0 41584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1
transform 1 0 41952 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1
transform 1 0 43240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1
transform -1 0 27416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1
transform -1 0 28704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1
transform 1 0 29072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1
transform -1 0 31924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1
transform -1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1
transform -1 0 34500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1
transform -1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1
transform 1 0 36156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1
transform 1 0 1380 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1
transform 1 0 1380 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1
transform 1 0 1380 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1
transform 1 0 1380 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1
transform 1 0 1380 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1
transform 1 0 1380 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1
transform 1 0 1380 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1
transform 1 0 1380 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1
transform 1 0 1380 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1
transform 1 0 1380 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1
transform 1 0 1380 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1
transform 1 0 1380 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1
transform 1 0 1380 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1
transform 1 0 1380 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1
transform 1 0 1380 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1
transform 1 0 1380 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1
transform -1 0 108560 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew86
timestamp 1
transform -1 0 105156 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  load_slew87
timestamp 1
transform 1 0 95036 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  load_slew88
timestamp 1
transform 1 0 104328 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  load_slew89
timestamp 1
transform -1 0 104604 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew90
timestamp 1
transform 1 0 104328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  load_slew91
timestamp 1
transform -1 0 104696 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  load_slew92
timestamp 1
transform 1 0 98164 0 1 66368
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  load_slew93
timestamp 1
transform -1 0 96876 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew94
timestamp 1
transform 1 0 104788 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  load_slew95
timestamp 1
transform 1 0 99084 0 -1 66368
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  load_slew96
timestamp 1
transform 1 0 99084 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  load_slew97
timestamp 1
transform 1 0 94944 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew98
timestamp 1
transform 1 0 101660 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  load_slew99
timestamp 1
transform 1 0 101660 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  load_slew100
timestamp 1
transform 1 0 99452 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  load_slew101
timestamp 1
transform -1 0 105248 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  load_slew102
timestamp 1
transform 1 0 96140 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew103
timestamp 1
transform 1 0 99084 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  load_slew104
timestamp 1
transform -1 0 104696 0 1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  load_slew105
timestamp 1
transform -1 0 105524 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  load_slew106
timestamp 1
transform -1 0 91172 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  load_slew107
timestamp 1
transform -1 0 104604 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew108
timestamp 1
transform -1 0 104696 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  load_slew109
timestamp 1
transform -1 0 104972 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  load_slew110
timestamp 1
transform 1 0 94024 0 1 67456
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  load_slew111
timestamp 1
transform -1 0 91632 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mem_i0_115
timestamp 1
transform -1 0 104604 0 1 59840
box -38 -48 314 592
use ram_256x16  mem_i0
timestamp 0
transform 1 0 10000 0 1 10000
box 0 0 1 1
use sky130_fd_sc_hd__conb_1  mem_i1_116
timestamp 1
transform -1 0 104604 0 1 119680
box -38 -48 314 592
use ram_256x16  mem_i1
timestamp 0
transform 1 0 10000 0 1 70000
box 0 0 1 1
use sky130_fd_sc_hd__buf_1  output52
timestamp 1
transform -1 0 1656 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output53
timestamp 1
transform 1 0 108284 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output54
timestamp 1
transform 1 0 108284 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output55
timestamp 1
transform 1 0 108284 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output56
timestamp 1
transform 1 0 108284 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output57
timestamp 1
transform 1 0 108284 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output58
timestamp 1
transform 1 0 108284 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output59
timestamp 1
transform -1 0 1656 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output60
timestamp 1
transform -1 0 1656 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output61
timestamp 1
transform -1 0 1656 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output62
timestamp 1
transform -1 0 1656 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output63
timestamp 1
transform -1 0 1656 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output64
timestamp 1
transform -1 0 1656 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output65
timestamp 1
transform 1 0 108284 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output66
timestamp 1
transform 1 0 108284 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output67
timestamp 1
transform 1 0 108284 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_230
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 108836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_231
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 108836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_232
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 108836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_233
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 108836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_234
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 108836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_235
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 108836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_236
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 108836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_237
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 108836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_238
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 108836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_239
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 108836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_459
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_673
timestamp 1
transform -1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_460
timestamp 1
transform 1 0 104052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_16
timestamp 1
transform -1 0 108836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_240
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_567
timestamp 1
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_461
timestamp 1
transform 1 0 104052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_17
timestamp 1
transform -1 0 108836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_241
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_568
timestamp 1
transform -1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_462
timestamp 1
transform 1 0 104052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_18
timestamp 1
transform -1 0 108836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_242
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_569
timestamp 1
transform -1 0 7912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_463
timestamp 1
transform 1 0 104052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_19
timestamp 1
transform -1 0 108836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Left_243
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Right_570
timestamp 1
transform -1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_464
timestamp 1
transform 1 0 104052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_20
timestamp 1
transform -1 0 108836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Left_244
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Right_571
timestamp 1
transform -1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_465
timestamp 1
transform 1 0 104052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_21
timestamp 1
transform -1 0 108836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Left_245
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Right_572
timestamp 1
transform -1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_466
timestamp 1
transform 1 0 104052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_22
timestamp 1
transform -1 0 108836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Left_246
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Right_573
timestamp 1
transform -1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_467
timestamp 1
transform 1 0 104052 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_23
timestamp 1
transform -1 0 108836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Left_247
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Right_574
timestamp 1
transform -1 0 7912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_468
timestamp 1
transform 1 0 104052 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_24
timestamp 1
transform -1 0 108836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Left_248
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Right_575
timestamp 1
transform -1 0 7912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_469
timestamp 1
transform 1 0 104052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_25
timestamp 1
transform -1 0 108836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Left_249
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Right_576
timestamp 1
transform -1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_470
timestamp 1
transform 1 0 104052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_26
timestamp 1
transform -1 0 108836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Left_250
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Right_577
timestamp 1
transform -1 0 7912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_471
timestamp 1
transform 1 0 104052 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_27
timestamp 1
transform -1 0 108836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Left_251
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Right_578
timestamp 1
transform -1 0 7912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_472
timestamp 1
transform 1 0 104052 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_28
timestamp 1
transform -1 0 108836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Left_252
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Right_579
timestamp 1
transform -1 0 7912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_473
timestamp 1
transform 1 0 104052 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_29
timestamp 1
transform -1 0 108836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Left_253
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Right_580
timestamp 1
transform -1 0 7912 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_474
timestamp 1
transform 1 0 104052 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_30
timestamp 1
transform -1 0 108836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Left_254
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Right_581
timestamp 1
transform -1 0 7912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_475
timestamp 1
transform 1 0 104052 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_31
timestamp 1
transform -1 0 108836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Left_255
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Right_582
timestamp 1
transform -1 0 7912 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_476
timestamp 1
transform 1 0 104052 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_32
timestamp 1
transform -1 0 108836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Left_256
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Right_583
timestamp 1
transform -1 0 7912 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_477
timestamp 1
transform 1 0 104052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_33
timestamp 1
transform -1 0 108836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Left_257
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Right_584
timestamp 1
transform -1 0 7912 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_478
timestamp 1
transform 1 0 104052 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_34
timestamp 1
transform -1 0 108836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Left_258
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Right_585
timestamp 1
transform -1 0 7912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_479
timestamp 1
transform 1 0 104052 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_35
timestamp 1
transform -1 0 108836 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Left_259
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Right_586
timestamp 1
transform -1 0 7912 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_480
timestamp 1
transform 1 0 104052 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_36
timestamp 1
transform -1 0 108836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Left_260
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Right_587
timestamp 1
transform -1 0 7912 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_481
timestamp 1
transform 1 0 104052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_37
timestamp 1
transform -1 0 108836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Left_261
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Right_588
timestamp 1
transform -1 0 7912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_482
timestamp 1
transform 1 0 104052 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_38
timestamp 1
transform -1 0 108836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Left_262
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Right_589
timestamp 1
transform -1 0 7912 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_483
timestamp 1
transform 1 0 104052 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_39
timestamp 1
transform -1 0 108836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Left_263
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Right_590
timestamp 1
transform -1 0 7912 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_484
timestamp 1
transform 1 0 104052 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_40
timestamp 1
transform -1 0 108836 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Left_264
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Right_591
timestamp 1
transform -1 0 7912 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_485
timestamp 1
transform 1 0 104052 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_41
timestamp 1
transform -1 0 108836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Left_265
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Right_592
timestamp 1
transform -1 0 7912 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_486
timestamp 1
transform 1 0 104052 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_42
timestamp 1
transform -1 0 108836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Left_266
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Right_593
timestamp 1
transform -1 0 7912 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_487
timestamp 1
transform 1 0 104052 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_43
timestamp 1
transform -1 0 108836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Left_267
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Right_594
timestamp 1
transform -1 0 7912 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_488
timestamp 1
transform 1 0 104052 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_44
timestamp 1
transform -1 0 108836 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Left_268
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Right_595
timestamp 1
transform -1 0 7912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_489
timestamp 1
transform 1 0 104052 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_45
timestamp 1
transform -1 0 108836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Left_269
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Right_596
timestamp 1
transform -1 0 7912 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_490
timestamp 1
transform 1 0 104052 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_46
timestamp 1
transform -1 0 108836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Left_270
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Right_597
timestamp 1
transform -1 0 7912 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_491
timestamp 1
transform 1 0 104052 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_47
timestamp 1
transform -1 0 108836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Left_271
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Right_598
timestamp 1
transform -1 0 7912 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_492
timestamp 1
transform 1 0 104052 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_48
timestamp 1
transform -1 0 108836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Left_272
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Right_599
timestamp 1
transform -1 0 7912 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_493
timestamp 1
transform 1 0 104052 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_49
timestamp 1
transform -1 0 108836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Left_273
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Right_600
timestamp 1
transform -1 0 7912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_494
timestamp 1
transform 1 0 104052 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_50
timestamp 1
transform -1 0 108836 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Left_274
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Right_601
timestamp 1
transform -1 0 7912 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_495
timestamp 1
transform 1 0 104052 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_51
timestamp 1
transform -1 0 108836 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Left_275
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Right_602
timestamp 1
transform -1 0 7912 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_496
timestamp 1
transform 1 0 104052 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_52
timestamp 1
transform -1 0 108836 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Left_276
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Right_603
timestamp 1
transform -1 0 7912 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_497
timestamp 1
transform 1 0 104052 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_53
timestamp 1
transform -1 0 108836 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Left_277
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Right_604
timestamp 1
transform -1 0 7912 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_498
timestamp 1
transform 1 0 104052 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_54
timestamp 1
transform -1 0 108836 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Left_278
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Right_605
timestamp 1
transform -1 0 7912 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_499
timestamp 1
transform 1 0 104052 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_55
timestamp 1
transform -1 0 108836 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Left_279
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Right_606
timestamp 1
transform -1 0 7912 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_500
timestamp 1
transform 1 0 104052 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_56
timestamp 1
transform -1 0 108836 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Left_280
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Right_607
timestamp 1
transform -1 0 7912 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_501
timestamp 1
transform 1 0 104052 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_57
timestamp 1
transform -1 0 108836 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Left_281
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Right_608
timestamp 1
transform -1 0 7912 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_502
timestamp 1
transform 1 0 104052 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_58
timestamp 1
transform -1 0 108836 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Left_282
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Right_609
timestamp 1
transform -1 0 7912 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_503
timestamp 1
transform 1 0 104052 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_59
timestamp 1
transform -1 0 108836 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Left_283
timestamp 1
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Right_610
timestamp 1
transform -1 0 7912 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_504
timestamp 1
transform 1 0 104052 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_60
timestamp 1
transform -1 0 108836 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Left_284
timestamp 1
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Right_611
timestamp 1
transform -1 0 7912 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_505
timestamp 1
transform 1 0 104052 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_61
timestamp 1
transform -1 0 108836 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Left_285
timestamp 1
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Right_612
timestamp 1
transform -1 0 7912 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_506
timestamp 1
transform 1 0 104052 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_62
timestamp 1
transform -1 0 108836 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Left_286
timestamp 1
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Right_613
timestamp 1
transform -1 0 7912 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_507
timestamp 1
transform 1 0 104052 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_63
timestamp 1
transform -1 0 108836 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Left_287
timestamp 1
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Right_614
timestamp 1
transform -1 0 7912 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_508
timestamp 1
transform 1 0 104052 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_64
timestamp 1
transform -1 0 108836 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Left_288
timestamp 1
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Right_615
timestamp 1
transform -1 0 7912 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_509
timestamp 1
transform 1 0 104052 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_65
timestamp 1
transform -1 0 108836 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Left_289
timestamp 1
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Right_616
timestamp 1
transform -1 0 7912 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_510
timestamp 1
transform 1 0 104052 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_66
timestamp 1
transform -1 0 108836 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Left_290
timestamp 1
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Right_617
timestamp 1
transform -1 0 7912 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_511
timestamp 1
transform 1 0 104052 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_67
timestamp 1
transform -1 0 108836 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Left_291
timestamp 1
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Right_618
timestamp 1
transform -1 0 7912 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_512
timestamp 1
transform 1 0 104052 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_68
timestamp 1
transform -1 0 108836 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Left_292
timestamp 1
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Right_619
timestamp 1
transform -1 0 7912 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_513
timestamp 1
transform 1 0 104052 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_69
timestamp 1
transform -1 0 108836 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Left_293
timestamp 1
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Right_620
timestamp 1
transform -1 0 7912 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_514
timestamp 1
transform 1 0 104052 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_70
timestamp 1
transform -1 0 108836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Left_294
timestamp 1
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Right_621
timestamp 1
transform -1 0 7912 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_515
timestamp 1
transform 1 0 104052 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_71
timestamp 1
transform -1 0 108836 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Left_295
timestamp 1
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Right_622
timestamp 1
transform -1 0 7912 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_516
timestamp 1
transform 1 0 104052 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_72
timestamp 1
transform -1 0 108836 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Left_296
timestamp 1
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Right_623
timestamp 1
transform -1 0 7912 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Left_517
timestamp 1
transform 1 0 104052 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Right_73
timestamp 1
transform -1 0 108836 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Left_297
timestamp 1
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Right_624
timestamp 1
transform -1 0 7912 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Left_518
timestamp 1
transform 1 0 104052 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Right_74
timestamp 1
transform -1 0 108836 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Left_298
timestamp 1
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Right_625
timestamp 1
transform -1 0 7912 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Left_519
timestamp 1
transform 1 0 104052 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Right_75
timestamp 1
transform -1 0 108836 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Left_299
timestamp 1
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Right_626
timestamp 1
transform -1 0 7912 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Left_520
timestamp 1
transform 1 0 104052 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Right_76
timestamp 1
transform -1 0 108836 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Left_300
timestamp 1
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Right_627
timestamp 1
transform -1 0 7912 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Left_521
timestamp 1
transform 1 0 104052 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Right_77
timestamp 1
transform -1 0 108836 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Left_301
timestamp 1
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Right_628
timestamp 1
transform -1 0 7912 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Left_522
timestamp 1
transform 1 0 104052 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Right_78
timestamp 1
transform -1 0 108836 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Left_302
timestamp 1
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Right_629
timestamp 1
transform -1 0 7912 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Left_523
timestamp 1
transform 1 0 104052 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Right_79
timestamp 1
transform -1 0 108836 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Left_303
timestamp 1
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Right_630
timestamp 1
transform -1 0 7912 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Left_524
timestamp 1
transform 1 0 104052 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Right_80
timestamp 1
transform -1 0 108836 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Left_304
timestamp 1
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Right_631
timestamp 1
transform -1 0 7912 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Left_525
timestamp 1
transform 1 0 104052 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Right_81
timestamp 1
transform -1 0 108836 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Left_305
timestamp 1
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Right_632
timestamp 1
transform -1 0 7912 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Left_526
timestamp 1
transform 1 0 104052 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Right_82
timestamp 1
transform -1 0 108836 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Left_306
timestamp 1
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Right_633
timestamp 1
transform -1 0 7912 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Left_527
timestamp 1
transform 1 0 104052 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Right_83
timestamp 1
transform -1 0 108836 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Left_307
timestamp 1
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Right_634
timestamp 1
transform -1 0 7912 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Left_528
timestamp 1
transform 1 0 104052 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Right_84
timestamp 1
transform -1 0 108836 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Left_308
timestamp 1
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Right_635
timestamp 1
transform -1 0 7912 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Left_529
timestamp 1
transform 1 0 104052 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Right_85
timestamp 1
transform -1 0 108836 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Left_309
timestamp 1
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Right_636
timestamp 1
transform -1 0 7912 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Left_530
timestamp 1
transform 1 0 104052 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Right_86
timestamp 1
transform -1 0 108836 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Left_310
timestamp 1
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Right_637
timestamp 1
transform -1 0 7912 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Left_531
timestamp 1
transform 1 0 104052 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Right_87
timestamp 1
transform -1 0 108836 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Left_311
timestamp 1
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Right_638
timestamp 1
transform -1 0 7912 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Left_532
timestamp 1
transform 1 0 104052 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Right_88
timestamp 1
transform -1 0 108836 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Left_312
timestamp 1
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Right_639
timestamp 1
transform -1 0 7912 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Left_533
timestamp 1
transform 1 0 104052 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Right_89
timestamp 1
transform -1 0 108836 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Left_313
timestamp 1
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Right_640
timestamp 1
transform -1 0 7912 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Left_534
timestamp 1
transform 1 0 104052 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Right_90
timestamp 1
transform -1 0 108836 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Left_314
timestamp 1
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Right_641
timestamp 1
transform -1 0 7912 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Left_535
timestamp 1
transform 1 0 104052 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Right_91
timestamp 1
transform -1 0 108836 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Left_315
timestamp 1
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Right_642
timestamp 1
transform -1 0 7912 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Left_536
timestamp 1
transform 1 0 104052 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Right_92
timestamp 1
transform -1 0 108836 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Left_316
timestamp 1
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Right_643
timestamp 1
transform -1 0 7912 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Left_537
timestamp 1
transform 1 0 104052 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Right_93
timestamp 1
transform -1 0 108836 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Left_317
timestamp 1
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Right_644
timestamp 1
transform -1 0 7912 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Left_538
timestamp 1
transform 1 0 104052 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Right_94
timestamp 1
transform -1 0 108836 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Left_318
timestamp 1
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Right_645
timestamp 1
transform -1 0 7912 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Left_539
timestamp 1
transform 1 0 104052 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Right_95
timestamp 1
transform -1 0 108836 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Left_319
timestamp 1
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Right_646
timestamp 1
transform -1 0 7912 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Left_540
timestamp 1
transform 1 0 104052 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Right_96
timestamp 1
transform -1 0 108836 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Left_320
timestamp 1
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Right_647
timestamp 1
transform -1 0 7912 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Left_541
timestamp 1
transform 1 0 104052 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Right_97
timestamp 1
transform -1 0 108836 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Left_321
timestamp 1
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Right_648
timestamp 1
transform -1 0 7912 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Left_542
timestamp 1
transform 1 0 104052 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Right_98
timestamp 1
transform -1 0 108836 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Left_322
timestamp 1
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Right_649
timestamp 1
transform -1 0 7912 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Left_543
timestamp 1
transform 1 0 104052 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Right_99
timestamp 1
transform -1 0 108836 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Left_323
timestamp 1
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Right_650
timestamp 1
transform -1 0 7912 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Left_544
timestamp 1
transform 1 0 104052 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Right_100
timestamp 1
transform -1 0 108836 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Left_324
timestamp 1
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Right_651
timestamp 1
transform -1 0 7912 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Left_545
timestamp 1
transform 1 0 104052 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Right_101
timestamp 1
transform -1 0 108836 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Left_325
timestamp 1
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Right_652
timestamp 1
transform -1 0 7912 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Left_546
timestamp 1
transform 1 0 104052 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Right_102
timestamp 1
transform -1 0 108836 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Left_326
timestamp 1
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Right_653
timestamp 1
transform -1 0 7912 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Left_547
timestamp 1
transform 1 0 104052 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Right_103
timestamp 1
transform -1 0 108836 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Left_327
timestamp 1
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Right_654
timestamp 1
transform -1 0 7912 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Left_548
timestamp 1
transform 1 0 104052 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Right_104
timestamp 1
transform -1 0 108836 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Left_328
timestamp 1
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Right_655
timestamp 1
transform -1 0 7912 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Left_549
timestamp 1
transform 1 0 104052 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Right_105
timestamp 1
transform -1 0 108836 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Left_329
timestamp 1
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Right_656
timestamp 1
transform -1 0 7912 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Left_550
timestamp 1
transform 1 0 104052 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Right_106
timestamp 1
transform -1 0 108836 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Left_330
timestamp 1
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Right_657
timestamp 1
transform -1 0 7912 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Left_551
timestamp 1
transform 1 0 104052 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Right_107
timestamp 1
transform -1 0 108836 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Left_331
timestamp 1
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Right_658
timestamp 1
transform -1 0 7912 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Left_552
timestamp 1
transform 1 0 104052 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Right_108
timestamp 1
transform -1 0 108836 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Left_332
timestamp 1
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Right_659
timestamp 1
transform -1 0 7912 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Left_553
timestamp 1
transform 1 0 104052 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Right_109
timestamp 1
transform -1 0 108836 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Left_333
timestamp 1
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Right_660
timestamp 1
transform -1 0 7912 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Left_554
timestamp 1
transform 1 0 104052 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Right_110
timestamp 1
transform -1 0 108836 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Left_334
timestamp 1
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Right_661
timestamp 1
transform -1 0 7912 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Left_555
timestamp 1
transform 1 0 104052 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Right_111
timestamp 1
transform -1 0 108836 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Left_335
timestamp 1
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Right_662
timestamp 1
transform -1 0 7912 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Left_556
timestamp 1
transform 1 0 104052 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Right_112
timestamp 1
transform -1 0 108836 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Left_336
timestamp 1
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Right_663
timestamp 1
transform -1 0 7912 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Left_557
timestamp 1
transform 1 0 104052 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Right_113
timestamp 1
transform -1 0 108836 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Left_337
timestamp 1
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Right_664
timestamp 1
transform -1 0 7912 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Left_558
timestamp 1
transform 1 0 104052 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Right_114
timestamp 1
transform -1 0 108836 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Left_338
timestamp 1
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Right_665
timestamp 1
transform -1 0 7912 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Left_559
timestamp 1
transform 1 0 104052 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Right_115
timestamp 1
transform -1 0 108836 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Left_339
timestamp 1
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Right_666
timestamp 1
transform -1 0 7912 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Left_560
timestamp 1
transform 1 0 104052 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Right_116
timestamp 1
transform -1 0 108836 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Left_340
timestamp 1
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Right_667
timestamp 1
transform -1 0 7912 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Left_561
timestamp 1
transform 1 0 104052 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Right_117
timestamp 1
transform -1 0 108836 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Left_341
timestamp 1
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Right_668
timestamp 1
transform -1 0 7912 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Left_562
timestamp 1
transform 1 0 104052 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Right_118
timestamp 1
transform -1 0 108836 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Left_342
timestamp 1
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Right_669
timestamp 1
transform -1 0 7912 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Left_563
timestamp 1
transform 1 0 104052 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Right_119
timestamp 1
transform -1 0 108836 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Left_343
timestamp 1
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Right_670
timestamp 1
transform -1 0 7912 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Left_564
timestamp 1
transform 1 0 104052 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Right_120
timestamp 1
transform -1 0 108836 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Left_344
timestamp 1
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Right_671
timestamp 1
transform -1 0 7912 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Left_565
timestamp 1
transform 1 0 104052 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Right_121
timestamp 1
transform -1 0 108836 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Left_345
timestamp 1
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Right_672
timestamp 1
transform -1 0 7912 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Left_566
timestamp 1
transform 1 0 104052 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Right_122
timestamp 1
transform -1 0 108836 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Left_347
timestamp 1
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Right_10
timestamp 1
transform -1 0 108836 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Left_348
timestamp 1
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Right_11
timestamp 1
transform -1 0 108836 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Left_349
timestamp 1
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Right_12
timestamp 1
transform -1 0 108836 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Left_350
timestamp 1
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Right_13
timestamp 1
transform -1 0 108836 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Left_346
timestamp 1
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Right_781
timestamp 1
transform -1 0 7912 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Left_674
timestamp 1
transform 1 0 104052 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Right_123
timestamp 1
transform -1 0 108836 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Left_351
timestamp 1
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Right_782
timestamp 1
transform -1 0 7912 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Left_675
timestamp 1
transform 1 0 104052 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Right_124
timestamp 1
transform -1 0 108836 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Left_352
timestamp 1
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Right_783
timestamp 1
transform -1 0 7912 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Left_676
timestamp 1
transform 1 0 104052 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Right_125
timestamp 1
transform -1 0 108836 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Left_353
timestamp 1
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Right_784
timestamp 1
transform -1 0 7912 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Left_677
timestamp 1
transform 1 0 104052 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Right_126
timestamp 1
transform -1 0 108836 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Left_354
timestamp 1
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Right_785
timestamp 1
transform -1 0 7912 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Left_678
timestamp 1
transform 1 0 104052 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Right_127
timestamp 1
transform -1 0 108836 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Left_355
timestamp 1
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Right_786
timestamp 1
transform -1 0 7912 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Left_679
timestamp 1
transform 1 0 104052 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Right_128
timestamp 1
transform -1 0 108836 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Left_356
timestamp 1
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Right_787
timestamp 1
transform -1 0 7912 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Left_680
timestamp 1
transform 1 0 104052 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Right_129
timestamp 1
transform -1 0 108836 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Left_357
timestamp 1
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Right_788
timestamp 1
transform -1 0 7912 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Left_681
timestamp 1
transform 1 0 104052 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Right_130
timestamp 1
transform -1 0 108836 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Left_358
timestamp 1
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Right_789
timestamp 1
transform -1 0 7912 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Left_682
timestamp 1
transform 1 0 104052 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Right_131
timestamp 1
transform -1 0 108836 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Left_359
timestamp 1
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Right_790
timestamp 1
transform -1 0 7912 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Left_683
timestamp 1
transform 1 0 104052 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Right_132
timestamp 1
transform -1 0 108836 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Left_360
timestamp 1
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Right_791
timestamp 1
transform -1 0 7912 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Left_684
timestamp 1
transform 1 0 104052 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Right_133
timestamp 1
transform -1 0 108836 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Left_361
timestamp 1
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Right_792
timestamp 1
transform -1 0 7912 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Left_685
timestamp 1
transform 1 0 104052 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Right_134
timestamp 1
transform -1 0 108836 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Left_362
timestamp 1
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Right_793
timestamp 1
transform -1 0 7912 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Left_686
timestamp 1
transform 1 0 104052 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Right_135
timestamp 1
transform -1 0 108836 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Left_363
timestamp 1
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Right_794
timestamp 1
transform -1 0 7912 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Left_687
timestamp 1
transform 1 0 104052 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Right_136
timestamp 1
transform -1 0 108836 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Left_364
timestamp 1
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Right_795
timestamp 1
transform -1 0 7912 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Left_688
timestamp 1
transform 1 0 104052 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Right_137
timestamp 1
transform -1 0 108836 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Left_365
timestamp 1
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Right_796
timestamp 1
transform -1 0 7912 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Left_689
timestamp 1
transform 1 0 104052 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Right_138
timestamp 1
transform -1 0 108836 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Left_366
timestamp 1
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Right_797
timestamp 1
transform -1 0 7912 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Left_690
timestamp 1
transform 1 0 104052 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Right_139
timestamp 1
transform -1 0 108836 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Left_367
timestamp 1
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Right_798
timestamp 1
transform -1 0 7912 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Left_691
timestamp 1
transform 1 0 104052 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Right_140
timestamp 1
transform -1 0 108836 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Left_368
timestamp 1
transform 1 0 1104 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Right_799
timestamp 1
transform -1 0 7912 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Left_692
timestamp 1
transform 1 0 104052 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Right_141
timestamp 1
transform -1 0 108836 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Left_369
timestamp 1
transform 1 0 1104 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Right_800
timestamp 1
transform -1 0 7912 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Left_693
timestamp 1
transform 1 0 104052 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Right_142
timestamp 1
transform -1 0 108836 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Left_370
timestamp 1
transform 1 0 1104 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Right_801
timestamp 1
transform -1 0 7912 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Left_694
timestamp 1
transform 1 0 104052 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Right_143
timestamp 1
transform -1 0 108836 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Left_371
timestamp 1
transform 1 0 1104 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Right_802
timestamp 1
transform -1 0 7912 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Left_695
timestamp 1
transform 1 0 104052 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Right_144
timestamp 1
transform -1 0 108836 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Left_372
timestamp 1
transform 1 0 1104 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Right_803
timestamp 1
transform -1 0 7912 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Left_696
timestamp 1
transform 1 0 104052 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Right_145
timestamp 1
transform -1 0 108836 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Left_373
timestamp 1
transform 1 0 1104 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Right_804
timestamp 1
transform -1 0 7912 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Left_697
timestamp 1
transform 1 0 104052 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Right_146
timestamp 1
transform -1 0 108836 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Left_374
timestamp 1
transform 1 0 1104 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Right_805
timestamp 1
transform -1 0 7912 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Left_698
timestamp 1
transform 1 0 104052 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Right_147
timestamp 1
transform -1 0 108836 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Left_375
timestamp 1
transform 1 0 1104 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Right_806
timestamp 1
transform -1 0 7912 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Left_699
timestamp 1
transform 1 0 104052 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Right_148
timestamp 1
transform -1 0 108836 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Left_376
timestamp 1
transform 1 0 1104 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Right_807
timestamp 1
transform -1 0 7912 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Left_700
timestamp 1
transform 1 0 104052 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Right_149
timestamp 1
transform -1 0 108836 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Left_377
timestamp 1
transform 1 0 1104 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Right_808
timestamp 1
transform -1 0 7912 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Left_701
timestamp 1
transform 1 0 104052 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Right_150
timestamp 1
transform -1 0 108836 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Left_378
timestamp 1
transform 1 0 1104 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Right_809
timestamp 1
transform -1 0 7912 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Left_702
timestamp 1
transform 1 0 104052 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Right_151
timestamp 1
transform -1 0 108836 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Left_379
timestamp 1
transform 1 0 1104 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Right_810
timestamp 1
transform -1 0 7912 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Left_703
timestamp 1
transform 1 0 104052 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Right_152
timestamp 1
transform -1 0 108836 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Left_380
timestamp 1
transform 1 0 1104 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Right_811
timestamp 1
transform -1 0 7912 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Left_704
timestamp 1
transform 1 0 104052 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Right_153
timestamp 1
transform -1 0 108836 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Left_381
timestamp 1
transform 1 0 1104 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Right_812
timestamp 1
transform -1 0 7912 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Left_705
timestamp 1
transform 1 0 104052 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Right_154
timestamp 1
transform -1 0 108836 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Left_382
timestamp 1
transform 1 0 1104 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Right_813
timestamp 1
transform -1 0 7912 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Left_706
timestamp 1
transform 1 0 104052 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Right_155
timestamp 1
transform -1 0 108836 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Left_383
timestamp 1
transform 1 0 1104 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Right_814
timestamp 1
transform -1 0 7912 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Left_707
timestamp 1
transform 1 0 104052 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Right_156
timestamp 1
transform -1 0 108836 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Left_384
timestamp 1
transform 1 0 1104 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Right_815
timestamp 1
transform -1 0 7912 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Left_708
timestamp 1
transform 1 0 104052 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Right_157
timestamp 1
transform -1 0 108836 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Left_385
timestamp 1
transform 1 0 1104 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Right_816
timestamp 1
transform -1 0 7912 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_2_Left_709
timestamp 1
transform 1 0 104052 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_2_Right_158
timestamp 1
transform -1 0 108836 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Left_386
timestamp 1
transform 1 0 1104 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Right_817
timestamp 1
transform -1 0 7912 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_2_Left_710
timestamp 1
transform 1 0 104052 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_2_Right_159
timestamp 1
transform -1 0 108836 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Left_387
timestamp 1
transform 1 0 1104 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Right_818
timestamp 1
transform -1 0 7912 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_2_Left_711
timestamp 1
transform 1 0 104052 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_2_Right_160
timestamp 1
transform -1 0 108836 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Left_388
timestamp 1
transform 1 0 1104 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Right_819
timestamp 1
transform -1 0 7912 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_2_Left_712
timestamp 1
transform 1 0 104052 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_2_Right_161
timestamp 1
transform -1 0 108836 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Left_389
timestamp 1
transform 1 0 1104 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Right_820
timestamp 1
transform -1 0 7912 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_2_Left_713
timestamp 1
transform 1 0 104052 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_2_Right_162
timestamp 1
transform -1 0 108836 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Left_390
timestamp 1
transform 1 0 1104 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Right_821
timestamp 1
transform -1 0 7912 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_2_Left_714
timestamp 1
transform 1 0 104052 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_2_Right_163
timestamp 1
transform -1 0 108836 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Left_391
timestamp 1
transform 1 0 1104 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Right_822
timestamp 1
transform -1 0 7912 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_2_Left_715
timestamp 1
transform 1 0 104052 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_2_Right_164
timestamp 1
transform -1 0 108836 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Left_392
timestamp 1
transform 1 0 1104 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Right_823
timestamp 1
transform -1 0 7912 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_2_Left_716
timestamp 1
transform 1 0 104052 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_2_Right_165
timestamp 1
transform -1 0 108836 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_1_Left_393
timestamp 1
transform 1 0 1104 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_1_Right_824
timestamp 1
transform -1 0 7912 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_2_Left_717
timestamp 1
transform 1 0 104052 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_2_Right_166
timestamp 1
transform -1 0 108836 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_1_Left_394
timestamp 1
transform 1 0 1104 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_1_Right_825
timestamp 1
transform -1 0 7912 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_2_Left_718
timestamp 1
transform 1 0 104052 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_2_Right_167
timestamp 1
transform -1 0 108836 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_1_Left_395
timestamp 1
transform 1 0 1104 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_1_Right_826
timestamp 1
transform -1 0 7912 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_2_Left_719
timestamp 1
transform 1 0 104052 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_2_Right_168
timestamp 1
transform -1 0 108836 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_1_Left_396
timestamp 1
transform 1 0 1104 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_1_Right_827
timestamp 1
transform -1 0 7912 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_2_Left_720
timestamp 1
transform 1 0 104052 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_2_Right_169
timestamp 1
transform -1 0 108836 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_1_Left_397
timestamp 1
transform 1 0 1104 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_1_Right_828
timestamp 1
transform -1 0 7912 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_2_Left_721
timestamp 1
transform 1 0 104052 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_2_Right_170
timestamp 1
transform -1 0 108836 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_1_Left_398
timestamp 1
transform 1 0 1104 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_1_Right_829
timestamp 1
transform -1 0 7912 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_2_Left_722
timestamp 1
transform 1 0 104052 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_2_Right_171
timestamp 1
transform -1 0 108836 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_1_Left_399
timestamp 1
transform 1 0 1104 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_1_Right_830
timestamp 1
transform -1 0 7912 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_2_Left_723
timestamp 1
transform 1 0 104052 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_2_Right_172
timestamp 1
transform -1 0 108836 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_1_Left_400
timestamp 1
transform 1 0 1104 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_1_Right_831
timestamp 1
transform -1 0 7912 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_2_Left_724
timestamp 1
transform 1 0 104052 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_2_Right_173
timestamp 1
transform -1 0 108836 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_1_Left_401
timestamp 1
transform 1 0 1104 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_1_Right_832
timestamp 1
transform -1 0 7912 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_2_Left_725
timestamp 1
transform 1 0 104052 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_2_Right_174
timestamp 1
transform -1 0 108836 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_1_Left_402
timestamp 1
transform 1 0 1104 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_1_Right_833
timestamp 1
transform -1 0 7912 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_2_Left_726
timestamp 1
transform 1 0 104052 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_2_Right_175
timestamp 1
transform -1 0 108836 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_1_Left_403
timestamp 1
transform 1 0 1104 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_1_Right_834
timestamp 1
transform -1 0 7912 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_2_Left_727
timestamp 1
transform 1 0 104052 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_2_Right_176
timestamp 1
transform -1 0 108836 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_1_Left_404
timestamp 1
transform 1 0 1104 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_1_Right_835
timestamp 1
transform -1 0 7912 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_2_Left_728
timestamp 1
transform 1 0 104052 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_2_Right_177
timestamp 1
transform -1 0 108836 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_1_Left_405
timestamp 1
transform 1 0 1104 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_1_Right_836
timestamp 1
transform -1 0 7912 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_2_Left_729
timestamp 1
transform 1 0 104052 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_2_Right_178
timestamp 1
transform -1 0 108836 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_1_Left_406
timestamp 1
transform 1 0 1104 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_1_Right_837
timestamp 1
transform -1 0 7912 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_2_Left_730
timestamp 1
transform 1 0 104052 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_2_Right_179
timestamp 1
transform -1 0 108836 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_1_Left_407
timestamp 1
transform 1 0 1104 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_1_Right_838
timestamp 1
transform -1 0 7912 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_2_Left_731
timestamp 1
transform 1 0 104052 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_2_Right_180
timestamp 1
transform -1 0 108836 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_1_Left_408
timestamp 1
transform 1 0 1104 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_1_Right_839
timestamp 1
transform -1 0 7912 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_2_Left_732
timestamp 1
transform 1 0 104052 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_2_Right_181
timestamp 1
transform -1 0 108836 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_1_Left_409
timestamp 1
transform 1 0 1104 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_1_Right_840
timestamp 1
transform -1 0 7912 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_2_Left_733
timestamp 1
transform 1 0 104052 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_2_Right_182
timestamp 1
transform -1 0 108836 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_1_Left_410
timestamp 1
transform 1 0 1104 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_1_Right_841
timestamp 1
transform -1 0 7912 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_2_Left_734
timestamp 1
transform 1 0 104052 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_2_Right_183
timestamp 1
transform -1 0 108836 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_1_Left_411
timestamp 1
transform 1 0 1104 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_1_Right_842
timestamp 1
transform -1 0 7912 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_2_Left_735
timestamp 1
transform 1 0 104052 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_2_Right_184
timestamp 1
transform -1 0 108836 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_1_Left_412
timestamp 1
transform 1 0 1104 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_1_Right_843
timestamp 1
transform -1 0 7912 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_2_Left_736
timestamp 1
transform 1 0 104052 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_2_Right_185
timestamp 1
transform -1 0 108836 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_1_Left_413
timestamp 1
transform 1 0 1104 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_1_Right_844
timestamp 1
transform -1 0 7912 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_2_Left_737
timestamp 1
transform 1 0 104052 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_2_Right_186
timestamp 1
transform -1 0 108836 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_1_Left_414
timestamp 1
transform 1 0 1104 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_1_Right_845
timestamp 1
transform -1 0 7912 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_2_Left_738
timestamp 1
transform 1 0 104052 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_2_Right_187
timestamp 1
transform -1 0 108836 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_1_Left_415
timestamp 1
transform 1 0 1104 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_1_Right_846
timestamp 1
transform -1 0 7912 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_2_Left_739
timestamp 1
transform 1 0 104052 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_2_Right_188
timestamp 1
transform -1 0 108836 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_1_Left_416
timestamp 1
transform 1 0 1104 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_1_Right_847
timestamp 1
transform -1 0 7912 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_2_Left_740
timestamp 1
transform 1 0 104052 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_2_Right_189
timestamp 1
transform -1 0 108836 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_1_Left_417
timestamp 1
transform 1 0 1104 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_1_Right_848
timestamp 1
transform -1 0 7912 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_2_Left_741
timestamp 1
transform 1 0 104052 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_2_Right_190
timestamp 1
transform -1 0 108836 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_1_Left_418
timestamp 1
transform 1 0 1104 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_1_Right_849
timestamp 1
transform -1 0 7912 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_2_Left_742
timestamp 1
transform 1 0 104052 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_2_Right_191
timestamp 1
transform -1 0 108836 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_1_Left_419
timestamp 1
transform 1 0 1104 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_1_Right_850
timestamp 1
transform -1 0 7912 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_2_Left_743
timestamp 1
transform 1 0 104052 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_2_Right_192
timestamp 1
transform -1 0 108836 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_1_Left_420
timestamp 1
transform 1 0 1104 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_1_Right_851
timestamp 1
transform -1 0 7912 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_2_Left_744
timestamp 1
transform 1 0 104052 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_2_Right_193
timestamp 1
transform -1 0 108836 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_1_Left_421
timestamp 1
transform 1 0 1104 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_1_Right_852
timestamp 1
transform -1 0 7912 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_2_Left_745
timestamp 1
transform 1 0 104052 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_2_Right_194
timestamp 1
transform -1 0 108836 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_1_Left_422
timestamp 1
transform 1 0 1104 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_1_Right_853
timestamp 1
transform -1 0 7912 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_2_Left_746
timestamp 1
transform 1 0 104052 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_2_Right_195
timestamp 1
transform -1 0 108836 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_1_Left_423
timestamp 1
transform 1 0 1104 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_1_Right_854
timestamp 1
transform -1 0 7912 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_2_Left_747
timestamp 1
transform 1 0 104052 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_2_Right_196
timestamp 1
transform -1 0 108836 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_1_Left_424
timestamp 1
transform 1 0 1104 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_1_Right_855
timestamp 1
transform -1 0 7912 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_2_Left_748
timestamp 1
transform 1 0 104052 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_2_Right_197
timestamp 1
transform -1 0 108836 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_1_Left_425
timestamp 1
transform 1 0 1104 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_1_Right_856
timestamp 1
transform -1 0 7912 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_2_Left_749
timestamp 1
transform 1 0 104052 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_2_Right_198
timestamp 1
transform -1 0 108836 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_1_Left_426
timestamp 1
transform 1 0 1104 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_1_Right_857
timestamp 1
transform -1 0 7912 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_2_Left_750
timestamp 1
transform 1 0 104052 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_2_Right_199
timestamp 1
transform -1 0 108836 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_1_Left_427
timestamp 1
transform 1 0 1104 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_1_Right_858
timestamp 1
transform -1 0 7912 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_2_Left_751
timestamp 1
transform 1 0 104052 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_2_Right_200
timestamp 1
transform -1 0 108836 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_1_Left_428
timestamp 1
transform 1 0 1104 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_1_Right_859
timestamp 1
transform -1 0 7912 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_2_Left_752
timestamp 1
transform 1 0 104052 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_2_Right_201
timestamp 1
transform -1 0 108836 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_1_Left_429
timestamp 1
transform 1 0 1104 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_1_Right_860
timestamp 1
transform -1 0 7912 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_2_Left_753
timestamp 1
transform 1 0 104052 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_2_Right_202
timestamp 1
transform -1 0 108836 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_1_Left_430
timestamp 1
transform 1 0 1104 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_1_Right_861
timestamp 1
transform -1 0 7912 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_2_Left_754
timestamp 1
transform 1 0 104052 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_2_Right_203
timestamp 1
transform -1 0 108836 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_1_Left_431
timestamp 1
transform 1 0 1104 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_1_Right_862
timestamp 1
transform -1 0 7912 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_2_Left_755
timestamp 1
transform 1 0 104052 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_2_Right_204
timestamp 1
transform -1 0 108836 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_1_Left_432
timestamp 1
transform 1 0 1104 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_1_Right_863
timestamp 1
transform -1 0 7912 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_2_Left_756
timestamp 1
transform 1 0 104052 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_2_Right_205
timestamp 1
transform -1 0 108836 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_1_Left_433
timestamp 1
transform 1 0 1104 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_1_Right_864
timestamp 1
transform -1 0 7912 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_2_Left_757
timestamp 1
transform 1 0 104052 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_2_Right_206
timestamp 1
transform -1 0 108836 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_1_Left_434
timestamp 1
transform 1 0 1104 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_1_Right_865
timestamp 1
transform -1 0 7912 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_2_Left_758
timestamp 1
transform 1 0 104052 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_2_Right_207
timestamp 1
transform -1 0 108836 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_1_Left_435
timestamp 1
transform 1 0 1104 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_1_Right_866
timestamp 1
transform -1 0 7912 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_2_Left_759
timestamp 1
transform 1 0 104052 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_2_Right_208
timestamp 1
transform -1 0 108836 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_1_Left_436
timestamp 1
transform 1 0 1104 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_1_Right_867
timestamp 1
transform -1 0 7912 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_2_Left_760
timestamp 1
transform 1 0 104052 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_2_Right_209
timestamp 1
transform -1 0 108836 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_1_Left_437
timestamp 1
transform 1 0 1104 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_1_Right_868
timestamp 1
transform -1 0 7912 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_2_Left_761
timestamp 1
transform 1 0 104052 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_2_Right_210
timestamp 1
transform -1 0 108836 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_1_Left_438
timestamp 1
transform 1 0 1104 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_1_Right_869
timestamp 1
transform -1 0 7912 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_2_Left_762
timestamp 1
transform 1 0 104052 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_2_Right_211
timestamp 1
transform -1 0 108836 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_1_Left_439
timestamp 1
transform 1 0 1104 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_1_Right_870
timestamp 1
transform -1 0 7912 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_2_Left_763
timestamp 1
transform 1 0 104052 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_2_Right_212
timestamp 1
transform -1 0 108836 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_1_Left_440
timestamp 1
transform 1 0 1104 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_1_Right_871
timestamp 1
transform -1 0 7912 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_2_Left_764
timestamp 1
transform 1 0 104052 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_2_Right_213
timestamp 1
transform -1 0 108836 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_1_Left_441
timestamp 1
transform 1 0 1104 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_1_Right_872
timestamp 1
transform -1 0 7912 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_2_Left_765
timestamp 1
transform 1 0 104052 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_2_Right_214
timestamp 1
transform -1 0 108836 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_1_Left_442
timestamp 1
transform 1 0 1104 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_1_Right_873
timestamp 1
transform -1 0 7912 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_2_Left_766
timestamp 1
transform 1 0 104052 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_2_Right_215
timestamp 1
transform -1 0 108836 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_1_Left_443
timestamp 1
transform 1 0 1104 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_1_Right_874
timestamp 1
transform -1 0 7912 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_2_Left_767
timestamp 1
transform 1 0 104052 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_2_Right_216
timestamp 1
transform -1 0 108836 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_1_Left_444
timestamp 1
transform 1 0 1104 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_1_Right_875
timestamp 1
transform -1 0 7912 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_2_Left_768
timestamp 1
transform 1 0 104052 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_2_Right_217
timestamp 1
transform -1 0 108836 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_1_Left_445
timestamp 1
transform 1 0 1104 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_1_Right_876
timestamp 1
transform -1 0 7912 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_2_Left_769
timestamp 1
transform 1 0 104052 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_2_Right_218
timestamp 1
transform -1 0 108836 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_1_Left_446
timestamp 1
transform 1 0 1104 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_1_Right_877
timestamp 1
transform -1 0 7912 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_2_Left_770
timestamp 1
transform 1 0 104052 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_2_Right_219
timestamp 1
transform -1 0 108836 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_1_Left_447
timestamp 1
transform 1 0 1104 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_1_Right_878
timestamp 1
transform -1 0 7912 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_2_Left_771
timestamp 1
transform 1 0 104052 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_2_Right_220
timestamp 1
transform -1 0 108836 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_1_Left_448
timestamp 1
transform 1 0 1104 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_1_Right_879
timestamp 1
transform -1 0 7912 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_2_Left_772
timestamp 1
transform 1 0 104052 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_2_Right_221
timestamp 1
transform -1 0 108836 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_1_Left_449
timestamp 1
transform 1 0 1104 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_1_Right_880
timestamp 1
transform -1 0 7912 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_2_Left_773
timestamp 1
transform 1 0 104052 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_2_Right_222
timestamp 1
transform -1 0 108836 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_1_Left_450
timestamp 1
transform 1 0 1104 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_1_Right_881
timestamp 1
transform -1 0 7912 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_2_Left_774
timestamp 1
transform 1 0 104052 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_2_Right_223
timestamp 1
transform -1 0 108836 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_1_Left_451
timestamp 1
transform 1 0 1104 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_1_Right_882
timestamp 1
transform -1 0 7912 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_2_Left_775
timestamp 1
transform 1 0 104052 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_2_Right_224
timestamp 1
transform -1 0 108836 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_1_Left_452
timestamp 1
transform 1 0 1104 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_1_Right_883
timestamp 1
transform -1 0 7912 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_2_Left_776
timestamp 1
transform 1 0 104052 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_2_Right_225
timestamp 1
transform -1 0 108836 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_1_Left_453
timestamp 1
transform 1 0 1104 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_1_Right_884
timestamp 1
transform -1 0 7912 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_2_Left_777
timestamp 1
transform 1 0 104052 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_2_Right_226
timestamp 1
transform -1 0 108836 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_1_Left_454
timestamp 1
transform 1 0 1104 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_1_Right_885
timestamp 1
transform -1 0 7912 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_2_Left_778
timestamp 1
transform 1 0 104052 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_2_Right_227
timestamp 1
transform -1 0 108836 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_1_Left_455
timestamp 1
transform 1 0 1104 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_1_Right_886
timestamp 1
transform -1 0 7912 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_2_Left_779
timestamp 1
transform 1 0 104052 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_2_Right_228
timestamp 1
transform -1 0 108836 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_1_Left_456
timestamp 1
transform 1 0 1104 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_1_Right_887
timestamp 1
transform -1 0 7912 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_2_Left_780
timestamp 1
transform 1 0 104052 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_2_Right_229
timestamp 1
transform -1 0 108836 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_228_Left_457
timestamp 1
transform 1 0 1104 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_228_Right_14
timestamp 1
transform -1 0 108836 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_229_Left_458
timestamp 1
transform 1 0 1104 0 -1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_229_Right_15
timestamp 1
transform -1 0 108836 0 -1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_888
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_889
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_890
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_891
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_892
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_893
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_894
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_895
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_896
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_897
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_898
timestamp 1
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_899
timestamp 1
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_900
timestamp 1
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_901
timestamp 1
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_902
timestamp 1
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_903
timestamp 1
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_904
timestamp 1
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_905
timestamp 1
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_906
timestamp 1
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_907
timestamp 1
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_908
timestamp 1
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_909
timestamp 1
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_910
timestamp 1
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_911
timestamp 1
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_912
timestamp 1
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_913
timestamp 1
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_914
timestamp 1
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_915
timestamp 1
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_916
timestamp 1
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_917
timestamp 1
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_918
timestamp 1
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_919
timestamp 1
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_920
timestamp 1
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_921
timestamp 1
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_922
timestamp 1
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_923
timestamp 1
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_924
timestamp 1
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_925
timestamp 1
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_926
timestamp 1
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_927
timestamp 1
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_928
timestamp 1
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_929
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_930
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_931
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_932
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_933
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_934
timestamp 1
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_935
timestamp 1
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_936
timestamp 1
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_937
timestamp 1
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_938
timestamp 1
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_939
timestamp 1
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_940
timestamp 1
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_941
timestamp 1
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_942
timestamp 1
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_943
timestamp 1
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_944
timestamp 1
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_945
timestamp 1
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_946
timestamp 1
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_947
timestamp 1
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_948
timestamp 1
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_949
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_950
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_951
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_952
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_953
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_954
timestamp 1
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_955
timestamp 1
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_956
timestamp 1
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_957
timestamp 1
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_958
timestamp 1
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_959
timestamp 1
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_960
timestamp 1
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_961
timestamp 1
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_962
timestamp 1
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_963
timestamp 1
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_964
timestamp 1
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_965
timestamp 1
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_966
timestamp 1
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_967
timestamp 1
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_968
timestamp 1
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_969
timestamp 1
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_970
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_971
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_972
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_973
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_974
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_975
timestamp 1
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_976
timestamp 1
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_977
timestamp 1
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_978
timestamp 1
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_979
timestamp 1
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_980
timestamp 1
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_981
timestamp 1
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_982
timestamp 1
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_983
timestamp 1
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_984
timestamp 1
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_985
timestamp 1
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_986
timestamp 1
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_987
timestamp 1
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_988
timestamp 1
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_989
timestamp 1
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_990
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_991
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_992
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_993
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_994
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_995
timestamp 1
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_996
timestamp 1
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_997
timestamp 1
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_998
timestamp 1
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_999
timestamp 1
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1000
timestamp 1
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1001
timestamp 1
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1002
timestamp 1
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1003
timestamp 1
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1004
timestamp 1
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1005
timestamp 1
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1006
timestamp 1
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1007
timestamp 1
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1008
timestamp 1
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1009
timestamp 1
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1010
timestamp 1
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1011
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1012
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1013
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1014
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1015
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1016
timestamp 1
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1017
timestamp 1
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1018
timestamp 1
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1019
timestamp 1
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1020
timestamp 1
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1021
timestamp 1
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1022
timestamp 1
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1023
timestamp 1
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1024
timestamp 1
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1025
timestamp 1
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1026
timestamp 1
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1027
timestamp 1
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1028
timestamp 1
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1029
timestamp 1
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1030
timestamp 1
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1031
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1032
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1033
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1034
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1035
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1036
timestamp 1
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1037
timestamp 1
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1038
timestamp 1
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1039
timestamp 1
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1040
timestamp 1
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1041
timestamp 1
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1042
timestamp 1
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1043
timestamp 1
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1044
timestamp 1
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1045
timestamp 1
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1046
timestamp 1
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1047
timestamp 1
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1048
timestamp 1
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1049
timestamp 1
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1050
timestamp 1
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1051
timestamp 1
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1052
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1053
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1054
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1055
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1056
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1057
timestamp 1
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1058
timestamp 1
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1059
timestamp 1
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1060
timestamp 1
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1061
timestamp 1
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1062
timestamp 1
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1063
timestamp 1
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1064
timestamp 1
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1065
timestamp 1
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1066
timestamp 1
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1067
timestamp 1
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1068
timestamp 1
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1069
timestamp 1
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1070
timestamp 1
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1071
timestamp 1
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1072
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1073
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1074
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1075
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1076
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1077
timestamp 1
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1078
timestamp 1
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1079
timestamp 1
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1080
timestamp 1
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1081
timestamp 1
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1082
timestamp 1
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1083
timestamp 1
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1084
timestamp 1
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1085
timestamp 1
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1086
timestamp 1
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1087
timestamp 1
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1088
timestamp 1
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1089
timestamp 1
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1090
timestamp 1
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1091
timestamp 1
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1092
timestamp 1
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1093
timestamp 1
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1094
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1095
timestamp 1
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1096
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1097
timestamp 1
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1098
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1099
timestamp 1
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1100
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1101
timestamp 1
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1102
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1103
timestamp 1
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1104
timestamp 1
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1105
timestamp 1
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1106
timestamp 1
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1107
timestamp 1
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1108
timestamp 1
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1109
timestamp 1
transform 1 0 44896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1110
timestamp 1
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1111
timestamp 1
transform 1 0 50048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1112
timestamp 1
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1113
timestamp 1
transform 1 0 55200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1114
timestamp 1
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1115
timestamp 1
transform 1 0 60352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1116
timestamp 1
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1117
timestamp 1
transform 1 0 65504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1118
timestamp 1
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1119
timestamp 1
transform 1 0 70656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1120
timestamp 1
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1121
timestamp 1
transform 1 0 75808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1122
timestamp 1
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1123
timestamp 1
transform 1 0 80960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1124
timestamp 1
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1125
timestamp 1
transform 1 0 86112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1126
timestamp 1
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1127
timestamp 1
transform 1 0 91264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1128
timestamp 1
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1129
timestamp 1
transform 1 0 96416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1130
timestamp 1
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1131
timestamp 1
transform 1 0 101568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1132
timestamp 1
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1133
timestamp 1
transform 1 0 106720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_1552
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_1553
timestamp 1
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_1_1134
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_1135
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_1554
timestamp 1
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_1_1136
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_1_1137
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_1555
timestamp 1
transform 1 0 106628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_1_1138
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_1_1139
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_1556
timestamp 1
transform 1 0 106628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_1_1140
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_1_1141
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_1557
timestamp 1
transform 1 0 106628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_1_1142
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_1_1143
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_1558
timestamp 1
transform 1 0 106628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_1_1144
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_1_1145
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_1559
timestamp 1
transform 1 0 106628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_1_1146
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_1_1147
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_1560
timestamp 1
transform 1 0 106628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_1_1148
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_1_1149
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_1561
timestamp 1
transform 1 0 106628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_1_1150
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_1_1151
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_1562
timestamp 1
transform 1 0 106628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_1_1152
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_1_1153
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_1563
timestamp 1
transform 1 0 106628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_1_1154
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_1_1155
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_1564
timestamp 1
transform 1 0 106628 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_1_1156
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_1_1157
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_1565
timestamp 1
transform 1 0 106628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_1_1158
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_1_1159
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_1566
timestamp 1
transform 1 0 106628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_1_1160
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_1_1161
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_1567
timestamp 1
transform 1 0 106628 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_1_1162
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_1_1163
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_1568
timestamp 1
transform 1 0 106628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_1_1164
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_1_1165
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_1569
timestamp 1
transform 1 0 106628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_1_1166
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_1_1167
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_1570
timestamp 1
transform 1 0 106628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_1_1168
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_1_1169
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_1571
timestamp 1
transform 1 0 106628 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_1_1170
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1_1171
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_1572
timestamp 1
transform 1 0 106628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1_1172
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1_1173
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_1573
timestamp 1
transform 1 0 106628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1_1174
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1_1175
timestamp 1
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_1574
timestamp 1
transform 1 0 106628 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1_1176
timestamp 1
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1_1177
timestamp 1
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_1575
timestamp 1
transform 1 0 106628 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1_1178
timestamp 1
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1_1179
timestamp 1
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_1576
timestamp 1
transform 1 0 106628 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1_1180
timestamp 1
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1_1181
timestamp 1
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_1577
timestamp 1
transform 1 0 106628 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1_1182
timestamp 1
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1_1183
timestamp 1
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_1578
timestamp 1
transform 1 0 106628 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1_1184
timestamp 1
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1_1185
timestamp 1
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_1579
timestamp 1
transform 1 0 106628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1_1186
timestamp 1
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1_1187
timestamp 1
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_1580
timestamp 1
transform 1 0 106628 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1_1188
timestamp 1
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1_1189
timestamp 1
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_1581
timestamp 1
transform 1 0 106628 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1_1190
timestamp 1
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1_1191
timestamp 1
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_1582
timestamp 1
transform 1 0 106628 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1_1192
timestamp 1
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1_1193
timestamp 1
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_1583
timestamp 1
transform 1 0 106628 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1_1194
timestamp 1
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1_1195
timestamp 1
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_1584
timestamp 1
transform 1 0 106628 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1_1196
timestamp 1
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1_1197
timestamp 1
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_1585
timestamp 1
transform 1 0 106628 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1_1198
timestamp 1
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1_1199
timestamp 1
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_1586
timestamp 1
transform 1 0 106628 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1_1200
timestamp 1
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1_1201
timestamp 1
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_1587
timestamp 1
transform 1 0 106628 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1_1202
timestamp 1
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1_1203
timestamp 1
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_1588
timestamp 1
transform 1 0 106628 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1_1204
timestamp 1
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1_1205
timestamp 1
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_1589
timestamp 1
transform 1 0 106628 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1_1206
timestamp 1
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1_1207
timestamp 1
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_1590
timestamp 1
transform 1 0 106628 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1_1208
timestamp 1
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1_1209
timestamp 1
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_1591
timestamp 1
transform 1 0 106628 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1_1210
timestamp 1
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1_1211
timestamp 1
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_1592
timestamp 1
transform 1 0 106628 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1_1212
timestamp 1
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1_1213
timestamp 1
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_1593
timestamp 1
transform 1 0 106628 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1_1214
timestamp 1
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1_1215
timestamp 1
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_1594
timestamp 1
transform 1 0 106628 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1_1216
timestamp 1
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1_1217
timestamp 1
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_1595
timestamp 1
transform 1 0 106628 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1_1218
timestamp 1
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1_1219
timestamp 1
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_1596
timestamp 1
transform 1 0 106628 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1_1220
timestamp 1
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1_1221
timestamp 1
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_1597
timestamp 1
transform 1 0 106628 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1_1222
timestamp 1
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1_1223
timestamp 1
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_1598
timestamp 1
transform 1 0 106628 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1_1224
timestamp 1
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1_1225
timestamp 1
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_1599
timestamp 1
transform 1 0 106628 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1_1226
timestamp 1
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1_1227
timestamp 1
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_1600
timestamp 1
transform 1 0 106628 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1_1228
timestamp 1
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1_1229
timestamp 1
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_1601
timestamp 1
transform 1 0 106628 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1_1230
timestamp 1
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1_1231
timestamp 1
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_1602
timestamp 1
transform 1 0 106628 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1_1232
timestamp 1
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1_1233
timestamp 1
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_1603
timestamp 1
transform 1 0 106628 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1_1234
timestamp 1
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1_1235
timestamp 1
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_1604
timestamp 1
transform 1 0 106628 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1_1236
timestamp 1
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1_1237
timestamp 1
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_1605
timestamp 1
transform 1 0 106628 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1_1238
timestamp 1
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1_1239
timestamp 1
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_1606
timestamp 1
transform 1 0 106628 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1241
timestamp 1
transform 1 0 3680 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1242
timestamp 1
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1243
timestamp 1
transform 1 0 8832 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1244
timestamp 1
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1245
timestamp 1
transform 1 0 13984 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1246
timestamp 1
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1247
timestamp 1
transform 1 0 19136 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1248
timestamp 1
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1249
timestamp 1
transform 1 0 24288 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1250
timestamp 1
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1251
timestamp 1
transform 1 0 29440 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1252
timestamp 1
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1253
timestamp 1
transform 1 0 34592 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1254
timestamp 1
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1255
timestamp 1
transform 1 0 39744 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1256
timestamp 1
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1257
timestamp 1
transform 1 0 44896 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1258
timestamp 1
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1259
timestamp 1
transform 1 0 50048 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1260
timestamp 1
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1261
timestamp 1
transform 1 0 55200 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1262
timestamp 1
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1263
timestamp 1
transform 1 0 60352 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1264
timestamp 1
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1265
timestamp 1
transform 1 0 65504 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1266
timestamp 1
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1267
timestamp 1
transform 1 0 70656 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1268
timestamp 1
transform 1 0 73232 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1269
timestamp 1
transform 1 0 75808 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1270
timestamp 1
transform 1 0 78384 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1271
timestamp 1
transform 1 0 80960 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1272
timestamp 1
transform 1 0 83536 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1273
timestamp 1
transform 1 0 86112 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1274
timestamp 1
transform 1 0 88688 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1275
timestamp 1
transform 1 0 91264 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1276
timestamp 1
transform 1 0 93840 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1277
timestamp 1
transform 1 0 96416 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1278
timestamp 1
transform 1 0 98992 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1279
timestamp 1
transform 1 0 101568 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1280
timestamp 1
transform 1 0 104144 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1281
timestamp 1
transform 1 0 106720 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1282
timestamp 1
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1283
timestamp 1
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1284
timestamp 1
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1285
timestamp 1
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1286
timestamp 1
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1287
timestamp 1
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1288
timestamp 1
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1289
timestamp 1
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1290
timestamp 1
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1291
timestamp 1
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1292
timestamp 1
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1293
timestamp 1
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1294
timestamp 1
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1295
timestamp 1
transform 1 0 70656 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1296
timestamp 1
transform 1 0 75808 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1297
timestamp 1
transform 1 0 80960 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1298
timestamp 1
transform 1 0 86112 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1299
timestamp 1
transform 1 0 91264 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1300
timestamp 1
transform 1 0 96416 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1301
timestamp 1
transform 1 0 101568 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1302
timestamp 1
transform 1 0 106720 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1303
timestamp 1
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1304
timestamp 1
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1305
timestamp 1
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1306
timestamp 1
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1307
timestamp 1
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1308
timestamp 1
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1309
timestamp 1
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1310
timestamp 1
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1311
timestamp 1
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1312
timestamp 1
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1313
timestamp 1
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1314
timestamp 1
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1315
timestamp 1
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1316
timestamp 1
transform 1 0 73232 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1317
timestamp 1
transform 1 0 78384 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1318
timestamp 1
transform 1 0 83536 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1319
timestamp 1
transform 1 0 88688 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1320
timestamp 1
transform 1 0 93840 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1321
timestamp 1
transform 1 0 98992 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1322
timestamp 1
transform 1 0 104144 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1323
timestamp 1
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1324
timestamp 1
transform 1 0 6256 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1325
timestamp 1
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1326
timestamp 1
transform 1 0 11408 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1327
timestamp 1
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1328
timestamp 1
transform 1 0 16560 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1329
timestamp 1
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1330
timestamp 1
transform 1 0 21712 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1331
timestamp 1
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1332
timestamp 1
transform 1 0 26864 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1333
timestamp 1
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1334
timestamp 1
transform 1 0 32016 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1335
timestamp 1
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1336
timestamp 1
transform 1 0 37168 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1337
timestamp 1
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1338
timestamp 1
transform 1 0 42320 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1339
timestamp 1
transform 1 0 44896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1340
timestamp 1
transform 1 0 47472 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1341
timestamp 1
transform 1 0 50048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1342
timestamp 1
transform 1 0 52624 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1343
timestamp 1
transform 1 0 55200 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1344
timestamp 1
transform 1 0 57776 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1345
timestamp 1
transform 1 0 60352 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1346
timestamp 1
transform 1 0 62928 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1347
timestamp 1
transform 1 0 65504 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1348
timestamp 1
transform 1 0 68080 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1349
timestamp 1
transform 1 0 70656 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1350
timestamp 1
transform 1 0 73232 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1351
timestamp 1
transform 1 0 75808 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1352
timestamp 1
transform 1 0 78384 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1353
timestamp 1
transform 1 0 80960 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1354
timestamp 1
transform 1 0 83536 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1355
timestamp 1
transform 1 0 86112 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1356
timestamp 1
transform 1 0 88688 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1357
timestamp 1
transform 1 0 91264 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1358
timestamp 1
transform 1 0 93840 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1359
timestamp 1
transform 1 0 96416 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1360
timestamp 1
transform 1 0 98992 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1361
timestamp 1
transform 1 0 101568 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1362
timestamp 1
transform 1 0 104144 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1363
timestamp 1
transform 1 0 106720 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1_1240
timestamp 1
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1_1364
timestamp 1
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2_1607
timestamp 1
transform 1 0 106628 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1_1365
timestamp 1
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1_1366
timestamp 1
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2_1608
timestamp 1
transform 1 0 106628 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1_1367
timestamp 1
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1_1368
timestamp 1
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2_1609
timestamp 1
transform 1 0 106628 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1_1369
timestamp 1
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1_1370
timestamp 1
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2_1610
timestamp 1
transform 1 0 106628 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1_1371
timestamp 1
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1_1372
timestamp 1
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2_1611
timestamp 1
transform 1 0 106628 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1_1373
timestamp 1
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1_1374
timestamp 1
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2_1612
timestamp 1
transform 1 0 106628 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1_1375
timestamp 1
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1_1376
timestamp 1
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2_1613
timestamp 1
transform 1 0 106628 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1_1377
timestamp 1
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1_1378
timestamp 1
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2_1614
timestamp 1
transform 1 0 106628 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1_1379
timestamp 1
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1_1380
timestamp 1
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2_1615
timestamp 1
transform 1 0 106628 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1_1381
timestamp 1
transform 1 0 6256 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1_1382
timestamp 1
transform 1 0 3680 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_1616
timestamp 1
transform 1 0 106628 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1_1383
timestamp 1
transform 1 0 6256 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1_1384
timestamp 1
transform 1 0 3680 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_1617
timestamp 1
transform 1 0 106628 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1_1385
timestamp 1
transform 1 0 6256 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1_1386
timestamp 1
transform 1 0 3680 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_1618
timestamp 1
transform 1 0 106628 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1_1387
timestamp 1
transform 1 0 6256 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1_1388
timestamp 1
transform 1 0 3680 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_1619
timestamp 1
transform 1 0 106628 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1_1389
timestamp 1
transform 1 0 6256 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1_1390
timestamp 1
transform 1 0 3680 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_1620
timestamp 1
transform 1 0 106628 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1_1391
timestamp 1
transform 1 0 6256 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1_1392
timestamp 1
transform 1 0 3680 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_1621
timestamp 1
transform 1 0 106628 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1_1393
timestamp 1
transform 1 0 6256 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1_1394
timestamp 1
transform 1 0 3680 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_1622
timestamp 1
transform 1 0 106628 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1_1395
timestamp 1
transform 1 0 6256 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1_1396
timestamp 1
transform 1 0 3680 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_1623
timestamp 1
transform 1 0 106628 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1_1397
timestamp 1
transform 1 0 6256 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1_1398
timestamp 1
transform 1 0 3680 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_2_1624
timestamp 1
transform 1 0 106628 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1_1399
timestamp 1
transform 1 0 6256 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1_1400
timestamp 1
transform 1 0 3680 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_2_1625
timestamp 1
transform 1 0 106628 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1_1401
timestamp 1
transform 1 0 6256 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1_1402
timestamp 1
transform 1 0 3680 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_2_1626
timestamp 1
transform 1 0 106628 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1_1403
timestamp 1
transform 1 0 6256 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1_1404
timestamp 1
transform 1 0 3680 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_2_1627
timestamp 1
transform 1 0 106628 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1_1405
timestamp 1
transform 1 0 6256 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1_1406
timestamp 1
transform 1 0 3680 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_2_1628
timestamp 1
transform 1 0 106628 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1_1407
timestamp 1
transform 1 0 6256 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1_1408
timestamp 1
transform 1 0 3680 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_2_1629
timestamp 1
transform 1 0 106628 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1_1409
timestamp 1
transform 1 0 6256 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1_1410
timestamp 1
transform 1 0 3680 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_2_1630
timestamp 1
transform 1 0 106628 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1_1411
timestamp 1
transform 1 0 6256 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1_1412
timestamp 1
transform 1 0 3680 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_2_1631
timestamp 1
transform 1 0 106628 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1_1413
timestamp 1
transform 1 0 6256 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1_1414
timestamp 1
transform 1 0 3680 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_2_1632
timestamp 1
transform 1 0 106628 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1_1415
timestamp 1
transform 1 0 6256 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1_1416
timestamp 1
transform 1 0 3680 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_2_1633
timestamp 1
transform 1 0 106628 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1_1417
timestamp 1
transform 1 0 6256 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1_1418
timestamp 1
transform 1 0 3680 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_2_1634
timestamp 1
transform 1 0 106628 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1_1419
timestamp 1
transform 1 0 6256 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1_1420
timestamp 1
transform 1 0 3680 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_2_1635
timestamp 1
transform 1 0 106628 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1_1421
timestamp 1
transform 1 0 6256 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_1_1422
timestamp 1
transform 1 0 3680 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2_1636
timestamp 1
transform 1 0 106628 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_1_1423
timestamp 1
transform 1 0 6256 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_1_1424
timestamp 1
transform 1 0 3680 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2_1637
timestamp 1
transform 1 0 106628 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_183_1_1425
timestamp 1
transform 1 0 6256 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_184_1_1426
timestamp 1
transform 1 0 3680 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_184_2_1638
timestamp 1
transform 1 0 106628 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_185_1_1427
timestamp 1
transform 1 0 6256 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_186_1_1428
timestamp 1
transform 1 0 3680 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_186_2_1639
timestamp 1
transform 1 0 106628 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_187_1_1429
timestamp 1
transform 1 0 6256 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_188_1_1430
timestamp 1
transform 1 0 3680 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_188_2_1640
timestamp 1
transform 1 0 106628 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_189_1_1431
timestamp 1
transform 1 0 6256 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_190_1_1432
timestamp 1
transform 1 0 3680 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_190_2_1641
timestamp 1
transform 1 0 106628 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_191_1_1433
timestamp 1
transform 1 0 6256 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_192_1_1434
timestamp 1
transform 1 0 3680 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_192_2_1642
timestamp 1
transform 1 0 106628 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_193_1_1435
timestamp 1
transform 1 0 6256 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_194_1_1436
timestamp 1
transform 1 0 3680 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_194_2_1643
timestamp 1
transform 1 0 106628 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_195_1_1437
timestamp 1
transform 1 0 6256 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_196_1_1438
timestamp 1
transform 1 0 3680 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_196_2_1644
timestamp 1
transform 1 0 106628 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_197_1_1439
timestamp 1
transform 1 0 6256 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_198_1_1440
timestamp 1
transform 1 0 3680 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_198_2_1645
timestamp 1
transform 1 0 106628 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_199_1_1441
timestamp 1
transform 1 0 6256 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_200_1_1442
timestamp 1
transform 1 0 3680 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_200_2_1646
timestamp 1
transform 1 0 106628 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_201_1_1443
timestamp 1
transform 1 0 6256 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_202_1_1444
timestamp 1
transform 1 0 3680 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_202_2_1647
timestamp 1
transform 1 0 106628 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_203_1_1445
timestamp 1
transform 1 0 6256 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_204_1_1446
timestamp 1
transform 1 0 3680 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_204_2_1648
timestamp 1
transform 1 0 106628 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_205_1_1447
timestamp 1
transform 1 0 6256 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_206_1_1448
timestamp 1
transform 1 0 3680 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_206_2_1649
timestamp 1
transform 1 0 106628 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_207_1_1449
timestamp 1
transform 1 0 6256 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_208_1_1450
timestamp 1
transform 1 0 3680 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_208_2_1650
timestamp 1
transform 1 0 106628 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_209_1_1451
timestamp 1
transform 1 0 6256 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_210_1_1452
timestamp 1
transform 1 0 3680 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_210_2_1651
timestamp 1
transform 1 0 106628 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_211_1_1453
timestamp 1
transform 1 0 6256 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_212_1_1454
timestamp 1
transform 1 0 3680 0 1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_212_2_1652
timestamp 1
transform 1 0 106628 0 1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_213_1_1455
timestamp 1
transform 1 0 6256 0 -1 118592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_214_1_1456
timestamp 1
transform 1 0 3680 0 1 118592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_214_2_1653
timestamp 1
transform 1 0 106628 0 1 118592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_215_1_1457
timestamp 1
transform 1 0 6256 0 -1 119680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_216_1_1458
timestamp 1
transform 1 0 3680 0 1 119680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_216_2_1654
timestamp 1
transform 1 0 106628 0 1 119680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_217_1_1459
timestamp 1
transform 1 0 6256 0 -1 120768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_218_1_1460
timestamp 1
transform 1 0 3680 0 1 120768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_218_2_1655
timestamp 1
transform 1 0 106628 0 1 120768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_219_1_1461
timestamp 1
transform 1 0 6256 0 -1 121856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_220_1_1462
timestamp 1
transform 1 0 3680 0 1 121856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_220_2_1656
timestamp 1
transform 1 0 106628 0 1 121856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_221_1_1463
timestamp 1
transform 1 0 6256 0 -1 122944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_222_1_1464
timestamp 1
transform 1 0 3680 0 1 122944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_222_2_1657
timestamp 1
transform 1 0 106628 0 1 122944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_223_1_1465
timestamp 1
transform 1 0 6256 0 -1 124032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_224_1_1466
timestamp 1
transform 1 0 3680 0 1 124032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_224_2_1658
timestamp 1
transform 1 0 106628 0 1 124032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_225_1_1467
timestamp 1
transform 1 0 6256 0 -1 125120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_226_1_1468
timestamp 1
transform 1 0 3680 0 1 125120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_226_2_1659
timestamp 1
transform 1 0 106628 0 1 125120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_227_1_1469
timestamp 1
transform 1 0 6256 0 -1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1470
timestamp 1
transform 1 0 3680 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1471
timestamp 1
transform 1 0 6256 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1472
timestamp 1
transform 1 0 8832 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1473
timestamp 1
transform 1 0 11408 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1474
timestamp 1
transform 1 0 13984 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1475
timestamp 1
transform 1 0 16560 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1476
timestamp 1
transform 1 0 19136 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1477
timestamp 1
transform 1 0 21712 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1478
timestamp 1
transform 1 0 24288 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1479
timestamp 1
transform 1 0 26864 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1480
timestamp 1
transform 1 0 29440 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1481
timestamp 1
transform 1 0 32016 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1482
timestamp 1
transform 1 0 34592 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1483
timestamp 1
transform 1 0 37168 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1484
timestamp 1
transform 1 0 39744 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1485
timestamp 1
transform 1 0 42320 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1486
timestamp 1
transform 1 0 44896 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1487
timestamp 1
transform 1 0 47472 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1488
timestamp 1
transform 1 0 50048 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1489
timestamp 1
transform 1 0 52624 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1490
timestamp 1
transform 1 0 55200 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1491
timestamp 1
transform 1 0 57776 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1492
timestamp 1
transform 1 0 60352 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1493
timestamp 1
transform 1 0 62928 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1494
timestamp 1
transform 1 0 65504 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1495
timestamp 1
transform 1 0 68080 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1496
timestamp 1
transform 1 0 70656 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1497
timestamp 1
transform 1 0 73232 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1498
timestamp 1
transform 1 0 75808 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1499
timestamp 1
transform 1 0 78384 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1500
timestamp 1
transform 1 0 80960 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1501
timestamp 1
transform 1 0 83536 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1502
timestamp 1
transform 1 0 86112 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1503
timestamp 1
transform 1 0 88688 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1504
timestamp 1
transform 1 0 91264 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1505
timestamp 1
transform 1 0 93840 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1506
timestamp 1
transform 1 0 96416 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1507
timestamp 1
transform 1 0 98992 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1508
timestamp 1
transform 1 0 101568 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1509
timestamp 1
transform 1 0 104144 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1510
timestamp 1
transform 1 0 106720 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1511
timestamp 1
transform 1 0 3680 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1512
timestamp 1
transform 1 0 6256 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1513
timestamp 1
transform 1 0 8832 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1514
timestamp 1
transform 1 0 11408 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1515
timestamp 1
transform 1 0 13984 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1516
timestamp 1
transform 1 0 16560 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1517
timestamp 1
transform 1 0 19136 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1518
timestamp 1
transform 1 0 21712 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1519
timestamp 1
transform 1 0 24288 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1520
timestamp 1
transform 1 0 26864 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1521
timestamp 1
transform 1 0 29440 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1522
timestamp 1
transform 1 0 32016 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1523
timestamp 1
transform 1 0 34592 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1524
timestamp 1
transform 1 0 37168 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1525
timestamp 1
transform 1 0 39744 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1526
timestamp 1
transform 1 0 42320 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1527
timestamp 1
transform 1 0 44896 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1528
timestamp 1
transform 1 0 47472 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1529
timestamp 1
transform 1 0 50048 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1530
timestamp 1
transform 1 0 52624 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1531
timestamp 1
transform 1 0 55200 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1532
timestamp 1
transform 1 0 57776 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1533
timestamp 1
transform 1 0 60352 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1534
timestamp 1
transform 1 0 62928 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1535
timestamp 1
transform 1 0 65504 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1536
timestamp 1
transform 1 0 68080 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1537
timestamp 1
transform 1 0 70656 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1538
timestamp 1
transform 1 0 73232 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1539
timestamp 1
transform 1 0 75808 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1540
timestamp 1
transform 1 0 78384 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1541
timestamp 1
transform 1 0 80960 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1542
timestamp 1
transform 1 0 83536 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1543
timestamp 1
transform 1 0 86112 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1544
timestamp 1
transform 1 0 88688 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1545
timestamp 1
transform 1 0 91264 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1546
timestamp 1
transform 1 0 93840 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1547
timestamp 1
transform 1 0 96416 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1548
timestamp 1
transform 1 0 98992 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1549
timestamp 1
transform 1 0 101568 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1550
timestamp 1
transform 1 0 104144 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1551
timestamp 1
transform 1 0 106720 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  wire68
timestamp 1
transform 1 0 61732 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire69
timestamp 1
transform 1 0 59248 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire70
timestamp 1
transform 1 0 58328 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire71
timestamp 1
transform -1 0 49864 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire72
timestamp 1
transform -1 0 48668 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire73
timestamp 1
transform -1 0 45356 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire74
timestamp 1
transform -1 0 41216 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire75
timestamp 1
transform 1 0 41216 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire76
timestamp 1
transform -1 0 37904 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire77
timestamp 1
transform 1 0 77188 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire78
timestamp 1
transform 1 0 71300 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire79
timestamp 1
transform 1 0 70196 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire80
timestamp 1
transform 1 0 66608 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire81
timestamp 1
transform 1 0 65596 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire82
timestamp 1
transform 1 0 63848 0 1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire83
timestamp 1
transform 1 0 35972 0 1 126208
box -38 -48 406 592
<< labels >>
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 addr00[0]
port 0 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 addr00[1]
port 1 nsew signal input
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 addr00[2]
port 2 nsew signal input
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 addr00[3]
port 3 nsew signal input
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 addr00[4]
port 4 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 addr00[5]
port 5 nsew signal input
flabel metal3 s 0 39448 800 39568 0 FreeSans 480 0 0 0 addr00[6]
port 6 nsew signal input
flabel metal3 s 0 41488 800 41608 0 FreeSans 480 0 0 0 addr00[7]
port 7 nsew signal input
flabel metal3 s 0 61208 800 61328 0 FreeSans 480 0 0 0 addr01[0]
port 8 nsew signal input
flabel metal3 s 0 70048 800 70168 0 FreeSans 480 0 0 0 addr01[1]
port 9 nsew signal input
flabel metal3 s 0 93848 800 93968 0 FreeSans 480 0 0 0 addr01[2]
port 10 nsew signal input
flabel metal3 s 0 95888 800 96008 0 FreeSans 480 0 0 0 addr01[3]
port 11 nsew signal input
flabel metal3 s 0 96568 800 96688 0 FreeSans 480 0 0 0 addr01[4]
port 12 nsew signal input
flabel metal3 s 0 98608 800 98728 0 FreeSans 480 0 0 0 addr01[5]
port 13 nsew signal input
flabel metal3 s 0 99288 800 99408 0 FreeSans 480 0 0 0 addr01[6]
port 14 nsew signal input
flabel metal3 s 0 101328 800 101448 0 FreeSans 480 0 0 0 addr01[7]
port 15 nsew signal input
flabel metal2 s 98550 129200 98606 130000 0 FreeSans 224 90 0 0 clk
port 16 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 csb00
port 17 nsew signal input
flabel metal3 s 0 75488 800 75608 0 FreeSans 480 0 0 0 csb01
port 18 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 din00[0]
port 19 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 din00[10]
port 20 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 din00[11]
port 21 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 din00[12]
port 22 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 din00[13]
port 23 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 din00[14]
port 24 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 din00[15]
port 25 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 din00[1]
port 26 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 din00[2]
port 27 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 din00[3]
port 28 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 din00[4]
port 29 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 din00[5]
port 30 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 din00[6]
port 31 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 din00[7]
port 32 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 din00[8]
port 33 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 din00[9]
port 34 nsew signal input
flabel metal3 s 0 68008 800 68128 0 FreeSans 480 0 0 0 din01[0]
port 35 nsew signal input
flabel metal3 s 0 69368 800 69488 0 FreeSans 480 0 0 0 din01[10]
port 36 nsew signal input
flabel metal3 s 0 71408 800 71528 0 FreeSans 480 0 0 0 din01[11]
port 37 nsew signal input
flabel metal3 s 0 72088 800 72208 0 FreeSans 480 0 0 0 din01[12]
port 38 nsew signal input
flabel metal3 s 0 72768 800 72888 0 FreeSans 480 0 0 0 din01[13]
port 39 nsew signal input
flabel metal3 s 0 68688 800 68808 0 FreeSans 480 0 0 0 din01[14]
port 40 nsew signal input
flabel metal3 s 0 73448 800 73568 0 FreeSans 480 0 0 0 din01[15]
port 41 nsew signal input
flabel metal3 s 0 74128 800 74248 0 FreeSans 480 0 0 0 din01[1]
port 42 nsew signal input
flabel metal3 s 0 61888 800 62008 0 FreeSans 480 0 0 0 din01[2]
port 43 nsew signal input
flabel metal3 s 0 76168 800 76288 0 FreeSans 480 0 0 0 din01[3]
port 44 nsew signal input
flabel metal3 s 0 67328 800 67448 0 FreeSans 480 0 0 0 din01[4]
port 45 nsew signal input
flabel metal3 s 0 76848 800 76968 0 FreeSans 480 0 0 0 din01[5]
port 46 nsew signal input
flabel metal3 s 0 77528 800 77648 0 FreeSans 480 0 0 0 din01[6]
port 47 nsew signal input
flabel metal3 s 0 70728 800 70848 0 FreeSans 480 0 0 0 din01[7]
port 48 nsew signal input
flabel metal3 s 0 74808 800 74928 0 FreeSans 480 0 0 0 din01[8]
port 49 nsew signal input
flabel metal3 s 0 78208 800 78328 0 FreeSans 480 0 0 0 din01[9]
port 50 nsew signal input
flabel metal3 s 109200 51008 110000 51128 0 FreeSans 480 0 0 0 rst
port 51 nsew signal input
flabel metal3 s 0 62568 800 62688 0 FreeSans 480 0 0 0 sine_out[0]
port 52 nsew signal output
flabel metal3 s 109200 63928 110000 64048 0 FreeSans 480 0 0 0 sine_out[10]
port 53 nsew signal output
flabel metal3 s 109200 69368 110000 69488 0 FreeSans 480 0 0 0 sine_out[11]
port 54 nsew signal output
flabel metal3 s 109200 65968 110000 66088 0 FreeSans 480 0 0 0 sine_out[12]
port 55 nsew signal output
flabel metal3 s 109200 65288 110000 65408 0 FreeSans 480 0 0 0 sine_out[13]
port 56 nsew signal output
flabel metal3 s 109200 68008 110000 68128 0 FreeSans 480 0 0 0 sine_out[14]
port 57 nsew signal output
flabel metal3 s 109200 67328 110000 67448 0 FreeSans 480 0 0 0 sine_out[15]
port 58 nsew signal output
flabel metal3 s 0 63928 800 64048 0 FreeSans 480 0 0 0 sine_out[1]
port 59 nsew signal output
flabel metal3 s 0 63248 800 63368 0 FreeSans 480 0 0 0 sine_out[2]
port 60 nsew signal output
flabel metal3 s 0 64608 800 64728 0 FreeSans 480 0 0 0 sine_out[3]
port 61 nsew signal output
flabel metal3 s 0 65968 800 66088 0 FreeSans 480 0 0 0 sine_out[4]
port 62 nsew signal output
flabel metal3 s 0 66648 800 66768 0 FreeSans 480 0 0 0 sine_out[5]
port 63 nsew signal output
flabel metal3 s 0 65288 800 65408 0 FreeSans 480 0 0 0 sine_out[6]
port 64 nsew signal output
flabel metal3 s 109200 64608 110000 64728 0 FreeSans 480 0 0 0 sine_out[7]
port 65 nsew signal output
flabel metal3 s 109200 66648 110000 66768 0 FreeSans 480 0 0 0 sine_out[8]
port 66 nsew signal output
flabel metal3 s 109200 68688 110000 68808 0 FreeSans 480 0 0 0 sine_out[9]
port 67 nsew signal output
flabel metal4 s 4208 2128 4528 127344 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 34928 2128 35248 7880 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 34928 65650 35248 67880 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 34928 125650 35248 127344 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 65648 2128 65968 8064 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 65648 65776 65968 68064 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 65648 125834 65968 127344 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 96368 2128 96688 8064 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 96368 65650 96688 68064 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 96368 125650 96688 127344 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal5 s 1056 5346 108884 5666 0 FreeSans 2560 0 0 0 vccd1
port 68 nsew power bidirectional
flabel metal5 s 1056 35982 108884 36302 0 FreeSans 2560 0 0 0 vccd1
port 68 nsew power bidirectional
flabel metal5 s 1056 66618 108884 66938 0 FreeSans 2560 0 0 0 vccd1
port 68 nsew power bidirectional
flabel metal5 s 1056 97254 108884 97574 0 FreeSans 2560 0 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 105916 7024 106236 66416 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 105916 67408 106236 126800 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal5 s 4208 125980 108884 126300 0 FreeSans 2560 0 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 4868 2128 5188 127344 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 8064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 35588 65650 35908 68064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 35588 125650 35908 127344 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 66308 2128 66628 8064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 66308 65650 66628 68064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 66308 125650 66628 127344 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 97028 2128 97348 8064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 97028 65650 97348 68064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 97028 125650 97348 127344 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal5 s 1056 6006 108884 6326 0 FreeSans 2560 0 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal5 s 1056 36642 108884 36962 0 FreeSans 2560 0 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal5 s 1056 67278 108884 67598 0 FreeSans 2560 0 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal5 s 1056 97914 108884 98234 0 FreeSans 2560 0 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 106652 7024 106972 66416 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 106652 67408 106972 126800 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal5 s 4208 126660 108884 126980 0 FreeSans 2560 0 0 0 vssd1
port 69 nsew ground bidirectional
rlabel via4 101806 97414 101806 97414 0 vccd1
rlabel via4 101110 98074 101110 98074 0 vssd1
rlabel metal1 33350 67320 33350 67320 0 _000_
rlabel metal2 85238 67082 85238 67082 0 _001_
rlabel metal2 74014 66708 74014 66708 0 _002_
rlabel metal2 89746 66572 89746 66572 0 _003_
rlabel metal2 75854 67082 75854 67082 0 _004_
rlabel metal1 75210 67286 75210 67286 0 _005_
rlabel metal1 86894 66470 86894 66470 0 _006_
rlabel metal2 32798 66266 32798 66266 0 _007_
rlabel metal2 32890 67320 32890 67320 0 _008_
rlabel metal2 24702 66946 24702 66946 0 _009_
rlabel metal1 21942 66504 21942 66504 0 _010_
rlabel metal1 44114 67048 44114 67048 0 _011_
rlabel metal2 44022 66912 44022 66912 0 _012_
rlabel metal2 70426 67031 70426 67031 0 _013_
rlabel metal2 79994 67184 79994 67184 0 _014_
rlabel metal2 75946 66096 75946 66096 0 _015_
rlabel metal1 91540 67150 91540 67150 0 _016_
rlabel metal1 105386 85578 105386 85578 0 _017_
rlabel via1 96823 65926 96823 65926 0 _018_
rlabel metal1 100004 65994 100004 65994 0 _019_
rlabel metal1 92138 66062 92138 66062 0 _020_
rlabel metal2 96094 65688 96094 65688 0 _021_
rlabel metal1 104788 45254 104788 45254 0 _022_
rlabel metal1 93196 66062 93196 66062 0 _023_
rlabel metal1 79258 66538 79258 66538 0 _024_
rlabel metal1 84134 66681 84134 66681 0 _025_
rlabel metal2 91770 66606 91770 66606 0 _026_
rlabel metal1 89861 66538 89861 66538 0 _027_
rlabel metal2 90298 66198 90298 66198 0 _028_
rlabel metal2 89746 66181 89746 66181 0 _029_
rlabel metal1 86848 66198 86848 66198 0 _030_
rlabel metal2 93610 67830 93610 67830 0 _031_
rlabel metal1 93157 66538 93157 66538 0 _032_
rlabel metal1 89654 67218 89654 67218 0 _033_
rlabel metal1 104512 80070 104512 80070 0 _034_
rlabel metal1 93702 68204 93702 68204 0 _035_
rlabel metal2 98210 67422 98210 67422 0 _036_
rlabel metal1 92046 67320 92046 67320 0 _037_
rlabel metal1 94477 66198 94477 66198 0 _038_
rlabel metal2 104742 41004 104742 41004 0 _039_
rlabel metal2 93518 67626 93518 67626 0 _040_
rlabel metal1 77142 67082 77142 67082 0 _041_
rlabel metal2 17342 66946 17342 66946 0 _042_
rlabel metal2 30590 66606 30590 66606 0 _043_
rlabel metal1 26680 66810 26680 66810 0 _044_
rlabel metal2 25806 66810 25806 66810 0 _045_
rlabel metal1 21673 66538 21673 66538 0 _046_
rlabel metal1 31878 66538 31878 66538 0 _047_
rlabel metal2 31050 66368 31050 66368 0 _048_
rlabel metal1 81551 67286 81551 67286 0 _049_
rlabel metal1 96002 67184 96002 67184 0 _050_
rlabel via1 104456 78642 104456 78642 0 _051_
rlabel metal1 104282 56882 104282 56882 0 _052_
rlabel metal1 101246 66130 101246 66130 0 _053_
rlabel metal1 104282 59534 104282 59534 0 _054_
rlabel metal1 103914 59602 103914 59602 0 _055_
rlabel metal2 104742 52224 104742 52224 0 _056_
rlabel metal1 104420 54842 104420 54842 0 _057_
rlabel metal1 105156 57018 105156 57018 0 _058_
rlabel metal2 23230 1520 23230 1520 0 addr00[0]
rlabel metal2 24518 1520 24518 1520 0 addr00[1]
rlabel metal2 1426 34323 1426 34323 0 addr00[2]
rlabel metal1 1380 35666 1380 35666 0 addr00[3]
rlabel metal2 1426 37009 1426 37009 0 addr00[4]
rlabel metal1 1334 38318 1334 38318 0 addr00[5]
rlabel metal2 1426 39763 1426 39763 0 addr00[6]
rlabel metal1 1334 41582 1334 41582 0 addr00[7]
rlabel metal1 1426 61778 1426 61778 0 addr01[0]
rlabel metal2 2254 70261 2254 70261 0 addr01[1]
rlabel metal1 1380 94418 1380 94418 0 addr01[2]
rlabel metal1 1334 95982 1334 95982 0 addr01[3]
rlabel metal1 1380 97070 1380 97070 0 addr01[4]
rlabel metal1 1380 98770 1380 98770 0 addr01[5]
rlabel metal2 1426 99603 1426 99603 0 addr01[6]
rlabel metal1 1334 101422 1334 101422 0 addr01[7]
rlabel metal1 100372 128350 100372 128350 0 clk
rlabel metal1 21574 66130 21574 66130 0 clknet_0_clk
rlabel metal1 17250 66130 17250 66130 0 clknet_2_0__leaf_clk
rlabel metal1 58006 66198 58006 66198 0 clknet_2_1__leaf_clk
rlabel metal1 106030 37978 106030 37978 0 clknet_2_2__leaf_clk
rlabel metal4 95890 123903 95890 123903 0 clknet_2_3__leaf_clk
rlabel metal1 1380 16082 1380 16082 0 csb00
rlabel metal2 1426 75735 1426 75735 0 csb01
rlabel metal2 25806 1520 25806 1520 0 din00[0]
rlabel metal2 37398 1520 37398 1520 0 din00[10]
rlabel metal2 38686 1520 38686 1520 0 din00[11]
rlabel metal2 39974 1520 39974 1520 0 din00[12]
rlabel metal2 41262 1520 41262 1520 0 din00[13]
rlabel metal2 41906 1520 41906 1520 0 din00[14]
rlabel metal2 43194 1520 43194 1520 0 din00[15]
rlabel metal2 27094 1520 27094 1520 0 din00[1]
rlabel metal2 28382 1520 28382 1520 0 din00[2]
rlabel metal2 29026 1520 29026 1520 0 din00[3]
rlabel metal2 30314 1520 30314 1520 0 din00[4]
rlabel metal2 31602 1520 31602 1520 0 din00[5]
rlabel metal2 32890 1520 32890 1520 0 din00[6]
rlabel metal2 34178 1520 34178 1520 0 din00[7]
rlabel metal2 35466 1520 35466 1520 0 din00[8]
rlabel metal2 36110 1520 36110 1520 0 din00[9]
rlabel metal1 1426 68306 1426 68306 0 din01[0]
rlabel metal1 1426 69802 1426 69802 0 din01[10]
rlabel metal1 1380 71570 1380 71570 0 din01[11]
rlabel metal1 1426 72658 1426 72658 0 din01[12]
rlabel metal2 1518 72947 1518 72947 0 din01[13]
rlabel metal1 1380 68714 1380 68714 0 din01[14]
rlabel metal1 1380 73746 1380 73746 0 din01[15]
rlabel metal1 1380 74154 1380 74154 0 din01[1]
rlabel metal2 1518 62067 1518 62067 0 din01[2]
rlabel metal1 1380 76330 1380 76330 0 din01[3]
rlabel metal1 1334 67626 1334 67626 0 din01[4]
rlabel metal1 1380 77010 1380 77010 0 din01[5]
rlabel metal1 1426 78098 1426 78098 0 din01[6]
rlabel metal1 1426 70890 1426 70890 0 din01[7]
rlabel metal1 1426 75242 1426 75242 0 din01[8]
rlabel metal1 1426 78506 1426 78506 0 din01[9]
rlabel metal4 23460 9118 23460 9118 0 net1
rlabel metal1 2208 70482 2208 70482 0 net10
rlabel metal1 100740 67286 100740 67286 0 net100
rlabel metal3 102279 85060 102279 85060 0 net101
rlabel metal1 104236 78506 104236 78506 0 net102
rlabel metal3 102279 25060 102279 25060 0 net103
rlabel metal4 86174 123835 86174 123835 0 net104
rlabel metal1 105294 78472 105294 78472 0 net105
rlabel metal4 86174 63983 86174 63983 0 net106
rlabel metal2 91586 67728 91586 67728 0 net107
rlabel metal4 87342 123767 87342 123767 0 net108
rlabel metal1 104650 85102 104650 85102 0 net109
rlabel metal2 8418 94095 8418 94095 0 net11
rlabel metal1 104190 78982 104190 78982 0 net110
rlabel metal2 91034 67065 91034 67065 0 net111
rlabel metal1 90160 66606 90160 66606 0 net112
rlabel metal1 104144 44302 104144 44302 0 net113
rlabel metal1 18492 66674 18492 66674 0 net114
rlabel metal3 102279 59738 102279 59738 0 net115
rlabel metal3 102279 119738 102279 119738 0 net116
rlabel metal4 90846 69854 90846 69854 0 net117
rlabel metal1 92138 66130 92138 66130 0 net118
rlabel metal2 105110 43894 105110 43894 0 net119
rlabel metal2 8418 95897 8418 95897 0 net12
rlabel metal2 8418 96985 8418 96985 0 net13
rlabel metal2 8418 98515 8418 98515 0 net14
rlabel metal2 8418 99603 8418 99603 0 net15
rlabel metal2 8418 101405 8418 101405 0 net16
rlabel metal2 9522 15699 9522 15699 0 net17
rlabel metal2 5566 75803 5566 75803 0 net18
rlabel metal4 25806 9934 25806 9934 0 net19
rlabel via3 24771 8228 24771 8228 0 net2
rlabel metal4 37486 9934 37486 9934 0 net20
rlabel metal4 38654 9934 38654 9934 0 net21
rlabel metal1 40020 2618 40020 2618 0 net22
rlabel metal4 40990 9934 40990 9934 0 net23
rlabel metal4 42158 9934 42158 9934 0 net24
rlabel metal3 43401 8228 43401 8228 0 net25
rlabel metal4 26956 9118 26956 9118 0 net26
rlabel metal3 28359 8228 28359 8228 0 net27
rlabel metal4 29310 9934 29310 9934 0 net28
rlabel metal4 30478 9934 30478 9934 0 net29
rlabel metal2 5566 34323 5566 34323 0 net3
rlabel via3 31717 8228 31717 8228 0 net30
rlabel metal4 32814 9934 32814 9934 0 net31
rlabel metal4 33982 9934 33982 9934 0 net32
rlabel metal1 35512 2618 35512 2618 0 net33
rlabel metal4 36318 9934 36318 9934 0 net34
rlabel metal1 1794 68170 1794 68170 0 net35
rlabel metal1 1794 69802 1794 69802 0 net36
rlabel metal2 1886 70686 1886 70686 0 net37
rlabel metal1 1794 72522 1794 72522 0 net38
rlabel metal1 1794 73202 1794 73202 0 net39
rlabel metal2 9522 35707 9522 35707 0 net4
rlabel metal1 1794 68714 1794 68714 0 net40
rlabel metal1 1748 73610 1748 73610 0 net41
rlabel metal2 1886 72896 1886 72896 0 net42
rlabel metal2 1886 63376 1886 63376 0 net43
rlabel metal1 1794 76330 1794 76330 0 net44
rlabel metal1 1978 67898 1978 67898 0 net45
rlabel metal1 1794 76874 1794 76874 0 net46
rlabel metal1 1794 77962 1794 77962 0 net47
rlabel metal1 1794 70958 1794 70958 0 net48
rlabel metal1 1794 75242 1794 75242 0 net49
rlabel metal1 1610 37128 1610 37128 0 net5
rlabel metal1 1794 78506 1794 78506 0 net50
rlabel metal1 106674 44846 106674 44846 0 net51
rlabel metal1 2622 63002 2622 63002 0 net52
rlabel via2 87998 66453 87998 66453 0 net53
rlabel metal2 85606 65688 85606 65688 0 net54
rlabel metal2 91218 65790 91218 65790 0 net55
rlabel metal1 91310 66538 91310 66538 0 net56
rlabel metal2 95910 68034 95910 68034 0 net57
rlabel metal1 93242 66742 93242 66742 0 net58
rlabel metal1 1702 64430 1702 64430 0 net59
rlabel via2 8418 38437 8418 38437 0 net6
rlabel metal1 2300 63478 2300 63478 0 net60
rlabel metal1 1702 65042 1702 65042 0 net61
rlabel metal1 1702 66130 1702 66130 0 net62
rlabel metal1 1702 67218 1702 67218 0 net63
rlabel metal1 1702 65518 1702 65518 0 net64
rlabel metal1 87584 67014 87584 67014 0 net65
rlabel via2 84686 66589 84686 66589 0 net66
rlabel metal2 88642 68000 88642 68000 0 net67
rlabel metal2 62238 126174 62238 126174 0 net68
rlabel metal2 59754 126208 59754 126208 0 net69
rlabel metal2 5566 39899 5566 39899 0 net7
rlabel metal1 58742 126446 58742 126446 0 net70
rlabel via2 44482 67133 44482 67133 0 net71
rlabel metal2 8050 96475 8050 96475 0 net72
rlabel metal2 45126 126174 45126 126174 0 net73
rlabel metal2 40986 126106 40986 126106 0 net74
rlabel metal2 41446 126140 41446 126140 0 net75
rlabel metal2 37674 126072 37674 126072 0 net76
rlabel metal1 77602 126378 77602 126378 0 net77
rlabel metal2 71806 126038 71806 126038 0 net78
rlabel metal2 70886 126004 70886 126004 0 net79
rlabel metal2 5566 41497 5566 41497 0 net8
rlabel metal2 67114 126072 67114 126072 0 net80
rlabel metal2 66010 126106 66010 126106 0 net81
rlabel metal2 64354 126140 64354 126140 0 net82
rlabel metal1 36340 126378 36340 126378 0 net83
rlabel metal1 44574 67184 44574 67184 0 net84
rlabel metal1 79488 67014 79488 67014 0 net85
rlabel metal4 90846 9934 90846 9934 0 net86
rlabel metal1 104972 56882 104972 56882 0 net87
rlabel metal1 104788 56406 104788 56406 0 net88
rlabel metal1 104420 56338 104420 56338 0 net89
rlabel metal1 1748 61846 1748 61846 0 net9
rlabel metal1 104696 37298 104696 37298 0 net90
rlabel metal1 104144 55386 104144 55386 0 net91
rlabel metal1 104420 57562 104420 57562 0 net92
rlabel metal4 90559 69786 90559 69786 0 net93
rlabel metal3 102279 22232 102279 22232 0 net94
rlabel metal1 104098 57494 104098 57494 0 net95
rlabel metal3 102279 82232 102279 82232 0 net96
rlabel metal2 99222 67524 99222 67524 0 net97
rlabel metal3 102026 23360 102026 23360 0 net98
rlabel metal3 102026 83360 102026 83360 0 net99
rlabel metal2 108514 51221 108514 51221 0 rst
rlabel metal3 751 62628 751 62628 0 sine_out[0]
rlabel metal2 108514 64141 108514 64141 0 sine_out[10]
rlabel metal2 108514 69581 108514 69581 0 sine_out[11]
rlabel via2 108514 66011 108514 66011 0 sine_out[12]
rlabel via2 108514 65365 108514 65365 0 sine_out[13]
rlabel via2 108514 68085 108514 68085 0 sine_out[14]
rlabel metal2 108514 67609 108514 67609 0 sine_out[15]
rlabel metal3 751 63988 751 63988 0 sine_out[1]
rlabel metal3 751 63308 751 63308 0 sine_out[2]
rlabel metal3 1050 64668 1050 64668 0 sine_out[3]
rlabel metal3 751 66028 751 66028 0 sine_out[4]
rlabel metal3 751 66708 751 66708 0 sine_out[5]
rlabel metal3 751 65348 751 65348 0 sine_out[6]
rlabel metal2 108514 64787 108514 64787 0 sine_out[7]
rlabel metal2 108514 66861 108514 66861 0 sine_out[8]
rlabel metal2 108514 68697 108514 68697 0 sine_out[9]
rlabel metal4 36107 63983 36107 63983 0 sine_out_temp0\[0\]
rlabel metal2 71898 65535 71898 65535 0 sine_out_temp0\[10\]
rlabel metal2 67574 66895 67574 66895 0 sine_out_temp0\[11\]
rlabel metal4 66059 63983 66059 63983 0 sine_out_temp0\[12\]
rlabel metal4 68555 63915 68555 63915 0 sine_out_temp0\[13\]
rlabel metal4 71051 63983 71051 63983 0 sine_out_temp0\[14\]
rlabel metal4 73547 63983 73547 63983 0 sine_out_temp0\[15\]
rlabel metal4 38603 63915 38603 63915 0 sine_out_temp0\[1\]
rlabel metal4 41099 63983 41099 63983 0 sine_out_temp0\[2\]
rlabel metal4 43595 63983 43595 63983 0 sine_out_temp0\[3\]
rlabel metal2 45770 66725 45770 66725 0 sine_out_temp0\[4\]
rlabel metal3 48047 64124 48047 64124 0 sine_out_temp0\[5\]
rlabel metal4 51071 64260 51071 64260 0 sine_out_temp0\[6\]
rlabel metal4 53579 63983 53579 63983 0 sine_out_temp0\[7\]
rlabel metal4 56075 63915 56075 63915 0 sine_out_temp0\[8\]
rlabel metal4 58571 63847 58571 63847 0 sine_out_temp0\[9\]
rlabel metal4 36107 123971 36107 123971 0 sine_out_temp1\[0\]
rlabel metal4 61088 123903 61088 123903 0 sine_out_temp1\[10\]
rlabel metal2 64446 125783 64446 125783 0 sine_out_temp1\[11\]
rlabel metal4 66059 123971 66059 123971 0 sine_out_temp1\[12\]
rlabel metal4 68555 123971 68555 123971 0 sine_out_temp1\[13\]
rlabel metal4 71051 123971 71051 123971 0 sine_out_temp1\[14\]
rlabel via2 77326 126395 77326 126395 0 sine_out_temp1\[15\]
rlabel metal4 38603 123971 38603 123971 0 sine_out_temp1\[1\]
rlabel metal4 41099 123971 41099 123971 0 sine_out_temp1\[2\]
rlabel metal4 43595 123903 43595 123903 0 sine_out_temp1\[3\]
rlabel metal2 45218 126191 45218 126191 0 sine_out_temp1\[4\]
rlabel metal4 48576 123971 48576 123971 0 sine_out_temp1\[5\]
rlabel metal4 51083 123903 51083 123903 0 sine_out_temp1\[6\]
rlabel metal2 56810 126191 56810 126191 0 sine_out_temp1\[7\]
rlabel metal4 56075 123903 56075 123903 0 sine_out_temp1\[8\]
rlabel metal4 58571 123903 58571 123903 0 sine_out_temp1\[9\]
rlabel metal1 91586 67728 91586 67728 0 tcout\[0\]
rlabel metal1 104650 78608 104650 78608 0 tcout\[1\]
rlabel metal2 90666 67932 90666 67932 0 tcout\[2\]
rlabel metal1 96968 67354 96968 67354 0 tcout\[3\]
rlabel metal2 93794 67354 93794 67354 0 tcout\[4\]
rlabel metal1 96738 66606 96738 66606 0 tcout\[5\]
rlabel metal1 104374 42194 104374 42194 0 tcout\[6\]
rlabel metal2 94990 67320 94990 67320 0 tcout\[7\]
rlabel metal2 77602 66368 77602 66368 0 tcout\[8\]
<< properties >>
string FIXED_BBOX 0 0 110000 130000
<< end >>
