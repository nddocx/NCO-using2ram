logic [0:255] [15:0]  sine_table0 = { 
16'h0000,
16'h0192,
16'h0324,
16'h04b6,
16'h0648,
16'h07d9,
16'h096a,
16'h0afb,
16'h0c8c,
16'h0e1c,
16'h0fab,
16'h113a,
16'h12c8,
16'h1455,
16'h15e2,
16'h176e,
16'h18f9,
16'h1a82,
16'h1c0b,
16'h1d93,
16'h1f1a,
16'h209f,
16'h2223,
16'h23a6,
16'h2528,
16'h26a8,
16'h2826,
16'h29a3,
16'h2b1f,
16'h2c99,
16'h2e11,
16'h2f87,
16'h30fb,
16'h326e,
16'h33df,
16'h354d,
16'h36ba,
16'h3824,
16'h398c,
16'h3af2,
16'h3c56,
16'h3db8,
16'h3f17,
16'h4073,
16'h41ce,
16'h4325,
16'h447a,
16'h45cd,
16'h471c,
16'h4869,
16'h49b4,
16'h4afb,
16'h4c3f,
16'h4d81,
16'h4ebf,
16'h4ffb,
16'h5133,
16'h5268,
16'h539b,
16'h54c9,
16'h55f5,
16'h571d,
16'h5842,
16'h5964,
16'h5a82,
16'h5b9c,
16'h5cb3,
16'h5dc7,
16'h5ed7,
16'h5fe3,
16'h60eb,
16'h61f0,
16'h62f1,
16'h63ee,
16'h64e8,
16'h65dd,
16'h66cf,
16'h67bc,
16'h68a6,
16'h698b,
16'h6a6d,
16'h6b4a,
16'h6c23,
16'h6cf8,
16'h6dc9,
16'h6e96,
16'h6f5e,
16'h7022,
16'h70e2,
16'h719d,
16'h7254,
16'h7307,
16'h73b5,
16'h745f,
16'h7504,
16'h75a5,
16'h7641,
16'h76d8,
16'h776b,
16'h77fa,
16'h7884,
16'h7909,
16'h7989,
16'h7a05,
16'h7a7c,
16'h7aee,
16'h7b5c,
16'h7bc5,
16'h7c29,
16'h7c88,
16'h7ce3,
16'h7d39,
16'h7d89,
16'h7dd5,
16'h7e1d,
16'h7e5f,
16'h7e9c,
16'h7ed5,
16'h7f09,
16'h7f37,
16'h7f61,
16'h7f86,
16'h7fa6,
16'h7fc1,
16'h7fd8,
16'h7fe9,
16'h7ff5,
16'h7ffd,
16'h7fff,
16'h7ffd,
16'h7ff5,
16'h7fe9,
16'h7fd8,
16'h7fc1,
16'h7fa6,
16'h7f86,
16'h7f61,
16'h7f37,
16'h7f09,
16'h7ed5,
16'h7e9c,
16'h7e5f,
16'h7e1d,
16'h7dd5,
16'h7d89,
16'h7d39,
16'h7ce3,
16'h7c88,
16'h7c29,
16'h7bc5,
16'h7b5c,
16'h7aee,
16'h7a7c,
16'h7a05,
16'h7989,
16'h7909,
16'h7884,
16'h77fa,
16'h776b,
16'h76d8,
16'h7641,
16'h75a5,
16'h7504,
16'h745f,
16'h73b5,
16'h7307,
16'h7254,
16'h719d,
16'h70e2,
16'h7022,
16'h6f5e,
16'h6e96,
16'h6dc9,
16'h6cf8,
16'h6c23,
16'h6b4a,
16'h6a6d,
16'h698b,
16'h68a6,
16'h67bc,
16'h66cf,
16'h65dd,
16'h64e8,
16'h63ee,
16'h62f1,
16'h61f0,
16'h60eb,
16'h5fe3,
16'h5ed7,
16'h5dc7,
16'h5cb3,
16'h5b9c,
16'h5a82,
16'h5964,
16'h5842,
16'h571d,
16'h55f5,
16'h54c9,
16'h539b,
16'h5268,
16'h5133,
16'h4ffb,
16'h4ebf,
16'h4d81,
16'h4c3f,
16'h4afb,
16'h49b4,
16'h4869,
16'h471c,
16'h45cd,
16'h447a,
16'h4325,
16'h41ce,
16'h4073,
16'h3f17,
16'h3db8,
16'h3c56,
16'h3af2,
16'h398c,
16'h3824,
16'h36ba,
16'h354d,
16'h33df,
16'h326e,
16'h30fb,
16'h2f87,
16'h2e11,
16'h2c99,
16'h2b1f,
16'h29a3,
16'h2826,
16'h26a8,
16'h2528,
16'h23a6,
16'h2223,
16'h209f,
16'h1f1a,
16'h1d93,
16'h1c0b,
16'h1a82,
16'h18f9,
16'h176e,
16'h15e2,
16'h1455,
16'h12c8,
16'h113a,
16'h0fab,
16'h0e1c,
16'h0c8c,
16'h0afb,
16'h096a,
16'h07d9,
16'h0648,
16'h04b6,
16'h0324,
16'h0192
};
