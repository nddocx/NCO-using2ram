magic
tech sky130A
magscale 1 2
timestamp 1741114801
<< viali >>
rect 47593 136221 47627 136255
rect 47961 136221 47995 136255
rect 53757 136221 53791 136255
rect 53941 136221 53975 136255
rect 38209 136153 38243 136187
rect 40693 136153 40727 136187
rect 42993 136153 43027 136187
rect 45293 136153 45327 136187
rect 47777 136153 47811 136187
rect 53573 136153 53607 136187
rect 55781 136153 55815 136187
rect 58173 136153 58207 136187
rect 60657 136153 60691 136187
rect 63141 136153 63175 136187
rect 64981 136153 65015 136187
rect 67557 136153 67591 136187
rect 69765 136153 69799 136187
rect 72157 136153 72191 136187
rect 74181 136153 74215 136187
rect 36093 136085 36127 136119
rect 38117 136085 38151 136119
rect 38393 136085 38427 136119
rect 40601 136085 40635 136119
rect 40877 136085 40911 136119
rect 42901 136085 42935 136119
rect 43177 136085 43211 136119
rect 45201 136085 45235 136119
rect 45477 136085 45511 136119
rect 55873 136085 55907 136119
rect 56149 136085 56183 136119
rect 58265 136085 58299 136119
rect 58541 136085 58575 136119
rect 60749 136085 60783 136119
rect 61025 136085 61059 136119
rect 63233 136085 63267 136119
rect 63509 136085 63543 136119
rect 65073 136085 65107 136119
rect 65349 136085 65383 136119
rect 67649 136085 67683 136119
rect 67925 136085 67959 136119
rect 69857 136085 69891 136119
rect 70133 136085 70167 136119
rect 72249 136085 72283 136119
rect 72525 136085 72559 136119
rect 74273 136085 74307 136119
rect 74549 136085 74583 136119
rect 86233 136085 86267 136119
rect 87337 136085 87371 136119
rect 95985 136085 96019 136119
rect 104357 129829 104391 129863
rect 1593 111333 1627 111367
rect 1409 111197 1443 111231
rect 1685 111197 1719 111231
rect 1409 109633 1443 109667
rect 1685 109633 1719 109667
rect 1593 109497 1627 109531
rect 1409 108545 1443 108579
rect 1685 108545 1719 108579
rect 1593 108409 1627 108443
rect 1593 106981 1627 107015
rect 1409 106845 1443 106879
rect 1685 106845 1719 106879
rect 1593 105893 1627 105927
rect 1409 105757 1443 105791
rect 1685 105757 1719 105791
rect 1409 104193 1443 104227
rect 1685 104193 1719 104227
rect 1593 104057 1627 104091
rect 104357 95285 104391 95319
rect 104357 93857 104391 93891
rect 104357 92565 104391 92599
rect 104357 91137 104391 91171
rect 105645 90933 105679 90967
rect 106197 90933 106231 90967
rect 104357 90389 104391 90423
rect 1501 88961 1535 88995
rect 1961 88961 1995 88995
rect 1685 88825 1719 88859
rect 1869 88825 1903 88859
rect 1501 87873 1535 87907
rect 1961 87873 1995 87907
rect 1685 87737 1719 87771
rect 1869 87737 1903 87771
rect 1501 87193 1535 87227
rect 1961 87193 1995 87227
rect 1593 87125 1627 87159
rect 1869 87125 1903 87159
rect 1501 86785 1535 86819
rect 1961 86785 1995 86819
rect 1685 86649 1719 86683
rect 1869 86649 1903 86683
rect 1409 86173 1443 86207
rect 1685 86173 1719 86207
rect 1593 86037 1627 86071
rect 1501 85017 1535 85051
rect 1961 85017 1995 85051
rect 1593 84949 1627 84983
rect 1777 84949 1811 84983
rect 1501 84609 1535 84643
rect 1961 84609 1995 84643
rect 1685 84473 1719 84507
rect 1777 84473 1811 84507
rect 1501 83929 1535 83963
rect 1685 83929 1719 83963
rect 1869 83929 1903 83963
rect 1961 83861 1995 83895
rect 1501 83521 1535 83555
rect 1961 83521 1995 83555
rect 1593 83317 1627 83351
rect 1869 83317 1903 83351
rect 1501 82433 1535 82467
rect 1961 82433 1995 82467
rect 1593 82229 1627 82263
rect 1869 82229 1903 82263
rect 1501 81753 1535 81787
rect 1961 81753 1995 81787
rect 1593 81685 1627 81719
rect 1869 81685 1903 81719
rect 1501 81345 1535 81379
rect 1961 81345 1995 81379
rect 1593 81141 1627 81175
rect 1777 81141 1811 81175
rect 1409 80733 1443 80767
rect 1685 80733 1719 80767
rect 2421 80597 2455 80631
rect 1409 80325 1443 80359
rect 1501 79577 1535 79611
rect 1685 79577 1719 79611
rect 1869 79577 1903 79611
rect 1961 79509 1995 79543
rect 1501 79169 1535 79203
rect 1961 79169 1995 79203
rect 108313 79169 108347 79203
rect 1685 79033 1719 79067
rect 1869 79033 1903 79067
rect 108129 78965 108163 78999
rect 108497 78965 108531 78999
rect 108313 78557 108347 78591
rect 1501 78489 1535 78523
rect 1685 78489 1719 78523
rect 1869 78489 1903 78523
rect 1961 78421 1995 78455
rect 108129 78421 108163 78455
rect 108497 78421 108531 78455
rect 1501 78081 1535 78115
rect 1961 78081 1995 78115
rect 108313 78081 108347 78115
rect 1685 77945 1719 77979
rect 1869 77945 1903 77979
rect 108129 77877 108163 77911
rect 108497 77877 108531 77911
rect 21833 77673 21867 77707
rect 27629 77673 27663 77707
rect 28181 77673 28215 77707
rect 29561 77673 29595 77707
rect 30481 77673 30515 77707
rect 30757 77673 30791 77707
rect 31677 77673 31711 77707
rect 32505 77673 32539 77707
rect 33701 77673 33735 77707
rect 33977 77673 34011 77707
rect 34713 77673 34747 77707
rect 34897 77673 34931 77707
rect 35817 77673 35851 77707
rect 70225 77673 70259 77707
rect 70409 77673 70443 77707
rect 70961 77673 70995 77707
rect 71973 77673 72007 77707
rect 74457 77673 74491 77707
rect 76665 77673 76699 77707
rect 78229 77673 78263 77707
rect 79241 77673 79275 77707
rect 80069 77673 80103 77707
rect 19809 77605 19843 77639
rect 24685 77605 24719 77639
rect 24869 77605 24903 77639
rect 25053 77605 25087 77639
rect 27261 77605 27295 77639
rect 38669 77605 38703 77639
rect 39681 77605 39715 77639
rect 39865 77605 39899 77639
rect 40877 77605 40911 77639
rect 41245 77605 41279 77639
rect 42165 77605 42199 77639
rect 43729 77605 43763 77639
rect 62497 77605 62531 77639
rect 63785 77605 63819 77639
rect 63969 77605 64003 77639
rect 67649 77605 67683 77639
rect 68937 77605 68971 77639
rect 69121 77605 69155 77639
rect 70501 77605 70535 77639
rect 71145 77605 71179 77639
rect 73445 77605 73479 77639
rect 77769 77605 77803 77639
rect 79885 77605 79919 77639
rect 80897 77605 80931 77639
rect 87337 77605 87371 77639
rect 90557 77605 90591 77639
rect 90741 77605 90775 77639
rect 93133 77605 93167 77639
rect 95709 77605 95743 77639
rect 21557 77537 21591 77571
rect 22293 77537 22327 77571
rect 22477 77537 22511 77571
rect 22753 77537 22787 77571
rect 31217 77537 31251 77571
rect 31401 77537 31435 77571
rect 32137 77537 32171 77571
rect 33149 77537 33183 77571
rect 33241 77537 33275 77571
rect 34161 77537 34195 77571
rect 35449 77537 35483 77571
rect 36093 77537 36127 77571
rect 37841 77537 37875 77571
rect 38485 77537 38519 77571
rect 40509 77537 40543 77571
rect 41153 77537 41187 77571
rect 43085 77537 43119 77571
rect 43821 77537 43855 77571
rect 61025 77537 61059 77571
rect 61853 77537 61887 77571
rect 63141 77537 63175 77571
rect 64061 77537 64095 77571
rect 65717 77537 65751 77571
rect 66637 77537 66671 77571
rect 68293 77537 68327 77571
rect 68477 77537 68511 77571
rect 69581 77537 69615 77571
rect 69765 77537 69799 77571
rect 71329 77537 71363 77571
rect 72065 77537 72099 77571
rect 73813 77537 73847 77571
rect 73997 77537 74031 77571
rect 76113 77537 76147 77571
rect 76205 77537 76239 77571
rect 78689 77537 78723 77571
rect 78781 77537 78815 77571
rect 79701 77537 79735 77571
rect 80253 77537 80287 77571
rect 80437 77537 80471 77571
rect 81633 77537 81667 77571
rect 85681 77537 85715 77571
rect 86233 77537 86267 77571
rect 86509 77537 86543 77571
rect 93961 77537 93995 77571
rect 95801 77537 95835 77571
rect 26801 77469 26835 77503
rect 27077 77469 27111 77503
rect 31125 77469 31159 77503
rect 31769 77469 31803 77503
rect 35265 77469 35299 77503
rect 35357 77469 35391 77503
rect 35909 77469 35943 77503
rect 36369 77469 36403 77503
rect 37013 77469 37047 77503
rect 37657 77469 37691 77503
rect 38209 77469 38243 77503
rect 40785 77469 40819 77503
rect 60565 77469 60599 77503
rect 61117 77469 61151 77503
rect 62773 77469 62807 77503
rect 63325 77469 63359 77503
rect 65349 77469 65383 77503
rect 65901 77469 65935 77503
rect 67925 77469 67959 77503
rect 68569 77469 68603 77503
rect 74641 77469 74675 77503
rect 75469 77469 75503 77503
rect 78873 77469 78907 77503
rect 80529 77469 80563 77503
rect 83381 77469 83415 77503
rect 83841 77469 83875 77503
rect 85957 77469 85991 77503
rect 86601 77469 86635 77503
rect 88809 77469 88843 77503
rect 91385 77469 91419 77503
rect 21281 77401 21315 77435
rect 26525 77401 26559 77435
rect 40233 77401 40267 77435
rect 42809 77401 42843 77435
rect 43361 77401 43395 77435
rect 60749 77401 60783 77435
rect 61209 77401 61243 77435
rect 63417 77401 63451 77435
rect 65165 77401 65199 77435
rect 65993 77401 66027 77435
rect 66545 77401 66579 77435
rect 71605 77401 71639 77435
rect 73537 77401 73571 77435
rect 74089 77401 74123 77435
rect 75009 77401 75043 77435
rect 75193 77401 75227 77435
rect 75377 77401 75411 77435
rect 75745 77401 75779 77435
rect 78045 77401 78079 77435
rect 83105 77401 83139 77435
rect 86969 77401 87003 77435
rect 87153 77401 87187 77435
rect 89085 77401 89119 77435
rect 91661 77401 91695 77435
rect 94237 77401 94271 77435
rect 16129 77333 16163 77367
rect 19625 77333 19659 77367
rect 24225 77333 24259 77367
rect 24409 77333 24443 77367
rect 27445 77333 27479 77367
rect 32321 77333 32355 77367
rect 32689 77333 32723 77367
rect 33057 77333 33091 77367
rect 33609 77333 33643 77367
rect 37289 77333 37323 77367
rect 37749 77333 37783 77367
rect 38301 77333 38335 77367
rect 40325 77333 40359 77367
rect 42441 77333 42475 77367
rect 42901 77333 42935 77367
rect 43453 77333 43487 77367
rect 61577 77333 61611 77367
rect 61761 77333 61795 77367
rect 66361 77333 66395 77367
rect 69305 77333 69339 77367
rect 69857 77333 69891 77367
rect 71513 77333 71547 77367
rect 76297 77333 76331 77367
rect 83657 77333 83691 77367
rect 84025 77333 84059 77367
rect 84209 77333 84243 77367
rect 90925 77333 90959 77367
rect 93317 77333 93351 77367
rect 27629 77129 27663 77163
rect 75837 77129 75871 77163
rect 81541 77129 81575 77163
rect 83933 77129 83967 77163
rect 88625 77129 88659 77163
rect 88901 77129 88935 77163
rect 92029 77129 92063 77163
rect 30297 77061 30331 77095
rect 69213 77061 69247 77095
rect 75653 77061 75687 77095
rect 91753 77061 91787 77095
rect 1501 76993 1535 77027
rect 1961 76993 1995 77027
rect 26433 76993 26467 77027
rect 27721 76993 27755 77027
rect 27905 76993 27939 77027
rect 30389 76993 30423 77027
rect 81633 76993 81667 77027
rect 84025 76993 84059 77027
rect 84117 76993 84151 77027
rect 85957 76993 85991 77027
rect 86601 76993 86635 77027
rect 86785 76993 86819 77027
rect 86877 76993 86911 77027
rect 89085 76993 89119 77027
rect 89453 76993 89487 77027
rect 91661 76993 91695 77027
rect 108313 76993 108347 77027
rect 22753 76925 22787 76959
rect 24317 76925 24351 76959
rect 24593 76925 24627 76959
rect 26157 76925 26191 76959
rect 87153 76925 87187 76959
rect 89729 76925 89763 76959
rect 1685 76857 1719 76891
rect 1869 76857 1903 76891
rect 69397 76857 69431 76891
rect 91201 76857 91235 76891
rect 91385 76857 91419 76891
rect 108497 76857 108531 76891
rect 22845 76789 22879 76823
rect 24685 76789 24719 76823
rect 26525 76789 26559 76823
rect 26801 76789 26835 76823
rect 30573 76789 30607 76823
rect 81817 76789 81851 76823
rect 84301 76789 84335 76823
rect 85865 76789 85899 76823
rect 86141 76789 86175 76823
rect 86417 76789 86451 76823
rect 91477 76789 91511 76823
rect 21557 76585 21591 76619
rect 23489 76585 23523 76619
rect 23581 76585 23615 76619
rect 24961 76585 24995 76619
rect 31585 76585 31619 76619
rect 82829 76585 82863 76619
rect 85773 76585 85807 76619
rect 85957 76585 85991 76619
rect 88533 76585 88567 76619
rect 88993 76585 89027 76619
rect 89821 76585 89855 76619
rect 24685 76517 24719 76551
rect 31033 76517 31067 76551
rect 88165 76517 88199 76551
rect 21741 76449 21775 76483
rect 22017 76449 22051 76483
rect 83013 76449 83047 76483
rect 85129 76449 85163 76483
rect 86233 76449 86267 76483
rect 1593 76381 1627 76415
rect 1777 76381 1811 76415
rect 29101 76381 29135 76415
rect 29285 76381 29319 76415
rect 31125 76381 31159 76415
rect 31309 76381 31343 76415
rect 31677 76381 31711 76415
rect 31861 76381 31895 76415
rect 32413 76381 32447 76415
rect 82277 76381 82311 76415
rect 82369 76381 82403 76415
rect 82737 76381 82771 76415
rect 85681 76381 85715 76415
rect 88073 76381 88107 76415
rect 88441 76381 88475 76415
rect 89729 76381 89763 76415
rect 108313 76381 108347 76415
rect 29009 76313 29043 76347
rect 32321 76313 32355 76347
rect 82461 76313 82495 76347
rect 83289 76313 83323 76347
rect 86509 76313 86543 76347
rect 88809 76313 88843 76347
rect 1409 76245 1443 76279
rect 32597 76245 32631 76279
rect 84761 76245 84795 76279
rect 84945 76245 84979 76279
rect 87981 76245 88015 76279
rect 89177 76245 89211 76279
rect 90005 76245 90039 76279
rect 108497 76245 108531 76279
rect 1777 76041 1811 76075
rect 83105 76041 83139 76075
rect 83933 76041 83967 76075
rect 90097 76041 90131 76075
rect 108129 76041 108163 76075
rect 108497 76041 108531 76075
rect 82921 75973 82955 76007
rect 83749 75973 83783 76007
rect 86417 75973 86451 76007
rect 90281 75973 90315 76007
rect 1593 75905 1627 75939
rect 83657 75905 83691 75939
rect 84301 75905 84335 75939
rect 90005 75905 90039 75939
rect 90373 75905 90407 75939
rect 90833 75905 90867 75939
rect 108313 75905 108347 75939
rect 84209 75837 84243 75871
rect 84577 75837 84611 75871
rect 86693 75837 86727 75871
rect 86969 75837 87003 75871
rect 88901 75837 88935 75871
rect 86049 75769 86083 75803
rect 88441 75769 88475 75803
rect 88625 75769 88659 75803
rect 91017 75769 91051 75803
rect 91201 75769 91235 75803
rect 1409 75701 1443 75735
rect 86325 75701 86359 75735
rect 90281 75701 90315 75735
rect 90557 75701 90591 75735
rect 86785 75497 86819 75531
rect 90649 75497 90683 75531
rect 86325 75429 86359 75463
rect 82737 75361 82771 75395
rect 85589 75361 85623 75395
rect 1593 75293 1627 75327
rect 82185 75293 82219 75327
rect 82461 75293 82495 75327
rect 85497 75293 85531 75327
rect 86233 75293 86267 75327
rect 86601 75293 86635 75327
rect 108313 75293 108347 75327
rect 81817 75225 81851 75259
rect 90833 75225 90867 75259
rect 108129 75225 108163 75259
rect 1409 75157 1443 75191
rect 1777 75157 1811 75191
rect 82093 75157 82127 75191
rect 82277 75157 82311 75191
rect 84209 75157 84243 75191
rect 84393 75157 84427 75191
rect 86969 75157 87003 75191
rect 90465 75157 90499 75191
rect 90633 75157 90667 75191
rect 108497 75157 108531 75191
rect 82553 74953 82587 74987
rect 1409 74341 1443 74375
rect 1593 74205 1627 74239
rect 1777 74205 1811 74239
rect 108129 74205 108163 74239
rect 108313 74205 108347 74239
rect 108497 74069 108531 74103
rect 1593 73729 1627 73763
rect 1777 73729 1811 73763
rect 108313 73729 108347 73763
rect 1409 73593 1443 73627
rect 108129 73525 108163 73559
rect 108497 73525 108531 73559
rect 1777 73321 1811 73355
rect 108129 73321 108163 73355
rect 90097 73253 90131 73287
rect 1593 73117 1627 73151
rect 90097 73117 90131 73151
rect 90281 73117 90315 73151
rect 108313 73117 108347 73151
rect 1409 72981 1443 73015
rect 108497 72981 108531 73015
rect 44649 72709 44683 72743
rect 75101 72709 75135 72743
rect 1501 72641 1535 72675
rect 1961 72641 1995 72675
rect 44189 72641 44223 72675
rect 46581 72641 46615 72675
rect 46397 72573 46431 72607
rect 73629 72573 73663 72607
rect 75377 72573 75411 72607
rect 1685 72505 1719 72539
rect 1869 72505 1903 72539
rect 46765 72437 46799 72471
rect 73445 72437 73479 72471
rect 44649 72233 44683 72267
rect 74181 72233 74215 72267
rect 74089 72029 74123 72063
rect 90741 72029 90775 72063
rect 91569 72029 91603 72063
rect 55873 71961 55907 71995
rect 56057 71961 56091 71995
rect 57805 71961 57839 71995
rect 91753 71961 91787 71995
rect 91937 71961 91971 71995
rect 92489 71961 92523 71995
rect 92673 71961 92707 71995
rect 92857 71961 92891 71995
rect 57989 71893 58023 71927
rect 74365 71893 74399 71927
rect 90557 71893 90591 71927
rect 91845 71893 91879 71927
rect 92121 71893 92155 71927
rect 90741 71689 90775 71723
rect 90925 71553 90959 71587
rect 91845 71553 91879 71587
rect 92029 71349 92063 71383
rect 92305 71349 92339 71383
rect 90465 71145 90499 71179
rect 77769 71009 77803 71043
rect 78137 71009 78171 71043
rect 88717 71009 88751 71043
rect 90557 71009 90591 71043
rect 77585 70941 77619 70975
rect 87889 70941 87923 70975
rect 88993 70873 89027 70907
rect 87981 70805 88015 70839
rect 78045 70601 78079 70635
rect 77769 70465 77803 70499
rect 77401 70397 77435 70431
rect 77861 70397 77895 70431
rect 89085 69173 89119 69207
rect 90741 68901 90775 68935
rect 89269 68833 89303 68867
rect 88993 68765 89027 68799
rect 89545 68765 89579 68799
rect 89821 68765 89855 68799
rect 90097 68765 90131 68799
rect 90189 68765 90223 68799
rect 90557 68765 90591 68799
rect 92213 68765 92247 68799
rect 92397 68765 92431 68799
rect 88717 68697 88751 68731
rect 90465 68629 90499 68663
rect 92305 68629 92339 68663
rect 86601 68289 86635 68323
rect 88993 68289 89027 68323
rect 86693 68085 86727 68119
rect 89085 68085 89119 68119
rect 90557 67881 90591 67915
rect 107945 67881 107979 67915
rect 108313 67881 108347 67915
rect 88809 67813 88843 67847
rect 92581 67813 92615 67847
rect 92857 67813 92891 67847
rect 86233 67677 86267 67711
rect 88625 67677 88659 67711
rect 89729 67677 89763 67711
rect 90189 67677 90223 67711
rect 90373 67677 90407 67711
rect 90925 67677 90959 67711
rect 91109 67677 91143 67711
rect 92397 67677 92431 67711
rect 108221 67677 108255 67711
rect 108497 67677 108531 67711
rect 86325 67609 86359 67643
rect 89453 67609 89487 67643
rect 89637 67609 89671 67643
rect 90097 67609 90131 67643
rect 89913 67541 89947 67575
rect 91017 67541 91051 67575
rect 88625 67337 88659 67371
rect 88809 67337 88843 67371
rect 91753 67337 91787 67371
rect 90281 67269 90315 67303
rect 83933 67201 83967 67235
rect 84393 67201 84427 67235
rect 88441 67201 88475 67235
rect 89361 67201 89395 67235
rect 89637 67201 89671 67235
rect 90005 67201 90039 67235
rect 88165 67133 88199 67167
rect 89453 67133 89487 67167
rect 83841 66997 83875 67031
rect 84485 66997 84519 67031
rect 86693 66997 86727 67031
rect 88993 66997 89027 67031
rect 89821 66997 89855 67031
rect 91937 66997 91971 67031
rect 83841 66793 83875 66827
rect 85773 66793 85807 66827
rect 91017 66793 91051 66827
rect 90005 66725 90039 66759
rect 90557 66725 90591 66759
rect 84025 66657 84059 66691
rect 87337 66657 87371 66691
rect 89177 66657 89211 66691
rect 89637 66589 89671 66623
rect 90189 66589 90223 66623
rect 90281 66589 90315 66623
rect 91017 66589 91051 66623
rect 91201 66589 91235 66623
rect 91569 66589 91603 66623
rect 91753 66589 91787 66623
rect 84301 66521 84335 66555
rect 88901 66521 88935 66555
rect 89361 66521 89395 66555
rect 90557 66521 90591 66555
rect 90741 66521 90775 66555
rect 90925 66521 90959 66555
rect 87429 66453 87463 66487
rect 89453 66453 89487 66487
rect 89821 66453 89855 66487
rect 90373 66453 90407 66487
rect 91385 66453 91419 66487
rect 91937 66453 91971 66487
rect 85221 66249 85255 66283
rect 88441 66249 88475 66283
rect 89269 66249 89303 66283
rect 91017 66249 91051 66283
rect 36093 66181 36127 66215
rect 38669 66181 38703 66215
rect 41153 66181 41187 66215
rect 43637 66181 43671 66215
rect 46121 66181 46155 66215
rect 48605 66181 48639 66215
rect 51089 66181 51123 66215
rect 53573 66181 53607 66215
rect 56149 66181 56183 66215
rect 58633 66181 58667 66215
rect 61117 66181 61151 66215
rect 63601 66181 63635 66215
rect 66085 66181 66119 66215
rect 68569 66181 68603 66215
rect 71053 66181 71087 66215
rect 73537 66181 73571 66215
rect 88073 66181 88107 66215
rect 88257 66181 88291 66215
rect 89545 66181 89579 66215
rect 90649 66181 90683 66215
rect 91553 66181 91587 66215
rect 91753 66181 91787 66215
rect 94329 66181 94363 66215
rect 94421 66181 94455 66215
rect 85681 66113 85715 66147
rect 87981 66113 88015 66147
rect 88349 66113 88383 66147
rect 89361 66113 89395 66147
rect 89729 66113 89763 66147
rect 89913 66113 89947 66147
rect 90373 66113 90407 66147
rect 90833 66113 90867 66147
rect 91201 66113 91235 66147
rect 91937 66113 91971 66147
rect 87705 66045 87739 66079
rect 88809 66045 88843 66079
rect 88993 66045 89027 66079
rect 89085 66045 89119 66079
rect 89453 66045 89487 66079
rect 90465 66045 90499 66079
rect 85405 65977 85439 66011
rect 88625 65977 88659 66011
rect 86233 65909 86267 65943
rect 90005 65909 90039 65943
rect 91385 65909 91419 65943
rect 91569 65909 91603 65943
rect 92029 65909 92063 65943
rect 92305 65909 92339 65943
rect 95893 65909 95927 65943
rect 96261 65909 96295 65943
rect 96537 65909 96571 65943
rect 7297 60673 7331 60707
rect 7481 60605 7515 60639
rect 6285 60265 6319 60299
rect 7573 60061 7607 60095
rect 104357 60061 104391 60095
rect 6929 59721 6963 59755
rect 7205 59653 7239 59687
rect 7573 41429 7607 41463
rect 7481 39797 7515 39831
rect 7573 38709 7607 38743
rect 7573 36601 7607 36635
rect 7481 35445 7515 35479
rect 7573 33881 7607 33915
rect 104357 25109 104391 25143
rect 104357 23817 104391 23851
rect 104357 22729 104391 22763
rect 7481 15317 7515 15351
rect 1593 14025 1627 14059
rect 1869 14025 1903 14059
rect 1501 13889 1535 13923
rect 1961 13889 1995 13923
rect 1593 13481 1627 13515
rect 1869 13481 1903 13515
rect 1501 13209 1535 13243
rect 1961 13209 1995 13243
rect 1685 12869 1719 12903
rect 1777 12869 1811 12903
rect 1501 12801 1535 12835
rect 1961 12801 1995 12835
rect 1593 11849 1627 11883
rect 1777 11849 1811 11883
rect 1501 11713 1535 11747
rect 1961 11713 1995 11747
rect 1593 11305 1627 11339
rect 1869 11305 1903 11339
rect 1501 11033 1535 11067
rect 1961 11033 1995 11067
rect 1593 10761 1627 10795
rect 1777 10761 1811 10795
rect 1501 10625 1535 10659
rect 1961 10625 1995 10659
rect 1501 9945 1535 9979
rect 1685 9945 1719 9979
rect 1869 9945 1903 9979
rect 1961 9877 1995 9911
rect 1501 8857 1535 8891
rect 1685 8857 1719 8891
rect 1869 8857 1903 8891
rect 1961 8789 1995 8823
rect 1961 8381 1995 8415
rect 2237 8381 2271 8415
rect 2421 8313 2455 8347
rect 1961 8041 1995 8075
rect 2145 7837 2179 7871
rect 1501 7769 1535 7803
rect 1685 7769 1719 7803
rect 1869 7769 1903 7803
rect 16129 7497 16163 7531
rect 23489 7497 23523 7531
rect 24685 7497 24719 7531
rect 25881 7497 25915 7531
rect 26985 7497 27019 7531
rect 28181 7497 28215 7531
rect 29561 7497 29595 7531
rect 30481 7497 30515 7531
rect 90557 7497 90591 7531
rect 90741 7497 90775 7531
rect 90925 7497 90959 7531
rect 1501 7361 1535 7395
rect 1961 7361 1995 7395
rect 1685 7225 1719 7259
rect 1869 7225 1903 7259
rect 1501 6273 1535 6307
rect 1961 6273 1995 6307
rect 1685 6137 1719 6171
rect 1869 6137 1903 6171
rect 1593 5865 1627 5899
rect 1777 5865 1811 5899
rect 1409 5661 1443 5695
rect 1869 5661 1903 5695
rect 1501 5185 1535 5219
rect 1961 5185 1995 5219
rect 1685 5049 1719 5083
rect 1869 5049 1903 5083
rect 31677 2601 31711 2635
rect 32965 2601 32999 2635
rect 34253 2601 34287 2635
rect 35541 2601 35575 2635
rect 36369 2601 36403 2635
rect 37473 2601 37507 2635
rect 38761 2601 38795 2635
rect 40049 2601 40083 2635
rect 41337 2601 41371 2635
rect 42165 2601 42199 2635
rect 43453 2601 43487 2635
rect 31861 2397 31895 2431
rect 33149 2397 33183 2431
rect 34437 2397 34471 2431
rect 35725 2397 35759 2431
rect 36185 2397 36219 2431
rect 37657 2397 37691 2431
rect 38945 2397 38979 2431
rect 40233 2397 40267 2431
rect 41521 2397 41555 2431
rect 41981 2397 42015 2431
rect 43269 2397 43303 2431
rect 31585 2261 31619 2295
rect 32873 2261 32907 2295
rect 34161 2261 34195 2295
rect 35449 2261 35483 2295
rect 36093 2261 36127 2295
rect 37381 2261 37415 2295
rect 38669 2261 38703 2295
rect 39957 2261 39991 2295
rect 41245 2261 41279 2295
rect 41889 2261 41923 2295
rect 43177 2261 43211 2295
<< metal1 >>
rect 1104 147450 108836 147472
rect 1104 147398 4214 147450
rect 4266 147398 4278 147450
rect 4330 147398 4342 147450
rect 4394 147398 4406 147450
rect 4458 147398 4470 147450
rect 4522 147398 34934 147450
rect 34986 147398 34998 147450
rect 35050 147398 35062 147450
rect 35114 147398 35126 147450
rect 35178 147398 35190 147450
rect 35242 147398 65654 147450
rect 65706 147398 65718 147450
rect 65770 147398 65782 147450
rect 65834 147398 65846 147450
rect 65898 147398 65910 147450
rect 65962 147398 96374 147450
rect 96426 147398 96438 147450
rect 96490 147398 96502 147450
rect 96554 147398 96566 147450
rect 96618 147398 96630 147450
rect 96682 147398 108836 147450
rect 1104 147376 108836 147398
rect 1104 146906 108836 146928
rect 1104 146854 4874 146906
rect 4926 146854 4938 146906
rect 4990 146854 5002 146906
rect 5054 146854 5066 146906
rect 5118 146854 5130 146906
rect 5182 146854 35594 146906
rect 35646 146854 35658 146906
rect 35710 146854 35722 146906
rect 35774 146854 35786 146906
rect 35838 146854 35850 146906
rect 35902 146854 66314 146906
rect 66366 146854 66378 146906
rect 66430 146854 66442 146906
rect 66494 146854 66506 146906
rect 66558 146854 66570 146906
rect 66622 146854 97034 146906
rect 97086 146854 97098 146906
rect 97150 146854 97162 146906
rect 97214 146854 97226 146906
rect 97278 146854 97290 146906
rect 97342 146854 108836 146906
rect 1104 146832 108836 146854
rect 1104 146362 108836 146384
rect 1104 146310 4214 146362
rect 4266 146310 4278 146362
rect 4330 146310 4342 146362
rect 4394 146310 4406 146362
rect 4458 146310 4470 146362
rect 4522 146310 34934 146362
rect 34986 146310 34998 146362
rect 35050 146310 35062 146362
rect 35114 146310 35126 146362
rect 35178 146310 35190 146362
rect 35242 146310 65654 146362
rect 65706 146310 65718 146362
rect 65770 146310 65782 146362
rect 65834 146310 65846 146362
rect 65898 146310 65910 146362
rect 65962 146310 96374 146362
rect 96426 146310 96438 146362
rect 96490 146310 96502 146362
rect 96554 146310 96566 146362
rect 96618 146310 96630 146362
rect 96682 146310 108836 146362
rect 1104 146288 108836 146310
rect 1104 145818 108836 145840
rect 1104 145766 4874 145818
rect 4926 145766 4938 145818
rect 4990 145766 5002 145818
rect 5054 145766 5066 145818
rect 5118 145766 5130 145818
rect 5182 145766 35594 145818
rect 35646 145766 35658 145818
rect 35710 145766 35722 145818
rect 35774 145766 35786 145818
rect 35838 145766 35850 145818
rect 35902 145766 66314 145818
rect 66366 145766 66378 145818
rect 66430 145766 66442 145818
rect 66494 145766 66506 145818
rect 66558 145766 66570 145818
rect 66622 145766 97034 145818
rect 97086 145766 97098 145818
rect 97150 145766 97162 145818
rect 97214 145766 97226 145818
rect 97278 145766 97290 145818
rect 97342 145766 108836 145818
rect 1104 145744 108836 145766
rect 1104 145274 108836 145296
rect 1104 145222 4214 145274
rect 4266 145222 4278 145274
rect 4330 145222 4342 145274
rect 4394 145222 4406 145274
rect 4458 145222 4470 145274
rect 4522 145222 34934 145274
rect 34986 145222 34998 145274
rect 35050 145222 35062 145274
rect 35114 145222 35126 145274
rect 35178 145222 35190 145274
rect 35242 145222 65654 145274
rect 65706 145222 65718 145274
rect 65770 145222 65782 145274
rect 65834 145222 65846 145274
rect 65898 145222 65910 145274
rect 65962 145222 96374 145274
rect 96426 145222 96438 145274
rect 96490 145222 96502 145274
rect 96554 145222 96566 145274
rect 96618 145222 96630 145274
rect 96682 145222 108836 145274
rect 1104 145200 108836 145222
rect 1104 144730 108836 144752
rect 1104 144678 4874 144730
rect 4926 144678 4938 144730
rect 4990 144678 5002 144730
rect 5054 144678 5066 144730
rect 5118 144678 5130 144730
rect 5182 144678 35594 144730
rect 35646 144678 35658 144730
rect 35710 144678 35722 144730
rect 35774 144678 35786 144730
rect 35838 144678 35850 144730
rect 35902 144678 66314 144730
rect 66366 144678 66378 144730
rect 66430 144678 66442 144730
rect 66494 144678 66506 144730
rect 66558 144678 66570 144730
rect 66622 144678 97034 144730
rect 97086 144678 97098 144730
rect 97150 144678 97162 144730
rect 97214 144678 97226 144730
rect 97278 144678 97290 144730
rect 97342 144678 108836 144730
rect 1104 144656 108836 144678
rect 1104 144186 108836 144208
rect 1104 144134 4214 144186
rect 4266 144134 4278 144186
rect 4330 144134 4342 144186
rect 4394 144134 4406 144186
rect 4458 144134 4470 144186
rect 4522 144134 34934 144186
rect 34986 144134 34998 144186
rect 35050 144134 35062 144186
rect 35114 144134 35126 144186
rect 35178 144134 35190 144186
rect 35242 144134 65654 144186
rect 65706 144134 65718 144186
rect 65770 144134 65782 144186
rect 65834 144134 65846 144186
rect 65898 144134 65910 144186
rect 65962 144134 96374 144186
rect 96426 144134 96438 144186
rect 96490 144134 96502 144186
rect 96554 144134 96566 144186
rect 96618 144134 96630 144186
rect 96682 144134 108836 144186
rect 1104 144112 108836 144134
rect 1104 143642 108836 143664
rect 1104 143590 4874 143642
rect 4926 143590 4938 143642
rect 4990 143590 5002 143642
rect 5054 143590 5066 143642
rect 5118 143590 5130 143642
rect 5182 143590 35594 143642
rect 35646 143590 35658 143642
rect 35710 143590 35722 143642
rect 35774 143590 35786 143642
rect 35838 143590 35850 143642
rect 35902 143590 66314 143642
rect 66366 143590 66378 143642
rect 66430 143590 66442 143642
rect 66494 143590 66506 143642
rect 66558 143590 66570 143642
rect 66622 143590 97034 143642
rect 97086 143590 97098 143642
rect 97150 143590 97162 143642
rect 97214 143590 97226 143642
rect 97278 143590 97290 143642
rect 97342 143590 108836 143642
rect 1104 143568 108836 143590
rect 1104 143098 108836 143120
rect 1104 143046 4214 143098
rect 4266 143046 4278 143098
rect 4330 143046 4342 143098
rect 4394 143046 4406 143098
rect 4458 143046 4470 143098
rect 4522 143046 34934 143098
rect 34986 143046 34998 143098
rect 35050 143046 35062 143098
rect 35114 143046 35126 143098
rect 35178 143046 35190 143098
rect 35242 143046 65654 143098
rect 65706 143046 65718 143098
rect 65770 143046 65782 143098
rect 65834 143046 65846 143098
rect 65898 143046 65910 143098
rect 65962 143046 96374 143098
rect 96426 143046 96438 143098
rect 96490 143046 96502 143098
rect 96554 143046 96566 143098
rect 96618 143046 96630 143098
rect 96682 143046 108836 143098
rect 1104 143024 108836 143046
rect 1104 142554 108836 142576
rect 1104 142502 4874 142554
rect 4926 142502 4938 142554
rect 4990 142502 5002 142554
rect 5054 142502 5066 142554
rect 5118 142502 5130 142554
rect 5182 142502 35594 142554
rect 35646 142502 35658 142554
rect 35710 142502 35722 142554
rect 35774 142502 35786 142554
rect 35838 142502 35850 142554
rect 35902 142502 66314 142554
rect 66366 142502 66378 142554
rect 66430 142502 66442 142554
rect 66494 142502 66506 142554
rect 66558 142502 66570 142554
rect 66622 142502 97034 142554
rect 97086 142502 97098 142554
rect 97150 142502 97162 142554
rect 97214 142502 97226 142554
rect 97278 142502 97290 142554
rect 97342 142502 108836 142554
rect 1104 142480 108836 142502
rect 1104 142010 108836 142032
rect 1104 141958 4214 142010
rect 4266 141958 4278 142010
rect 4330 141958 4342 142010
rect 4394 141958 4406 142010
rect 4458 141958 4470 142010
rect 4522 141958 34934 142010
rect 34986 141958 34998 142010
rect 35050 141958 35062 142010
rect 35114 141958 35126 142010
rect 35178 141958 35190 142010
rect 35242 141958 65654 142010
rect 65706 141958 65718 142010
rect 65770 141958 65782 142010
rect 65834 141958 65846 142010
rect 65898 141958 65910 142010
rect 65962 141958 96374 142010
rect 96426 141958 96438 142010
rect 96490 141958 96502 142010
rect 96554 141958 96566 142010
rect 96618 141958 96630 142010
rect 96682 141958 108836 142010
rect 1104 141936 108836 141958
rect 1104 141466 108836 141488
rect 1104 141414 4874 141466
rect 4926 141414 4938 141466
rect 4990 141414 5002 141466
rect 5054 141414 5066 141466
rect 5118 141414 5130 141466
rect 5182 141414 35594 141466
rect 35646 141414 35658 141466
rect 35710 141414 35722 141466
rect 35774 141414 35786 141466
rect 35838 141414 35850 141466
rect 35902 141414 66314 141466
rect 66366 141414 66378 141466
rect 66430 141414 66442 141466
rect 66494 141414 66506 141466
rect 66558 141414 66570 141466
rect 66622 141414 97034 141466
rect 97086 141414 97098 141466
rect 97150 141414 97162 141466
rect 97214 141414 97226 141466
rect 97278 141414 97290 141466
rect 97342 141414 108836 141466
rect 1104 141392 108836 141414
rect 1104 140922 108836 140944
rect 1104 140870 4214 140922
rect 4266 140870 4278 140922
rect 4330 140870 4342 140922
rect 4394 140870 4406 140922
rect 4458 140870 4470 140922
rect 4522 140870 34934 140922
rect 34986 140870 34998 140922
rect 35050 140870 35062 140922
rect 35114 140870 35126 140922
rect 35178 140870 35190 140922
rect 35242 140870 65654 140922
rect 65706 140870 65718 140922
rect 65770 140870 65782 140922
rect 65834 140870 65846 140922
rect 65898 140870 65910 140922
rect 65962 140870 96374 140922
rect 96426 140870 96438 140922
rect 96490 140870 96502 140922
rect 96554 140870 96566 140922
rect 96618 140870 96630 140922
rect 96682 140870 108836 140922
rect 1104 140848 108836 140870
rect 1104 140378 108836 140400
rect 1104 140326 4874 140378
rect 4926 140326 4938 140378
rect 4990 140326 5002 140378
rect 5054 140326 5066 140378
rect 5118 140326 5130 140378
rect 5182 140326 35594 140378
rect 35646 140326 35658 140378
rect 35710 140326 35722 140378
rect 35774 140326 35786 140378
rect 35838 140326 35850 140378
rect 35902 140326 66314 140378
rect 66366 140326 66378 140378
rect 66430 140326 66442 140378
rect 66494 140326 66506 140378
rect 66558 140326 66570 140378
rect 66622 140326 97034 140378
rect 97086 140326 97098 140378
rect 97150 140326 97162 140378
rect 97214 140326 97226 140378
rect 97278 140326 97290 140378
rect 97342 140326 108836 140378
rect 1104 140304 108836 140326
rect 1104 139834 108836 139856
rect 1104 139782 4214 139834
rect 4266 139782 4278 139834
rect 4330 139782 4342 139834
rect 4394 139782 4406 139834
rect 4458 139782 4470 139834
rect 4522 139782 34934 139834
rect 34986 139782 34998 139834
rect 35050 139782 35062 139834
rect 35114 139782 35126 139834
rect 35178 139782 35190 139834
rect 35242 139782 65654 139834
rect 65706 139782 65718 139834
rect 65770 139782 65782 139834
rect 65834 139782 65846 139834
rect 65898 139782 65910 139834
rect 65962 139782 96374 139834
rect 96426 139782 96438 139834
rect 96490 139782 96502 139834
rect 96554 139782 96566 139834
rect 96618 139782 96630 139834
rect 96682 139782 108836 139834
rect 1104 139760 108836 139782
rect 1104 139290 108836 139312
rect 1104 139238 4874 139290
rect 4926 139238 4938 139290
rect 4990 139238 5002 139290
rect 5054 139238 5066 139290
rect 5118 139238 5130 139290
rect 5182 139238 35594 139290
rect 35646 139238 35658 139290
rect 35710 139238 35722 139290
rect 35774 139238 35786 139290
rect 35838 139238 35850 139290
rect 35902 139238 66314 139290
rect 66366 139238 66378 139290
rect 66430 139238 66442 139290
rect 66494 139238 66506 139290
rect 66558 139238 66570 139290
rect 66622 139238 97034 139290
rect 97086 139238 97098 139290
rect 97150 139238 97162 139290
rect 97214 139238 97226 139290
rect 97278 139238 97290 139290
rect 97342 139238 108836 139290
rect 1104 139216 108836 139238
rect 1104 138746 108836 138768
rect 1104 138694 4214 138746
rect 4266 138694 4278 138746
rect 4330 138694 4342 138746
rect 4394 138694 4406 138746
rect 4458 138694 4470 138746
rect 4522 138694 34934 138746
rect 34986 138694 34998 138746
rect 35050 138694 35062 138746
rect 35114 138694 35126 138746
rect 35178 138694 35190 138746
rect 35242 138694 65654 138746
rect 65706 138694 65718 138746
rect 65770 138694 65782 138746
rect 65834 138694 65846 138746
rect 65898 138694 65910 138746
rect 65962 138694 96374 138746
rect 96426 138694 96438 138746
rect 96490 138694 96502 138746
rect 96554 138694 96566 138746
rect 96618 138694 96630 138746
rect 96682 138694 108836 138746
rect 1104 138672 108836 138694
rect 1104 138202 108836 138224
rect 1104 138150 4874 138202
rect 4926 138150 4938 138202
rect 4990 138150 5002 138202
rect 5054 138150 5066 138202
rect 5118 138150 5130 138202
rect 5182 138150 35594 138202
rect 35646 138150 35658 138202
rect 35710 138150 35722 138202
rect 35774 138150 35786 138202
rect 35838 138150 35850 138202
rect 35902 138150 66314 138202
rect 66366 138150 66378 138202
rect 66430 138150 66442 138202
rect 66494 138150 66506 138202
rect 66558 138150 66570 138202
rect 66622 138150 97034 138202
rect 97086 138150 97098 138202
rect 97150 138150 97162 138202
rect 97214 138150 97226 138202
rect 97278 138150 97290 138202
rect 97342 138150 108836 138202
rect 1104 138128 108836 138150
rect 1104 137658 108836 137680
rect 1104 137606 4214 137658
rect 4266 137606 4278 137658
rect 4330 137606 4342 137658
rect 4394 137606 4406 137658
rect 4458 137606 4470 137658
rect 4522 137606 34934 137658
rect 34986 137606 34998 137658
rect 35050 137606 35062 137658
rect 35114 137606 35126 137658
rect 35178 137606 35190 137658
rect 35242 137606 65654 137658
rect 65706 137606 65718 137658
rect 65770 137606 65782 137658
rect 65834 137606 65846 137658
rect 65898 137606 65910 137658
rect 65962 137606 96374 137658
rect 96426 137606 96438 137658
rect 96490 137606 96502 137658
rect 96554 137606 96566 137658
rect 96618 137606 96630 137658
rect 96682 137606 108836 137658
rect 1104 137584 108836 137606
rect 1104 137114 108836 137136
rect 1104 137062 4874 137114
rect 4926 137062 4938 137114
rect 4990 137062 5002 137114
rect 5054 137062 5066 137114
rect 5118 137062 5130 137114
rect 5182 137062 35594 137114
rect 35646 137062 35658 137114
rect 35710 137062 35722 137114
rect 35774 137062 35786 137114
rect 35838 137062 35850 137114
rect 35902 137062 66314 137114
rect 66366 137062 66378 137114
rect 66430 137062 66442 137114
rect 66494 137062 66506 137114
rect 66558 137062 66570 137114
rect 66622 137062 97034 137114
rect 97086 137062 97098 137114
rect 97150 137062 97162 137114
rect 97214 137062 97226 137114
rect 97278 137062 97290 137114
rect 97342 137062 108836 137114
rect 1104 137040 108836 137062
rect 1104 136570 108836 136592
rect 1104 136518 4214 136570
rect 4266 136518 4278 136570
rect 4330 136518 4342 136570
rect 4394 136518 4406 136570
rect 4458 136518 4470 136570
rect 4522 136518 34934 136570
rect 34986 136518 34998 136570
rect 35050 136518 35062 136570
rect 35114 136518 35126 136570
rect 35178 136518 35190 136570
rect 35242 136518 65654 136570
rect 65706 136518 65718 136570
rect 65770 136518 65782 136570
rect 65834 136518 65846 136570
rect 65898 136518 65910 136570
rect 65962 136518 96374 136570
rect 96426 136518 96438 136570
rect 96490 136518 96502 136570
rect 96554 136518 96566 136570
rect 96618 136518 96630 136570
rect 96682 136518 105922 136570
rect 105974 136518 105986 136570
rect 106038 136518 106050 136570
rect 106102 136518 106114 136570
rect 106166 136518 106178 136570
rect 106230 136518 108836 136570
rect 1104 136496 108836 136518
rect 47581 136255 47639 136261
rect 47581 136252 47593 136255
rect 26206 136224 47593 136252
rect 9490 136076 9496 136128
rect 9548 136116 9554 136128
rect 26206 136116 26234 136224
rect 47581 136221 47593 136224
rect 47627 136252 47639 136255
rect 47949 136255 48007 136261
rect 47949 136252 47961 136255
rect 47627 136224 47961 136252
rect 47627 136221 47639 136224
rect 47581 136215 47639 136221
rect 47949 136221 47961 136224
rect 47995 136221 48007 136255
rect 47949 136215 48007 136221
rect 53745 136255 53803 136261
rect 53745 136221 53757 136255
rect 53791 136252 53803 136255
rect 53929 136255 53987 136261
rect 53929 136252 53941 136255
rect 53791 136224 53941 136252
rect 53791 136221 53803 136224
rect 53745 136215 53803 136221
rect 53929 136221 53941 136224
rect 53975 136252 53987 136255
rect 101950 136252 101956 136264
rect 53975 136224 101956 136252
rect 53975 136221 53987 136224
rect 53929 136215 53987 136221
rect 101950 136212 101956 136224
rect 102008 136212 102014 136264
rect 38194 136144 38200 136196
rect 38252 136144 38258 136196
rect 40678 136144 40684 136196
rect 40736 136144 40742 136196
rect 42978 136144 42984 136196
rect 43036 136144 43042 136196
rect 45281 136187 45339 136193
rect 45281 136153 45293 136187
rect 45327 136184 45339 136187
rect 46014 136184 46020 136196
rect 45327 136156 46020 136184
rect 45327 136153 45339 136156
rect 45281 136147 45339 136153
rect 46014 136144 46020 136156
rect 46072 136144 46078 136196
rect 47765 136187 47823 136193
rect 47765 136153 47777 136187
rect 47811 136184 47823 136187
rect 48498 136184 48504 136196
rect 47811 136156 48504 136184
rect 47811 136153 47823 136156
rect 47765 136147 47823 136153
rect 48498 136144 48504 136156
rect 48556 136144 48562 136196
rect 52362 136144 52368 136196
rect 52420 136184 52426 136196
rect 53561 136187 53619 136193
rect 53561 136184 53573 136187
rect 52420 136156 53573 136184
rect 52420 136144 52426 136156
rect 53561 136153 53573 136156
rect 53607 136153 53619 136187
rect 53561 136147 53619 136153
rect 55766 136144 55772 136196
rect 55824 136144 55830 136196
rect 58158 136144 58164 136196
rect 58216 136144 58222 136196
rect 60642 136144 60648 136196
rect 60700 136144 60706 136196
rect 63126 136144 63132 136196
rect 63184 136144 63190 136196
rect 64414 136144 64420 136196
rect 64472 136184 64478 136196
rect 64969 136187 65027 136193
rect 64969 136184 64981 136187
rect 64472 136156 64981 136184
rect 64472 136144 64478 136156
rect 64969 136153 64981 136156
rect 65015 136153 65027 136187
rect 64969 136147 65027 136153
rect 67542 136144 67548 136196
rect 67600 136144 67606 136196
rect 69750 136144 69756 136196
rect 69808 136144 69814 136196
rect 72142 136144 72148 136196
rect 72200 136144 72206 136196
rect 74166 136144 74172 136196
rect 74224 136144 74230 136196
rect 9548 136088 26234 136116
rect 9548 136076 9554 136088
rect 36078 136076 36084 136128
rect 36136 136076 36142 136128
rect 38102 136076 38108 136128
rect 38160 136116 38166 136128
rect 38381 136119 38439 136125
rect 38381 136116 38393 136119
rect 38160 136088 38393 136116
rect 38160 136076 38166 136088
rect 38381 136085 38393 136088
rect 38427 136085 38439 136119
rect 38381 136079 38439 136085
rect 40586 136076 40592 136128
rect 40644 136116 40650 136128
rect 40865 136119 40923 136125
rect 40865 136116 40877 136119
rect 40644 136088 40877 136116
rect 40644 136076 40650 136088
rect 40865 136085 40877 136088
rect 40911 136085 40923 136119
rect 40865 136079 40923 136085
rect 42886 136076 42892 136128
rect 42944 136116 42950 136128
rect 43165 136119 43223 136125
rect 43165 136116 43177 136119
rect 42944 136088 43177 136116
rect 42944 136076 42950 136088
rect 43165 136085 43177 136088
rect 43211 136085 43223 136119
rect 43165 136079 43223 136085
rect 45186 136076 45192 136128
rect 45244 136116 45250 136128
rect 45465 136119 45523 136125
rect 45465 136116 45477 136119
rect 45244 136088 45477 136116
rect 45244 136076 45250 136088
rect 45465 136085 45477 136088
rect 45511 136085 45523 136119
rect 45465 136079 45523 136085
rect 55861 136119 55919 136125
rect 55861 136085 55873 136119
rect 55907 136116 55919 136119
rect 56134 136116 56140 136128
rect 55907 136088 56140 136116
rect 55907 136085 55919 136088
rect 55861 136079 55919 136085
rect 56134 136076 56140 136088
rect 56192 136076 56198 136128
rect 58253 136119 58311 136125
rect 58253 136085 58265 136119
rect 58299 136116 58311 136119
rect 58526 136116 58532 136128
rect 58299 136088 58532 136116
rect 58299 136085 58311 136088
rect 58253 136079 58311 136085
rect 58526 136076 58532 136088
rect 58584 136076 58590 136128
rect 60737 136119 60795 136125
rect 60737 136085 60749 136119
rect 60783 136116 60795 136119
rect 61010 136116 61016 136128
rect 60783 136088 61016 136116
rect 60783 136085 60795 136088
rect 60737 136079 60795 136085
rect 61010 136076 61016 136088
rect 61068 136076 61074 136128
rect 63221 136119 63279 136125
rect 63221 136085 63233 136119
rect 63267 136116 63279 136119
rect 63494 136116 63500 136128
rect 63267 136088 63500 136116
rect 63267 136085 63279 136088
rect 63221 136079 63279 136085
rect 63494 136076 63500 136088
rect 63552 136076 63558 136128
rect 65061 136119 65119 136125
rect 65061 136085 65073 136119
rect 65107 136116 65119 136119
rect 65334 136116 65340 136128
rect 65107 136088 65340 136116
rect 65107 136085 65119 136088
rect 65061 136079 65119 136085
rect 65334 136076 65340 136088
rect 65392 136076 65398 136128
rect 67637 136119 67695 136125
rect 67637 136085 67649 136119
rect 67683 136116 67695 136119
rect 67910 136116 67916 136128
rect 67683 136088 67916 136116
rect 67683 136085 67695 136088
rect 67637 136079 67695 136085
rect 67910 136076 67916 136088
rect 67968 136076 67974 136128
rect 69845 136119 69903 136125
rect 69845 136085 69857 136119
rect 69891 136116 69903 136119
rect 70118 136116 70124 136128
rect 69891 136088 70124 136116
rect 69891 136085 69903 136088
rect 69845 136079 69903 136085
rect 70118 136076 70124 136088
rect 70176 136076 70182 136128
rect 72237 136119 72295 136125
rect 72237 136085 72249 136119
rect 72283 136116 72295 136119
rect 72510 136116 72516 136128
rect 72283 136088 72516 136116
rect 72283 136085 72295 136088
rect 72237 136079 72295 136085
rect 72510 136076 72516 136088
rect 72568 136076 72574 136128
rect 74261 136119 74319 136125
rect 74261 136085 74273 136119
rect 74307 136116 74319 136119
rect 74537 136119 74595 136125
rect 74537 136116 74549 136119
rect 74307 136088 74549 136116
rect 74307 136085 74319 136088
rect 74261 136079 74319 136085
rect 74537 136085 74549 136088
rect 74583 136116 74595 136119
rect 77754 136116 77760 136128
rect 74583 136088 77760 136116
rect 74583 136085 74595 136088
rect 74537 136079 74595 136085
rect 77754 136076 77760 136088
rect 77812 136076 77818 136128
rect 86126 136076 86132 136128
rect 86184 136116 86190 136128
rect 86221 136119 86279 136125
rect 86221 136116 86233 136119
rect 86184 136088 86233 136116
rect 86184 136076 86190 136088
rect 86221 136085 86233 136088
rect 86267 136085 86279 136119
rect 86221 136079 86279 136085
rect 87322 136076 87328 136128
rect 87380 136076 87386 136128
rect 95970 136076 95976 136128
rect 96028 136076 96034 136128
rect 1104 136026 108836 136048
rect 1104 135974 4874 136026
rect 4926 135974 4938 136026
rect 4990 135974 5002 136026
rect 5054 135974 5066 136026
rect 5118 135974 5130 136026
rect 5182 135974 35594 136026
rect 35646 135974 35658 136026
rect 35710 135974 35722 136026
rect 35774 135974 35786 136026
rect 35838 135974 35850 136026
rect 35902 135974 66314 136026
rect 66366 135974 66378 136026
rect 66430 135974 66442 136026
rect 66494 135974 66506 136026
rect 66558 135974 66570 136026
rect 66622 135974 97034 136026
rect 97086 135974 97098 136026
rect 97150 135974 97162 136026
rect 97214 135974 97226 136026
rect 97278 135974 97290 136026
rect 97342 135974 106658 136026
rect 106710 135974 106722 136026
rect 106774 135974 106786 136026
rect 106838 135974 106850 136026
rect 106902 135974 106914 136026
rect 106966 135974 108836 136026
rect 1104 135952 108836 135974
rect 8110 135872 8116 135924
rect 8168 135912 8174 135924
rect 45186 135912 45192 135924
rect 8168 135884 45192 135912
rect 8168 135872 8174 135884
rect 45186 135872 45192 135884
rect 45244 135872 45250 135924
rect 56134 135872 56140 135924
rect 56192 135912 56198 135924
rect 102134 135912 102140 135924
rect 56192 135884 102140 135912
rect 56192 135872 56198 135884
rect 102134 135872 102140 135884
rect 102192 135872 102198 135924
rect 8202 135804 8208 135856
rect 8260 135844 8266 135856
rect 42886 135844 42892 135856
rect 8260 135816 42892 135844
rect 8260 135804 8266 135816
rect 42886 135804 42892 135816
rect 42944 135804 42950 135856
rect 58526 135804 58532 135856
rect 58584 135844 58590 135856
rect 103974 135844 103980 135856
rect 58584 135816 103980 135844
rect 58584 135804 58590 135816
rect 103974 135804 103980 135816
rect 104032 135804 104038 135856
rect 9582 135736 9588 135788
rect 9640 135776 9646 135788
rect 40586 135776 40592 135788
rect 9640 135748 40592 135776
rect 9640 135736 9646 135748
rect 40586 135736 40592 135748
rect 40644 135736 40650 135788
rect 61010 135736 61016 135788
rect 61068 135776 61074 135788
rect 102318 135776 102324 135788
rect 61068 135748 102324 135776
rect 61068 135736 61074 135748
rect 102318 135736 102324 135748
rect 102376 135736 102382 135788
rect 8018 135668 8024 135720
rect 8076 135708 8082 135720
rect 38102 135708 38108 135720
rect 8076 135680 38108 135708
rect 8076 135668 8082 135680
rect 38102 135668 38108 135680
rect 38160 135668 38166 135720
rect 63494 135668 63500 135720
rect 63552 135708 63558 135720
rect 102410 135708 102416 135720
rect 63552 135680 102416 135708
rect 63552 135668 63558 135680
rect 102410 135668 102416 135680
rect 102468 135668 102474 135720
rect 65334 135600 65340 135652
rect 65392 135640 65398 135652
rect 103606 135640 103612 135652
rect 65392 135612 103612 135640
rect 65392 135600 65398 135612
rect 103606 135600 103612 135612
rect 103664 135600 103670 135652
rect 67910 135532 67916 135584
rect 67968 135572 67974 135584
rect 103698 135572 103704 135584
rect 67968 135544 103704 135572
rect 67968 135532 67974 135544
rect 103698 135532 103704 135544
rect 103756 135532 103762 135584
rect 1104 135482 7912 135504
rect 1104 135430 4214 135482
rect 4266 135430 4278 135482
rect 4330 135430 4342 135482
rect 4394 135430 4406 135482
rect 4458 135430 4470 135482
rect 4522 135430 7912 135482
rect 70118 135464 70124 135516
rect 70176 135504 70182 135516
rect 102502 135504 102508 135516
rect 70176 135476 102508 135504
rect 70176 135464 70182 135476
rect 102502 135464 102508 135476
rect 102560 135464 102566 135516
rect 104052 135482 108836 135504
rect 1104 135408 7912 135430
rect 72510 135396 72516 135448
rect 72568 135436 72574 135448
rect 103882 135436 103888 135448
rect 72568 135408 103888 135436
rect 72568 135396 72574 135408
rect 103882 135396 103888 135408
rect 103940 135396 103946 135448
rect 104052 135430 105922 135482
rect 105974 135430 105986 135482
rect 106038 135430 106050 135482
rect 106102 135430 106114 135482
rect 106166 135430 106178 135482
rect 106230 135430 108836 135482
rect 104052 135408 108836 135430
rect 77754 135328 77760 135380
rect 77812 135368 77818 135380
rect 103790 135368 103796 135380
rect 77812 135340 103796 135368
rect 77812 135328 77818 135340
rect 103790 135328 103796 135340
rect 103848 135328 103854 135380
rect 1104 134938 7912 134960
rect 1104 134886 4874 134938
rect 4926 134886 4938 134938
rect 4990 134886 5002 134938
rect 5054 134886 5066 134938
rect 5118 134886 5130 134938
rect 5182 134886 7912 134938
rect 1104 134864 7912 134886
rect 104052 134938 108836 134960
rect 104052 134886 106658 134938
rect 106710 134886 106722 134938
rect 106774 134886 106786 134938
rect 106838 134886 106850 134938
rect 106902 134886 106914 134938
rect 106966 134886 108836 134938
rect 104052 134864 108836 134886
rect 95970 134512 95976 134564
rect 96028 134552 96034 134564
rect 103514 134552 103520 134564
rect 96028 134524 103520 134552
rect 96028 134512 96034 134524
rect 103514 134512 103520 134524
rect 103572 134512 103578 134564
rect 1104 134394 7912 134416
rect 1104 134342 4214 134394
rect 4266 134342 4278 134394
rect 4330 134342 4342 134394
rect 4394 134342 4406 134394
rect 4458 134342 4470 134394
rect 4522 134342 7912 134394
rect 1104 134320 7912 134342
rect 104052 134394 108836 134416
rect 104052 134342 105922 134394
rect 105974 134342 105986 134394
rect 106038 134342 106050 134394
rect 106102 134342 106114 134394
rect 106166 134342 106178 134394
rect 106230 134342 108836 134394
rect 104052 134320 108836 134342
rect 87322 133968 87328 134020
rect 87380 134008 87386 134020
rect 102226 134008 102232 134020
rect 87380 133980 102232 134008
rect 87380 133968 87386 133980
rect 102226 133968 102232 133980
rect 102284 133968 102290 134020
rect 7926 133900 7932 133952
rect 7984 133940 7990 133952
rect 36078 133940 36084 133952
rect 7984 133912 36084 133940
rect 7984 133900 7990 133912
rect 36078 133900 36084 133912
rect 36136 133900 36142 133952
rect 86126 133900 86132 133952
rect 86184 133940 86190 133952
rect 102594 133940 102600 133952
rect 86184 133912 102600 133940
rect 86184 133900 86190 133912
rect 102594 133900 102600 133912
rect 102652 133900 102658 133952
rect 1104 133850 7912 133872
rect 1104 133798 4874 133850
rect 4926 133798 4938 133850
rect 4990 133798 5002 133850
rect 5054 133798 5066 133850
rect 5118 133798 5130 133850
rect 5182 133798 7912 133850
rect 1104 133776 7912 133798
rect 104052 133850 108836 133872
rect 104052 133798 106658 133850
rect 106710 133798 106722 133850
rect 106774 133798 106786 133850
rect 106838 133798 106850 133850
rect 106902 133798 106914 133850
rect 106966 133798 108836 133850
rect 104052 133776 108836 133798
rect 1104 133306 7912 133328
rect 1104 133254 4214 133306
rect 4266 133254 4278 133306
rect 4330 133254 4342 133306
rect 4394 133254 4406 133306
rect 4458 133254 4470 133306
rect 4522 133254 7912 133306
rect 1104 133232 7912 133254
rect 104052 133306 108836 133328
rect 104052 133254 105922 133306
rect 105974 133254 105986 133306
rect 106038 133254 106050 133306
rect 106102 133254 106114 133306
rect 106166 133254 106178 133306
rect 106230 133254 108836 133306
rect 104052 133232 108836 133254
rect 1104 132762 7912 132784
rect 1104 132710 4874 132762
rect 4926 132710 4938 132762
rect 4990 132710 5002 132762
rect 5054 132710 5066 132762
rect 5118 132710 5130 132762
rect 5182 132710 7912 132762
rect 1104 132688 7912 132710
rect 104052 132762 108836 132784
rect 104052 132710 106658 132762
rect 106710 132710 106722 132762
rect 106774 132710 106786 132762
rect 106838 132710 106850 132762
rect 106902 132710 106914 132762
rect 106966 132710 108836 132762
rect 104052 132688 108836 132710
rect 1104 132218 7912 132240
rect 1104 132166 4214 132218
rect 4266 132166 4278 132218
rect 4330 132166 4342 132218
rect 4394 132166 4406 132218
rect 4458 132166 4470 132218
rect 4522 132166 7912 132218
rect 1104 132144 7912 132166
rect 104052 132218 108836 132240
rect 104052 132166 105922 132218
rect 105974 132166 105986 132218
rect 106038 132166 106050 132218
rect 106102 132166 106114 132218
rect 106166 132166 106178 132218
rect 106230 132166 108836 132218
rect 104052 132144 108836 132166
rect 1104 131674 7912 131696
rect 1104 131622 4874 131674
rect 4926 131622 4938 131674
rect 4990 131622 5002 131674
rect 5054 131622 5066 131674
rect 5118 131622 5130 131674
rect 5182 131622 7912 131674
rect 1104 131600 7912 131622
rect 104052 131674 108836 131696
rect 104052 131622 106658 131674
rect 106710 131622 106722 131674
rect 106774 131622 106786 131674
rect 106838 131622 106850 131674
rect 106902 131622 106914 131674
rect 106966 131622 108836 131674
rect 104052 131600 108836 131622
rect 1104 131130 7912 131152
rect 1104 131078 4214 131130
rect 4266 131078 4278 131130
rect 4330 131078 4342 131130
rect 4394 131078 4406 131130
rect 4458 131078 4470 131130
rect 4522 131078 7912 131130
rect 1104 131056 7912 131078
rect 104052 131130 108836 131152
rect 104052 131078 105922 131130
rect 105974 131078 105986 131130
rect 106038 131078 106050 131130
rect 106102 131078 106114 131130
rect 106166 131078 106178 131130
rect 106230 131078 108836 131130
rect 104052 131056 108836 131078
rect 1104 130586 7912 130608
rect 1104 130534 4874 130586
rect 4926 130534 4938 130586
rect 4990 130534 5002 130586
rect 5054 130534 5066 130586
rect 5118 130534 5130 130586
rect 5182 130534 7912 130586
rect 1104 130512 7912 130534
rect 104052 130586 108836 130608
rect 104052 130534 106658 130586
rect 106710 130534 106722 130586
rect 106774 130534 106786 130586
rect 106838 130534 106850 130586
rect 106902 130534 106914 130586
rect 106966 130534 108836 130586
rect 104052 130512 108836 130534
rect 1104 130042 7912 130064
rect 1104 129990 4214 130042
rect 4266 129990 4278 130042
rect 4330 129990 4342 130042
rect 4394 129990 4406 130042
rect 4458 129990 4470 130042
rect 4522 129990 7912 130042
rect 1104 129968 7912 129990
rect 104052 130042 108836 130064
rect 104052 129990 105922 130042
rect 105974 129990 105986 130042
rect 106038 129990 106050 130042
rect 106102 129990 106114 130042
rect 106166 129990 106178 130042
rect 106230 129990 108836 130042
rect 104052 129968 108836 129990
rect 104342 129820 104348 129872
rect 104400 129820 104406 129872
rect 1104 129498 7912 129520
rect 1104 129446 4874 129498
rect 4926 129446 4938 129498
rect 4990 129446 5002 129498
rect 5054 129446 5066 129498
rect 5118 129446 5130 129498
rect 5182 129446 7912 129498
rect 1104 129424 7912 129446
rect 104052 129498 108836 129520
rect 104052 129446 106658 129498
rect 106710 129446 106722 129498
rect 106774 129446 106786 129498
rect 106838 129446 106850 129498
rect 106902 129446 106914 129498
rect 106966 129446 108836 129498
rect 104052 129424 108836 129446
rect 1104 128954 7912 128976
rect 1104 128902 4214 128954
rect 4266 128902 4278 128954
rect 4330 128902 4342 128954
rect 4394 128902 4406 128954
rect 4458 128902 4470 128954
rect 4522 128902 7912 128954
rect 1104 128880 7912 128902
rect 104052 128954 108836 128976
rect 104052 128902 105922 128954
rect 105974 128902 105986 128954
rect 106038 128902 106050 128954
rect 106102 128902 106114 128954
rect 106166 128902 106178 128954
rect 106230 128902 108836 128954
rect 104052 128880 108836 128902
rect 1104 128410 7912 128432
rect 1104 128358 4874 128410
rect 4926 128358 4938 128410
rect 4990 128358 5002 128410
rect 5054 128358 5066 128410
rect 5118 128358 5130 128410
rect 5182 128358 7912 128410
rect 1104 128336 7912 128358
rect 104052 128410 108836 128432
rect 104052 128358 106658 128410
rect 106710 128358 106722 128410
rect 106774 128358 106786 128410
rect 106838 128358 106850 128410
rect 106902 128358 106914 128410
rect 106966 128358 108836 128410
rect 104052 128336 108836 128358
rect 1104 127866 7912 127888
rect 1104 127814 4214 127866
rect 4266 127814 4278 127866
rect 4330 127814 4342 127866
rect 4394 127814 4406 127866
rect 4458 127814 4470 127866
rect 4522 127814 7912 127866
rect 1104 127792 7912 127814
rect 104052 127866 108836 127888
rect 104052 127814 105922 127866
rect 105974 127814 105986 127866
rect 106038 127814 106050 127866
rect 106102 127814 106114 127866
rect 106166 127814 106178 127866
rect 106230 127814 108836 127866
rect 104052 127792 108836 127814
rect 1104 127322 7912 127344
rect 1104 127270 4874 127322
rect 4926 127270 4938 127322
rect 4990 127270 5002 127322
rect 5054 127270 5066 127322
rect 5118 127270 5130 127322
rect 5182 127270 7912 127322
rect 1104 127248 7912 127270
rect 104052 127322 108836 127344
rect 104052 127270 106658 127322
rect 106710 127270 106722 127322
rect 106774 127270 106786 127322
rect 106838 127270 106850 127322
rect 106902 127270 106914 127322
rect 106966 127270 108836 127322
rect 104052 127248 108836 127270
rect 1104 126778 7912 126800
rect 1104 126726 4214 126778
rect 4266 126726 4278 126778
rect 4330 126726 4342 126778
rect 4394 126726 4406 126778
rect 4458 126726 4470 126778
rect 4522 126726 7912 126778
rect 1104 126704 7912 126726
rect 104052 126778 108836 126800
rect 104052 126726 105922 126778
rect 105974 126726 105986 126778
rect 106038 126726 106050 126778
rect 106102 126726 106114 126778
rect 106166 126726 106178 126778
rect 106230 126726 108836 126778
rect 104052 126704 108836 126726
rect 1104 126234 7912 126256
rect 1104 126182 4874 126234
rect 4926 126182 4938 126234
rect 4990 126182 5002 126234
rect 5054 126182 5066 126234
rect 5118 126182 5130 126234
rect 5182 126182 7912 126234
rect 1104 126160 7912 126182
rect 104052 126234 108836 126256
rect 104052 126182 106658 126234
rect 106710 126182 106722 126234
rect 106774 126182 106786 126234
rect 106838 126182 106850 126234
rect 106902 126182 106914 126234
rect 106966 126182 108836 126234
rect 104052 126160 108836 126182
rect 1104 125690 7912 125712
rect 1104 125638 4214 125690
rect 4266 125638 4278 125690
rect 4330 125638 4342 125690
rect 4394 125638 4406 125690
rect 4458 125638 4470 125690
rect 4522 125638 7912 125690
rect 1104 125616 7912 125638
rect 104052 125690 108836 125712
rect 104052 125638 105922 125690
rect 105974 125638 105986 125690
rect 106038 125638 106050 125690
rect 106102 125638 106114 125690
rect 106166 125638 106178 125690
rect 106230 125638 108836 125690
rect 104052 125616 108836 125638
rect 1104 125146 7912 125168
rect 1104 125094 4874 125146
rect 4926 125094 4938 125146
rect 4990 125094 5002 125146
rect 5054 125094 5066 125146
rect 5118 125094 5130 125146
rect 5182 125094 7912 125146
rect 1104 125072 7912 125094
rect 104052 125146 108836 125168
rect 104052 125094 106658 125146
rect 106710 125094 106722 125146
rect 106774 125094 106786 125146
rect 106838 125094 106850 125146
rect 106902 125094 106914 125146
rect 106966 125094 108836 125146
rect 104052 125072 108836 125094
rect 1104 124602 7912 124624
rect 1104 124550 4214 124602
rect 4266 124550 4278 124602
rect 4330 124550 4342 124602
rect 4394 124550 4406 124602
rect 4458 124550 4470 124602
rect 4522 124550 7912 124602
rect 1104 124528 7912 124550
rect 104052 124602 108836 124624
rect 104052 124550 105922 124602
rect 105974 124550 105986 124602
rect 106038 124550 106050 124602
rect 106102 124550 106114 124602
rect 106166 124550 106178 124602
rect 106230 124550 108836 124602
rect 104052 124528 108836 124550
rect 1104 124058 7912 124080
rect 1104 124006 4874 124058
rect 4926 124006 4938 124058
rect 4990 124006 5002 124058
rect 5054 124006 5066 124058
rect 5118 124006 5130 124058
rect 5182 124006 7912 124058
rect 1104 123984 7912 124006
rect 104052 124058 108836 124080
rect 104052 124006 106658 124058
rect 106710 124006 106722 124058
rect 106774 124006 106786 124058
rect 106838 124006 106850 124058
rect 106902 124006 106914 124058
rect 106966 124006 108836 124058
rect 104052 123984 108836 124006
rect 1104 123514 7912 123536
rect 1104 123462 4214 123514
rect 4266 123462 4278 123514
rect 4330 123462 4342 123514
rect 4394 123462 4406 123514
rect 4458 123462 4470 123514
rect 4522 123462 7912 123514
rect 1104 123440 7912 123462
rect 104052 123514 108836 123536
rect 104052 123462 105922 123514
rect 105974 123462 105986 123514
rect 106038 123462 106050 123514
rect 106102 123462 106114 123514
rect 106166 123462 106178 123514
rect 106230 123462 108836 123514
rect 104052 123440 108836 123462
rect 1104 122970 7912 122992
rect 1104 122918 4874 122970
rect 4926 122918 4938 122970
rect 4990 122918 5002 122970
rect 5054 122918 5066 122970
rect 5118 122918 5130 122970
rect 5182 122918 7912 122970
rect 1104 122896 7912 122918
rect 104052 122970 108836 122992
rect 104052 122918 106658 122970
rect 106710 122918 106722 122970
rect 106774 122918 106786 122970
rect 106838 122918 106850 122970
rect 106902 122918 106914 122970
rect 106966 122918 108836 122970
rect 104052 122896 108836 122918
rect 1104 122426 7912 122448
rect 1104 122374 4214 122426
rect 4266 122374 4278 122426
rect 4330 122374 4342 122426
rect 4394 122374 4406 122426
rect 4458 122374 4470 122426
rect 4522 122374 7912 122426
rect 1104 122352 7912 122374
rect 104052 122426 108836 122448
rect 104052 122374 105922 122426
rect 105974 122374 105986 122426
rect 106038 122374 106050 122426
rect 106102 122374 106114 122426
rect 106166 122374 106178 122426
rect 106230 122374 108836 122426
rect 104052 122352 108836 122374
rect 1104 121882 7912 121904
rect 1104 121830 4874 121882
rect 4926 121830 4938 121882
rect 4990 121830 5002 121882
rect 5054 121830 5066 121882
rect 5118 121830 5130 121882
rect 5182 121830 7912 121882
rect 1104 121808 7912 121830
rect 104052 121882 108836 121904
rect 104052 121830 106658 121882
rect 106710 121830 106722 121882
rect 106774 121830 106786 121882
rect 106838 121830 106850 121882
rect 106902 121830 106914 121882
rect 106966 121830 108836 121882
rect 104052 121808 108836 121830
rect 1104 121338 7912 121360
rect 1104 121286 4214 121338
rect 4266 121286 4278 121338
rect 4330 121286 4342 121338
rect 4394 121286 4406 121338
rect 4458 121286 4470 121338
rect 4522 121286 7912 121338
rect 1104 121264 7912 121286
rect 104052 121338 108836 121360
rect 104052 121286 105922 121338
rect 105974 121286 105986 121338
rect 106038 121286 106050 121338
rect 106102 121286 106114 121338
rect 106166 121286 106178 121338
rect 106230 121286 108836 121338
rect 104052 121264 108836 121286
rect 1104 120794 7912 120816
rect 1104 120742 4874 120794
rect 4926 120742 4938 120794
rect 4990 120742 5002 120794
rect 5054 120742 5066 120794
rect 5118 120742 5130 120794
rect 5182 120742 7912 120794
rect 1104 120720 7912 120742
rect 104052 120794 108836 120816
rect 104052 120742 106658 120794
rect 106710 120742 106722 120794
rect 106774 120742 106786 120794
rect 106838 120742 106850 120794
rect 106902 120742 106914 120794
rect 106966 120742 108836 120794
rect 104052 120720 108836 120742
rect 1104 120250 7912 120272
rect 1104 120198 4214 120250
rect 4266 120198 4278 120250
rect 4330 120198 4342 120250
rect 4394 120198 4406 120250
rect 4458 120198 4470 120250
rect 4522 120198 7912 120250
rect 1104 120176 7912 120198
rect 104052 120250 108836 120272
rect 104052 120198 105922 120250
rect 105974 120198 105986 120250
rect 106038 120198 106050 120250
rect 106102 120198 106114 120250
rect 106166 120198 106178 120250
rect 106230 120198 108836 120250
rect 104052 120176 108836 120198
rect 1104 119706 7912 119728
rect 1104 119654 4874 119706
rect 4926 119654 4938 119706
rect 4990 119654 5002 119706
rect 5054 119654 5066 119706
rect 5118 119654 5130 119706
rect 5182 119654 7912 119706
rect 1104 119632 7912 119654
rect 104052 119706 108836 119728
rect 104052 119654 106658 119706
rect 106710 119654 106722 119706
rect 106774 119654 106786 119706
rect 106838 119654 106850 119706
rect 106902 119654 106914 119706
rect 106966 119654 108836 119706
rect 104052 119632 108836 119654
rect 1104 119162 7912 119184
rect 1104 119110 4214 119162
rect 4266 119110 4278 119162
rect 4330 119110 4342 119162
rect 4394 119110 4406 119162
rect 4458 119110 4470 119162
rect 4522 119110 7912 119162
rect 1104 119088 7912 119110
rect 104052 119162 108836 119184
rect 104052 119110 105922 119162
rect 105974 119110 105986 119162
rect 106038 119110 106050 119162
rect 106102 119110 106114 119162
rect 106166 119110 106178 119162
rect 106230 119110 108836 119162
rect 104052 119088 108836 119110
rect 1104 118618 7912 118640
rect 1104 118566 4874 118618
rect 4926 118566 4938 118618
rect 4990 118566 5002 118618
rect 5054 118566 5066 118618
rect 5118 118566 5130 118618
rect 5182 118566 7912 118618
rect 1104 118544 7912 118566
rect 104052 118618 108836 118640
rect 104052 118566 106658 118618
rect 106710 118566 106722 118618
rect 106774 118566 106786 118618
rect 106838 118566 106850 118618
rect 106902 118566 106914 118618
rect 106966 118566 108836 118618
rect 104052 118544 108836 118566
rect 1104 118074 7912 118096
rect 1104 118022 4214 118074
rect 4266 118022 4278 118074
rect 4330 118022 4342 118074
rect 4394 118022 4406 118074
rect 4458 118022 4470 118074
rect 4522 118022 7912 118074
rect 1104 118000 7912 118022
rect 104052 118074 108836 118096
rect 104052 118022 105922 118074
rect 105974 118022 105986 118074
rect 106038 118022 106050 118074
rect 106102 118022 106114 118074
rect 106166 118022 106178 118074
rect 106230 118022 108836 118074
rect 104052 118000 108836 118022
rect 1104 117530 7912 117552
rect 1104 117478 4874 117530
rect 4926 117478 4938 117530
rect 4990 117478 5002 117530
rect 5054 117478 5066 117530
rect 5118 117478 5130 117530
rect 5182 117478 7912 117530
rect 1104 117456 7912 117478
rect 104052 117530 108836 117552
rect 104052 117478 106658 117530
rect 106710 117478 106722 117530
rect 106774 117478 106786 117530
rect 106838 117478 106850 117530
rect 106902 117478 106914 117530
rect 106966 117478 108836 117530
rect 104052 117456 108836 117478
rect 1104 116986 7912 117008
rect 1104 116934 4214 116986
rect 4266 116934 4278 116986
rect 4330 116934 4342 116986
rect 4394 116934 4406 116986
rect 4458 116934 4470 116986
rect 4522 116934 7912 116986
rect 1104 116912 7912 116934
rect 104052 116986 108836 117008
rect 104052 116934 105922 116986
rect 105974 116934 105986 116986
rect 106038 116934 106050 116986
rect 106102 116934 106114 116986
rect 106166 116934 106178 116986
rect 106230 116934 108836 116986
rect 104052 116912 108836 116934
rect 1104 116442 7912 116464
rect 1104 116390 4874 116442
rect 4926 116390 4938 116442
rect 4990 116390 5002 116442
rect 5054 116390 5066 116442
rect 5118 116390 5130 116442
rect 5182 116390 7912 116442
rect 1104 116368 7912 116390
rect 104052 116442 108836 116464
rect 104052 116390 106658 116442
rect 106710 116390 106722 116442
rect 106774 116390 106786 116442
rect 106838 116390 106850 116442
rect 106902 116390 106914 116442
rect 106966 116390 108836 116442
rect 104052 116368 108836 116390
rect 1104 115898 7912 115920
rect 1104 115846 4214 115898
rect 4266 115846 4278 115898
rect 4330 115846 4342 115898
rect 4394 115846 4406 115898
rect 4458 115846 4470 115898
rect 4522 115846 7912 115898
rect 1104 115824 7912 115846
rect 104052 115898 108836 115920
rect 104052 115846 105922 115898
rect 105974 115846 105986 115898
rect 106038 115846 106050 115898
rect 106102 115846 106114 115898
rect 106166 115846 106178 115898
rect 106230 115846 108836 115898
rect 104052 115824 108836 115846
rect 1104 115354 7912 115376
rect 1104 115302 4874 115354
rect 4926 115302 4938 115354
rect 4990 115302 5002 115354
rect 5054 115302 5066 115354
rect 5118 115302 5130 115354
rect 5182 115302 7912 115354
rect 1104 115280 7912 115302
rect 104052 115354 108836 115376
rect 104052 115302 106658 115354
rect 106710 115302 106722 115354
rect 106774 115302 106786 115354
rect 106838 115302 106850 115354
rect 106902 115302 106914 115354
rect 106966 115302 108836 115354
rect 104052 115280 108836 115302
rect 1104 114810 7912 114832
rect 1104 114758 4214 114810
rect 4266 114758 4278 114810
rect 4330 114758 4342 114810
rect 4394 114758 4406 114810
rect 4458 114758 4470 114810
rect 4522 114758 7912 114810
rect 1104 114736 7912 114758
rect 104052 114810 108836 114832
rect 104052 114758 105922 114810
rect 105974 114758 105986 114810
rect 106038 114758 106050 114810
rect 106102 114758 106114 114810
rect 106166 114758 106178 114810
rect 106230 114758 108836 114810
rect 104052 114736 108836 114758
rect 1104 114266 7912 114288
rect 1104 114214 4874 114266
rect 4926 114214 4938 114266
rect 4990 114214 5002 114266
rect 5054 114214 5066 114266
rect 5118 114214 5130 114266
rect 5182 114214 7912 114266
rect 1104 114192 7912 114214
rect 104052 114266 108836 114288
rect 104052 114214 106658 114266
rect 106710 114214 106722 114266
rect 106774 114214 106786 114266
rect 106838 114214 106850 114266
rect 106902 114214 106914 114266
rect 106966 114214 108836 114266
rect 104052 114192 108836 114214
rect 1104 113722 7912 113744
rect 1104 113670 4214 113722
rect 4266 113670 4278 113722
rect 4330 113670 4342 113722
rect 4394 113670 4406 113722
rect 4458 113670 4470 113722
rect 4522 113670 7912 113722
rect 1104 113648 7912 113670
rect 104052 113722 108836 113744
rect 104052 113670 105922 113722
rect 105974 113670 105986 113722
rect 106038 113670 106050 113722
rect 106102 113670 106114 113722
rect 106166 113670 106178 113722
rect 106230 113670 108836 113722
rect 104052 113648 108836 113670
rect 1104 113178 7912 113200
rect 1104 113126 4874 113178
rect 4926 113126 4938 113178
rect 4990 113126 5002 113178
rect 5054 113126 5066 113178
rect 5118 113126 5130 113178
rect 5182 113126 7912 113178
rect 1104 113104 7912 113126
rect 104052 113178 108836 113200
rect 104052 113126 106658 113178
rect 106710 113126 106722 113178
rect 106774 113126 106786 113178
rect 106838 113126 106850 113178
rect 106902 113126 106914 113178
rect 106966 113126 108836 113178
rect 104052 113104 108836 113126
rect 1104 112634 7912 112656
rect 1104 112582 4214 112634
rect 4266 112582 4278 112634
rect 4330 112582 4342 112634
rect 4394 112582 4406 112634
rect 4458 112582 4470 112634
rect 4522 112582 7912 112634
rect 1104 112560 7912 112582
rect 104052 112634 108836 112656
rect 104052 112582 105922 112634
rect 105974 112582 105986 112634
rect 106038 112582 106050 112634
rect 106102 112582 106114 112634
rect 106166 112582 106178 112634
rect 106230 112582 108836 112634
rect 104052 112560 108836 112582
rect 1104 112090 7912 112112
rect 1104 112038 4874 112090
rect 4926 112038 4938 112090
rect 4990 112038 5002 112090
rect 5054 112038 5066 112090
rect 5118 112038 5130 112090
rect 5182 112038 7912 112090
rect 1104 112016 7912 112038
rect 104052 112090 108836 112112
rect 104052 112038 106658 112090
rect 106710 112038 106722 112090
rect 106774 112038 106786 112090
rect 106838 112038 106850 112090
rect 106902 112038 106914 112090
rect 106966 112038 108836 112090
rect 104052 112016 108836 112038
rect 1104 111546 7912 111568
rect 1104 111494 4214 111546
rect 4266 111494 4278 111546
rect 4330 111494 4342 111546
rect 4394 111494 4406 111546
rect 4458 111494 4470 111546
rect 4522 111494 7912 111546
rect 1104 111472 7912 111494
rect 104052 111546 108836 111568
rect 104052 111494 105922 111546
rect 105974 111494 105986 111546
rect 106038 111494 106050 111546
rect 106102 111494 106114 111546
rect 106166 111494 106178 111546
rect 106230 111494 108836 111546
rect 104052 111472 108836 111494
rect 1581 111367 1639 111373
rect 1581 111333 1593 111367
rect 1627 111364 1639 111367
rect 8386 111364 8392 111376
rect 1627 111336 8392 111364
rect 1627 111333 1639 111336
rect 1581 111327 1639 111333
rect 8386 111324 8392 111336
rect 8444 111324 8450 111376
rect 1302 111188 1308 111240
rect 1360 111228 1366 111240
rect 1397 111231 1455 111237
rect 1397 111228 1409 111231
rect 1360 111200 1409 111228
rect 1360 111188 1366 111200
rect 1397 111197 1409 111200
rect 1443 111228 1455 111231
rect 1673 111231 1731 111237
rect 1673 111228 1685 111231
rect 1443 111200 1685 111228
rect 1443 111197 1455 111200
rect 1397 111191 1455 111197
rect 1673 111197 1685 111200
rect 1719 111197 1731 111231
rect 1673 111191 1731 111197
rect 1104 111002 7912 111024
rect 1104 110950 4874 111002
rect 4926 110950 4938 111002
rect 4990 110950 5002 111002
rect 5054 110950 5066 111002
rect 5118 110950 5130 111002
rect 5182 110950 7912 111002
rect 1104 110928 7912 110950
rect 104052 111002 108836 111024
rect 104052 110950 106658 111002
rect 106710 110950 106722 111002
rect 106774 110950 106786 111002
rect 106838 110950 106850 111002
rect 106902 110950 106914 111002
rect 106966 110950 108836 111002
rect 104052 110928 108836 110950
rect 1104 110458 7912 110480
rect 1104 110406 4214 110458
rect 4266 110406 4278 110458
rect 4330 110406 4342 110458
rect 4394 110406 4406 110458
rect 4458 110406 4470 110458
rect 4522 110406 7912 110458
rect 1104 110384 7912 110406
rect 104052 110458 108836 110480
rect 104052 110406 105922 110458
rect 105974 110406 105986 110458
rect 106038 110406 106050 110458
rect 106102 110406 106114 110458
rect 106166 110406 106178 110458
rect 106230 110406 108836 110458
rect 104052 110384 108836 110406
rect 1104 109914 7912 109936
rect 1104 109862 4874 109914
rect 4926 109862 4938 109914
rect 4990 109862 5002 109914
rect 5054 109862 5066 109914
rect 5118 109862 5130 109914
rect 5182 109862 7912 109914
rect 1104 109840 7912 109862
rect 104052 109914 108836 109936
rect 104052 109862 106658 109914
rect 106710 109862 106722 109914
rect 106774 109862 106786 109914
rect 106838 109862 106850 109914
rect 106902 109862 106914 109914
rect 106966 109862 108836 109914
rect 104052 109840 108836 109862
rect 1302 109624 1308 109676
rect 1360 109664 1366 109676
rect 1397 109667 1455 109673
rect 1397 109664 1409 109667
rect 1360 109636 1409 109664
rect 1360 109624 1366 109636
rect 1397 109633 1409 109636
rect 1443 109664 1455 109667
rect 1673 109667 1731 109673
rect 1673 109664 1685 109667
rect 1443 109636 1685 109664
rect 1443 109633 1455 109636
rect 1397 109627 1455 109633
rect 1673 109633 1685 109636
rect 1719 109633 1731 109667
rect 1673 109627 1731 109633
rect 1581 109531 1639 109537
rect 1581 109497 1593 109531
rect 1627 109528 1639 109531
rect 8386 109528 8392 109540
rect 1627 109500 8392 109528
rect 1627 109497 1639 109500
rect 1581 109491 1639 109497
rect 8386 109488 8392 109500
rect 8444 109488 8450 109540
rect 1104 109370 7912 109392
rect 1104 109318 4214 109370
rect 4266 109318 4278 109370
rect 4330 109318 4342 109370
rect 4394 109318 4406 109370
rect 4458 109318 4470 109370
rect 4522 109318 7912 109370
rect 1104 109296 7912 109318
rect 104052 109370 108836 109392
rect 104052 109318 105922 109370
rect 105974 109318 105986 109370
rect 106038 109318 106050 109370
rect 106102 109318 106114 109370
rect 106166 109318 106178 109370
rect 106230 109318 108836 109370
rect 104052 109296 108836 109318
rect 1104 108826 7912 108848
rect 1104 108774 4874 108826
rect 4926 108774 4938 108826
rect 4990 108774 5002 108826
rect 5054 108774 5066 108826
rect 5118 108774 5130 108826
rect 5182 108774 7912 108826
rect 1104 108752 7912 108774
rect 104052 108826 108836 108848
rect 104052 108774 106658 108826
rect 106710 108774 106722 108826
rect 106774 108774 106786 108826
rect 106838 108774 106850 108826
rect 106902 108774 106914 108826
rect 106966 108774 108836 108826
rect 104052 108752 108836 108774
rect 1302 108536 1308 108588
rect 1360 108576 1366 108588
rect 1397 108579 1455 108585
rect 1397 108576 1409 108579
rect 1360 108548 1409 108576
rect 1360 108536 1366 108548
rect 1397 108545 1409 108548
rect 1443 108576 1455 108579
rect 1673 108579 1731 108585
rect 1673 108576 1685 108579
rect 1443 108548 1685 108576
rect 1443 108545 1455 108548
rect 1397 108539 1455 108545
rect 1673 108545 1685 108548
rect 1719 108545 1731 108579
rect 1673 108539 1731 108545
rect 1581 108443 1639 108449
rect 1581 108409 1593 108443
rect 1627 108440 1639 108443
rect 8386 108440 8392 108452
rect 1627 108412 8392 108440
rect 1627 108409 1639 108412
rect 1581 108403 1639 108409
rect 8386 108400 8392 108412
rect 8444 108400 8450 108452
rect 1104 108282 7912 108304
rect 1104 108230 4214 108282
rect 4266 108230 4278 108282
rect 4330 108230 4342 108282
rect 4394 108230 4406 108282
rect 4458 108230 4470 108282
rect 4522 108230 7912 108282
rect 1104 108208 7912 108230
rect 104052 108282 108836 108304
rect 104052 108230 105922 108282
rect 105974 108230 105986 108282
rect 106038 108230 106050 108282
rect 106102 108230 106114 108282
rect 106166 108230 106178 108282
rect 106230 108230 108836 108282
rect 104052 108208 108836 108230
rect 1104 107738 7912 107760
rect 1104 107686 4874 107738
rect 4926 107686 4938 107738
rect 4990 107686 5002 107738
rect 5054 107686 5066 107738
rect 5118 107686 5130 107738
rect 5182 107686 7912 107738
rect 1104 107664 7912 107686
rect 104052 107738 108836 107760
rect 104052 107686 106658 107738
rect 106710 107686 106722 107738
rect 106774 107686 106786 107738
rect 106838 107686 106850 107738
rect 106902 107686 106914 107738
rect 106966 107686 108836 107738
rect 104052 107664 108836 107686
rect 1104 107194 7912 107216
rect 1104 107142 4214 107194
rect 4266 107142 4278 107194
rect 4330 107142 4342 107194
rect 4394 107142 4406 107194
rect 4458 107142 4470 107194
rect 4522 107142 7912 107194
rect 1104 107120 7912 107142
rect 104052 107194 108836 107216
rect 104052 107142 105922 107194
rect 105974 107142 105986 107194
rect 106038 107142 106050 107194
rect 106102 107142 106114 107194
rect 106166 107142 106178 107194
rect 106230 107142 108836 107194
rect 104052 107120 108836 107142
rect 1581 107015 1639 107021
rect 1581 106981 1593 107015
rect 1627 107012 1639 107015
rect 8386 107012 8392 107024
rect 1627 106984 8392 107012
rect 1627 106981 1639 106984
rect 1581 106975 1639 106981
rect 8386 106972 8392 106984
rect 8444 106972 8450 107024
rect 1210 106836 1216 106888
rect 1268 106876 1274 106888
rect 1397 106879 1455 106885
rect 1397 106876 1409 106879
rect 1268 106848 1409 106876
rect 1268 106836 1274 106848
rect 1397 106845 1409 106848
rect 1443 106876 1455 106879
rect 1673 106879 1731 106885
rect 1673 106876 1685 106879
rect 1443 106848 1685 106876
rect 1443 106845 1455 106848
rect 1397 106839 1455 106845
rect 1673 106845 1685 106848
rect 1719 106845 1731 106879
rect 1673 106839 1731 106845
rect 1104 106650 7912 106672
rect 1104 106598 4874 106650
rect 4926 106598 4938 106650
rect 4990 106598 5002 106650
rect 5054 106598 5066 106650
rect 5118 106598 5130 106650
rect 5182 106598 7912 106650
rect 1104 106576 7912 106598
rect 104052 106650 108836 106672
rect 104052 106598 106658 106650
rect 106710 106598 106722 106650
rect 106774 106598 106786 106650
rect 106838 106598 106850 106650
rect 106902 106598 106914 106650
rect 106966 106598 108836 106650
rect 104052 106576 108836 106598
rect 1104 106106 7912 106128
rect 1104 106054 4214 106106
rect 4266 106054 4278 106106
rect 4330 106054 4342 106106
rect 4394 106054 4406 106106
rect 4458 106054 4470 106106
rect 4522 106054 7912 106106
rect 1104 106032 7912 106054
rect 104052 106106 108836 106128
rect 104052 106054 105922 106106
rect 105974 106054 105986 106106
rect 106038 106054 106050 106106
rect 106102 106054 106114 106106
rect 106166 106054 106178 106106
rect 106230 106054 108836 106106
rect 104052 106032 108836 106054
rect 1581 105927 1639 105933
rect 1581 105893 1593 105927
rect 1627 105924 1639 105927
rect 8386 105924 8392 105936
rect 1627 105896 8392 105924
rect 1627 105893 1639 105896
rect 1581 105887 1639 105893
rect 8386 105884 8392 105896
rect 8444 105884 8450 105936
rect 1302 105748 1308 105800
rect 1360 105788 1366 105800
rect 1397 105791 1455 105797
rect 1397 105788 1409 105791
rect 1360 105760 1409 105788
rect 1360 105748 1366 105760
rect 1397 105757 1409 105760
rect 1443 105788 1455 105791
rect 1673 105791 1731 105797
rect 1673 105788 1685 105791
rect 1443 105760 1685 105788
rect 1443 105757 1455 105760
rect 1397 105751 1455 105757
rect 1673 105757 1685 105760
rect 1719 105757 1731 105791
rect 1673 105751 1731 105757
rect 1104 105562 7912 105584
rect 1104 105510 4874 105562
rect 4926 105510 4938 105562
rect 4990 105510 5002 105562
rect 5054 105510 5066 105562
rect 5118 105510 5130 105562
rect 5182 105510 7912 105562
rect 1104 105488 7912 105510
rect 104052 105562 108836 105584
rect 104052 105510 106658 105562
rect 106710 105510 106722 105562
rect 106774 105510 106786 105562
rect 106838 105510 106850 105562
rect 106902 105510 106914 105562
rect 106966 105510 108836 105562
rect 104052 105488 108836 105510
rect 1104 105018 7912 105040
rect 1104 104966 4214 105018
rect 4266 104966 4278 105018
rect 4330 104966 4342 105018
rect 4394 104966 4406 105018
rect 4458 104966 4470 105018
rect 4522 104966 7912 105018
rect 1104 104944 7912 104966
rect 104052 105018 108836 105040
rect 104052 104966 105922 105018
rect 105974 104966 105986 105018
rect 106038 104966 106050 105018
rect 106102 104966 106114 105018
rect 106166 104966 106178 105018
rect 106230 104966 108836 105018
rect 104052 104944 108836 104966
rect 1104 104474 7912 104496
rect 1104 104422 4874 104474
rect 4926 104422 4938 104474
rect 4990 104422 5002 104474
rect 5054 104422 5066 104474
rect 5118 104422 5130 104474
rect 5182 104422 7912 104474
rect 1104 104400 7912 104422
rect 104052 104474 108836 104496
rect 104052 104422 106658 104474
rect 106710 104422 106722 104474
rect 106774 104422 106786 104474
rect 106838 104422 106850 104474
rect 106902 104422 106914 104474
rect 106966 104422 108836 104474
rect 104052 104400 108836 104422
rect 1302 104184 1308 104236
rect 1360 104224 1366 104236
rect 1397 104227 1455 104233
rect 1397 104224 1409 104227
rect 1360 104196 1409 104224
rect 1360 104184 1366 104196
rect 1397 104193 1409 104196
rect 1443 104224 1455 104227
rect 1673 104227 1731 104233
rect 1673 104224 1685 104227
rect 1443 104196 1685 104224
rect 1443 104193 1455 104196
rect 1397 104187 1455 104193
rect 1673 104193 1685 104196
rect 1719 104193 1731 104227
rect 1673 104187 1731 104193
rect 1581 104091 1639 104097
rect 1581 104057 1593 104091
rect 1627 104088 1639 104091
rect 8386 104088 8392 104100
rect 1627 104060 8392 104088
rect 1627 104057 1639 104060
rect 1581 104051 1639 104057
rect 8386 104048 8392 104060
rect 8444 104048 8450 104100
rect 1104 103930 7912 103952
rect 1104 103878 4214 103930
rect 4266 103878 4278 103930
rect 4330 103878 4342 103930
rect 4394 103878 4406 103930
rect 4458 103878 4470 103930
rect 4522 103878 7912 103930
rect 1104 103856 7912 103878
rect 104052 103930 108836 103952
rect 104052 103878 105922 103930
rect 105974 103878 105986 103930
rect 106038 103878 106050 103930
rect 106102 103878 106114 103930
rect 106166 103878 106178 103930
rect 106230 103878 108836 103930
rect 104052 103856 108836 103878
rect 1104 103386 7912 103408
rect 1104 103334 4874 103386
rect 4926 103334 4938 103386
rect 4990 103334 5002 103386
rect 5054 103334 5066 103386
rect 5118 103334 5130 103386
rect 5182 103334 7912 103386
rect 1104 103312 7912 103334
rect 104052 103386 108836 103408
rect 104052 103334 106658 103386
rect 106710 103334 106722 103386
rect 106774 103334 106786 103386
rect 106838 103334 106850 103386
rect 106902 103334 106914 103386
rect 106966 103334 108836 103386
rect 104052 103312 108836 103334
rect 1104 102842 7912 102864
rect 1104 102790 4214 102842
rect 4266 102790 4278 102842
rect 4330 102790 4342 102842
rect 4394 102790 4406 102842
rect 4458 102790 4470 102842
rect 4522 102790 7912 102842
rect 1104 102768 7912 102790
rect 104052 102842 108836 102864
rect 104052 102790 105922 102842
rect 105974 102790 105986 102842
rect 106038 102790 106050 102842
rect 106102 102790 106114 102842
rect 106166 102790 106178 102842
rect 106230 102790 108836 102842
rect 104052 102768 108836 102790
rect 1104 102298 7912 102320
rect 1104 102246 4874 102298
rect 4926 102246 4938 102298
rect 4990 102246 5002 102298
rect 5054 102246 5066 102298
rect 5118 102246 5130 102298
rect 5182 102246 7912 102298
rect 1104 102224 7912 102246
rect 104052 102298 108836 102320
rect 104052 102246 106658 102298
rect 106710 102246 106722 102298
rect 106774 102246 106786 102298
rect 106838 102246 106850 102298
rect 106902 102246 106914 102298
rect 106966 102246 108836 102298
rect 104052 102224 108836 102246
rect 1104 101754 7912 101776
rect 1104 101702 4214 101754
rect 4266 101702 4278 101754
rect 4330 101702 4342 101754
rect 4394 101702 4406 101754
rect 4458 101702 4470 101754
rect 4522 101702 7912 101754
rect 1104 101680 7912 101702
rect 104052 101754 108836 101776
rect 104052 101702 105922 101754
rect 105974 101702 105986 101754
rect 106038 101702 106050 101754
rect 106102 101702 106114 101754
rect 106166 101702 106178 101754
rect 106230 101702 108836 101754
rect 104052 101680 108836 101702
rect 1104 101210 7912 101232
rect 1104 101158 4874 101210
rect 4926 101158 4938 101210
rect 4990 101158 5002 101210
rect 5054 101158 5066 101210
rect 5118 101158 5130 101210
rect 5182 101158 7912 101210
rect 1104 101136 7912 101158
rect 104052 101210 108836 101232
rect 104052 101158 106658 101210
rect 106710 101158 106722 101210
rect 106774 101158 106786 101210
rect 106838 101158 106850 101210
rect 106902 101158 106914 101210
rect 106966 101158 108836 101210
rect 104052 101136 108836 101158
rect 1104 100666 7912 100688
rect 1104 100614 4214 100666
rect 4266 100614 4278 100666
rect 4330 100614 4342 100666
rect 4394 100614 4406 100666
rect 4458 100614 4470 100666
rect 4522 100614 7912 100666
rect 1104 100592 7912 100614
rect 104052 100666 108836 100688
rect 104052 100614 105922 100666
rect 105974 100614 105986 100666
rect 106038 100614 106050 100666
rect 106102 100614 106114 100666
rect 106166 100614 106178 100666
rect 106230 100614 108836 100666
rect 104052 100592 108836 100614
rect 1104 100122 7912 100144
rect 1104 100070 4874 100122
rect 4926 100070 4938 100122
rect 4990 100070 5002 100122
rect 5054 100070 5066 100122
rect 5118 100070 5130 100122
rect 5182 100070 7912 100122
rect 1104 100048 7912 100070
rect 104052 100122 108836 100144
rect 104052 100070 106658 100122
rect 106710 100070 106722 100122
rect 106774 100070 106786 100122
rect 106838 100070 106850 100122
rect 106902 100070 106914 100122
rect 106966 100070 108836 100122
rect 104052 100048 108836 100070
rect 1104 99578 7912 99600
rect 1104 99526 4214 99578
rect 4266 99526 4278 99578
rect 4330 99526 4342 99578
rect 4394 99526 4406 99578
rect 4458 99526 4470 99578
rect 4522 99526 7912 99578
rect 1104 99504 7912 99526
rect 104052 99578 108836 99600
rect 104052 99526 105922 99578
rect 105974 99526 105986 99578
rect 106038 99526 106050 99578
rect 106102 99526 106114 99578
rect 106166 99526 106178 99578
rect 106230 99526 108836 99578
rect 104052 99504 108836 99526
rect 1104 99034 7912 99056
rect 1104 98982 4874 99034
rect 4926 98982 4938 99034
rect 4990 98982 5002 99034
rect 5054 98982 5066 99034
rect 5118 98982 5130 99034
rect 5182 98982 7912 99034
rect 1104 98960 7912 98982
rect 104052 99034 108836 99056
rect 104052 98982 106658 99034
rect 106710 98982 106722 99034
rect 106774 98982 106786 99034
rect 106838 98982 106850 99034
rect 106902 98982 106914 99034
rect 106966 98982 108836 99034
rect 104052 98960 108836 98982
rect 1104 98490 7912 98512
rect 1104 98438 4214 98490
rect 4266 98438 4278 98490
rect 4330 98438 4342 98490
rect 4394 98438 4406 98490
rect 4458 98438 4470 98490
rect 4522 98438 7912 98490
rect 1104 98416 7912 98438
rect 104052 98490 108836 98512
rect 104052 98438 105922 98490
rect 105974 98438 105986 98490
rect 106038 98438 106050 98490
rect 106102 98438 106114 98490
rect 106166 98438 106178 98490
rect 106230 98438 108836 98490
rect 104052 98416 108836 98438
rect 1104 97946 7912 97968
rect 1104 97894 4874 97946
rect 4926 97894 4938 97946
rect 4990 97894 5002 97946
rect 5054 97894 5066 97946
rect 5118 97894 5130 97946
rect 5182 97894 7912 97946
rect 1104 97872 7912 97894
rect 104052 97946 108836 97968
rect 104052 97894 106658 97946
rect 106710 97894 106722 97946
rect 106774 97894 106786 97946
rect 106838 97894 106850 97946
rect 106902 97894 106914 97946
rect 106966 97894 108836 97946
rect 104052 97872 108836 97894
rect 1104 97402 7912 97424
rect 1104 97350 4214 97402
rect 4266 97350 4278 97402
rect 4330 97350 4342 97402
rect 4394 97350 4406 97402
rect 4458 97350 4470 97402
rect 4522 97350 7912 97402
rect 1104 97328 7912 97350
rect 104052 97402 108836 97424
rect 104052 97350 105922 97402
rect 105974 97350 105986 97402
rect 106038 97350 106050 97402
rect 106102 97350 106114 97402
rect 106166 97350 106178 97402
rect 106230 97350 108836 97402
rect 104052 97328 108836 97350
rect 1104 96858 7912 96880
rect 1104 96806 4874 96858
rect 4926 96806 4938 96858
rect 4990 96806 5002 96858
rect 5054 96806 5066 96858
rect 5118 96806 5130 96858
rect 5182 96806 7912 96858
rect 1104 96784 7912 96806
rect 104052 96858 108836 96880
rect 104052 96806 106658 96858
rect 106710 96806 106722 96858
rect 106774 96806 106786 96858
rect 106838 96806 106850 96858
rect 106902 96806 106914 96858
rect 106966 96806 108836 96858
rect 104052 96784 108836 96806
rect 1104 96314 7912 96336
rect 1104 96262 4214 96314
rect 4266 96262 4278 96314
rect 4330 96262 4342 96314
rect 4394 96262 4406 96314
rect 4458 96262 4470 96314
rect 4522 96262 7912 96314
rect 1104 96240 7912 96262
rect 104052 96314 108836 96336
rect 104052 96262 105922 96314
rect 105974 96262 105986 96314
rect 106038 96262 106050 96314
rect 106102 96262 106114 96314
rect 106166 96262 106178 96314
rect 106230 96262 108836 96314
rect 104052 96240 108836 96262
rect 1104 95770 7912 95792
rect 1104 95718 4874 95770
rect 4926 95718 4938 95770
rect 4990 95718 5002 95770
rect 5054 95718 5066 95770
rect 5118 95718 5130 95770
rect 5182 95718 7912 95770
rect 1104 95696 7912 95718
rect 104052 95770 108836 95792
rect 104052 95718 106658 95770
rect 106710 95718 106722 95770
rect 106774 95718 106786 95770
rect 106838 95718 106850 95770
rect 106902 95718 106914 95770
rect 106966 95718 108836 95770
rect 104052 95696 108836 95718
rect 102686 95276 102692 95328
rect 102744 95316 102750 95328
rect 104345 95319 104403 95325
rect 104345 95316 104357 95319
rect 102744 95288 104357 95316
rect 102744 95276 102750 95288
rect 104345 95285 104357 95288
rect 104391 95285 104403 95319
rect 104345 95279 104403 95285
rect 1104 95226 7912 95248
rect 1104 95174 4214 95226
rect 4266 95174 4278 95226
rect 4330 95174 4342 95226
rect 4394 95174 4406 95226
rect 4458 95174 4470 95226
rect 4522 95174 7912 95226
rect 1104 95152 7912 95174
rect 104052 95226 108836 95248
rect 104052 95174 105922 95226
rect 105974 95174 105986 95226
rect 106038 95174 106050 95226
rect 106102 95174 106114 95226
rect 106166 95174 106178 95226
rect 106230 95174 108836 95226
rect 104052 95152 108836 95174
rect 1104 94682 7912 94704
rect 1104 94630 4874 94682
rect 4926 94630 4938 94682
rect 4990 94630 5002 94682
rect 5054 94630 5066 94682
rect 5118 94630 5130 94682
rect 5182 94630 7912 94682
rect 1104 94608 7912 94630
rect 104052 94682 108836 94704
rect 104052 94630 106658 94682
rect 106710 94630 106722 94682
rect 106774 94630 106786 94682
rect 106838 94630 106850 94682
rect 106902 94630 106914 94682
rect 106966 94630 108836 94682
rect 104052 94608 108836 94630
rect 1104 94138 7912 94160
rect 1104 94086 4214 94138
rect 4266 94086 4278 94138
rect 4330 94086 4342 94138
rect 4394 94086 4406 94138
rect 4458 94086 4470 94138
rect 4522 94086 7912 94138
rect 1104 94064 7912 94086
rect 104052 94138 108836 94160
rect 104052 94086 105922 94138
rect 105974 94086 105986 94138
rect 106038 94086 106050 94138
rect 106102 94086 106114 94138
rect 106166 94086 106178 94138
rect 106230 94086 108836 94138
rect 104052 94064 108836 94086
rect 103054 93848 103060 93900
rect 103112 93888 103118 93900
rect 104345 93891 104403 93897
rect 104345 93888 104357 93891
rect 103112 93860 104357 93888
rect 103112 93848 103118 93860
rect 104345 93857 104357 93860
rect 104391 93857 104403 93891
rect 104345 93851 104403 93857
rect 1104 93594 7912 93616
rect 1104 93542 4874 93594
rect 4926 93542 4938 93594
rect 4990 93542 5002 93594
rect 5054 93542 5066 93594
rect 5118 93542 5130 93594
rect 5182 93542 7912 93594
rect 1104 93520 7912 93542
rect 104052 93594 108836 93616
rect 104052 93542 106658 93594
rect 106710 93542 106722 93594
rect 106774 93542 106786 93594
rect 106838 93542 106850 93594
rect 106902 93542 106914 93594
rect 106966 93542 108836 93594
rect 104052 93520 108836 93542
rect 1104 93050 7912 93072
rect 1104 92998 4214 93050
rect 4266 92998 4278 93050
rect 4330 92998 4342 93050
rect 4394 92998 4406 93050
rect 4458 92998 4470 93050
rect 4522 92998 7912 93050
rect 1104 92976 7912 92998
rect 104052 93050 108836 93072
rect 104052 92998 105922 93050
rect 105974 92998 105986 93050
rect 106038 92998 106050 93050
rect 106102 92998 106114 93050
rect 106166 92998 106178 93050
rect 106230 92998 108836 93050
rect 104052 92976 108836 92998
rect 102962 92556 102968 92608
rect 103020 92596 103026 92608
rect 104345 92599 104403 92605
rect 104345 92596 104357 92599
rect 103020 92568 104357 92596
rect 103020 92556 103026 92568
rect 104345 92565 104357 92568
rect 104391 92565 104403 92599
rect 104345 92559 104403 92565
rect 1104 92506 7912 92528
rect 1104 92454 4874 92506
rect 4926 92454 4938 92506
rect 4990 92454 5002 92506
rect 5054 92454 5066 92506
rect 5118 92454 5130 92506
rect 5182 92454 7912 92506
rect 1104 92432 7912 92454
rect 104052 92506 108836 92528
rect 104052 92454 106658 92506
rect 106710 92454 106722 92506
rect 106774 92454 106786 92506
rect 106838 92454 106850 92506
rect 106902 92454 106914 92506
rect 106966 92454 108836 92506
rect 104052 92432 108836 92454
rect 1104 91962 7912 91984
rect 1104 91910 4214 91962
rect 4266 91910 4278 91962
rect 4330 91910 4342 91962
rect 4394 91910 4406 91962
rect 4458 91910 4470 91962
rect 4522 91910 7912 91962
rect 1104 91888 7912 91910
rect 104052 91962 108836 91984
rect 104052 91910 105922 91962
rect 105974 91910 105986 91962
rect 106038 91910 106050 91962
rect 106102 91910 106114 91962
rect 106166 91910 106178 91962
rect 106230 91910 108836 91962
rect 104052 91888 108836 91910
rect 1104 91418 7912 91440
rect 1104 91366 4874 91418
rect 4926 91366 4938 91418
rect 4990 91366 5002 91418
rect 5054 91366 5066 91418
rect 5118 91366 5130 91418
rect 5182 91366 7912 91418
rect 1104 91344 7912 91366
rect 104052 91418 108836 91440
rect 104052 91366 106658 91418
rect 106710 91366 106722 91418
rect 106774 91366 106786 91418
rect 106838 91366 106850 91418
rect 106902 91366 106914 91418
rect 106966 91366 108836 91418
rect 104052 91344 108836 91366
rect 104342 91128 104348 91180
rect 104400 91128 104406 91180
rect 103514 90924 103520 90976
rect 103572 90964 103578 90976
rect 104158 90964 104164 90976
rect 103572 90936 104164 90964
rect 103572 90924 103578 90936
rect 104158 90924 104164 90936
rect 104216 90964 104222 90976
rect 105633 90967 105691 90973
rect 105633 90964 105645 90967
rect 104216 90936 105645 90964
rect 104216 90924 104222 90936
rect 105633 90933 105645 90936
rect 105679 90964 105691 90967
rect 106185 90967 106243 90973
rect 106185 90964 106197 90967
rect 105679 90936 106197 90964
rect 105679 90933 105691 90936
rect 105633 90927 105691 90933
rect 106185 90933 106197 90936
rect 106231 90933 106243 90967
rect 106185 90927 106243 90933
rect 1104 90874 7912 90896
rect 1104 90822 4214 90874
rect 4266 90822 4278 90874
rect 4330 90822 4342 90874
rect 4394 90822 4406 90874
rect 4458 90822 4470 90874
rect 4522 90822 7912 90874
rect 1104 90800 7912 90822
rect 104052 90874 108836 90896
rect 104052 90822 105922 90874
rect 105974 90822 105986 90874
rect 106038 90822 106050 90874
rect 106102 90822 106114 90874
rect 106166 90822 106178 90874
rect 106230 90822 108836 90874
rect 104052 90800 108836 90822
rect 104342 90380 104348 90432
rect 104400 90380 104406 90432
rect 1104 90330 7912 90352
rect 1104 90278 4874 90330
rect 4926 90278 4938 90330
rect 4990 90278 5002 90330
rect 5054 90278 5066 90330
rect 5118 90278 5130 90330
rect 5182 90278 7912 90330
rect 1104 90256 7912 90278
rect 104052 90330 108836 90352
rect 104052 90278 106658 90330
rect 106710 90278 106722 90330
rect 106774 90278 106786 90330
rect 106838 90278 106850 90330
rect 106902 90278 106914 90330
rect 106966 90278 108836 90330
rect 104052 90256 108836 90278
rect 1104 89786 7912 89808
rect 1104 89734 4214 89786
rect 4266 89734 4278 89786
rect 4330 89734 4342 89786
rect 4394 89734 4406 89786
rect 4458 89734 4470 89786
rect 4522 89734 7912 89786
rect 1104 89712 7912 89734
rect 104052 89786 108836 89808
rect 104052 89734 105922 89786
rect 105974 89734 105986 89786
rect 106038 89734 106050 89786
rect 106102 89734 106114 89786
rect 106166 89734 106178 89786
rect 106230 89734 108836 89786
rect 104052 89712 108836 89734
rect 1104 89242 7912 89264
rect 1104 89190 4874 89242
rect 4926 89190 4938 89242
rect 4990 89190 5002 89242
rect 5054 89190 5066 89242
rect 5118 89190 5130 89242
rect 5182 89190 7912 89242
rect 1104 89168 7912 89190
rect 104052 89242 108836 89264
rect 104052 89190 106658 89242
rect 106710 89190 106722 89242
rect 106774 89190 106786 89242
rect 106838 89190 106850 89242
rect 106902 89190 106914 89242
rect 106966 89190 108836 89242
rect 104052 89168 108836 89190
rect 1302 88952 1308 89004
rect 1360 88992 1366 89004
rect 1489 88995 1547 89001
rect 1489 88992 1501 88995
rect 1360 88964 1501 88992
rect 1360 88952 1366 88964
rect 1489 88961 1501 88964
rect 1535 88992 1547 88995
rect 1949 88995 2007 89001
rect 1949 88992 1961 88995
rect 1535 88964 1961 88992
rect 1535 88961 1547 88964
rect 1489 88955 1547 88961
rect 1949 88961 1961 88964
rect 1995 88961 2007 88995
rect 1949 88955 2007 88961
rect 1673 88859 1731 88865
rect 1673 88825 1685 88859
rect 1719 88856 1731 88859
rect 1857 88859 1915 88865
rect 1857 88856 1869 88859
rect 1719 88828 1869 88856
rect 1719 88825 1731 88828
rect 1673 88819 1731 88825
rect 1857 88825 1869 88828
rect 1903 88856 1915 88859
rect 7558 88856 7564 88868
rect 1903 88828 7564 88856
rect 1903 88825 1915 88828
rect 1857 88819 1915 88825
rect 7558 88816 7564 88828
rect 7616 88816 7622 88868
rect 1104 88698 7912 88720
rect 1104 88646 4214 88698
rect 4266 88646 4278 88698
rect 4330 88646 4342 88698
rect 4394 88646 4406 88698
rect 4458 88646 4470 88698
rect 4522 88646 7912 88698
rect 1104 88624 7912 88646
rect 104052 88698 108836 88720
rect 104052 88646 105922 88698
rect 105974 88646 105986 88698
rect 106038 88646 106050 88698
rect 106102 88646 106114 88698
rect 106166 88646 106178 88698
rect 106230 88646 108836 88698
rect 104052 88624 108836 88646
rect 1104 88154 7912 88176
rect 1104 88102 4874 88154
rect 4926 88102 4938 88154
rect 4990 88102 5002 88154
rect 5054 88102 5066 88154
rect 5118 88102 5130 88154
rect 5182 88102 7912 88154
rect 1104 88080 7912 88102
rect 104052 88154 108836 88176
rect 104052 88102 106658 88154
rect 106710 88102 106722 88154
rect 106774 88102 106786 88154
rect 106838 88102 106850 88154
rect 106902 88102 106914 88154
rect 106966 88102 108836 88154
rect 104052 88080 108836 88102
rect 1210 87864 1216 87916
rect 1268 87904 1274 87916
rect 1489 87907 1547 87913
rect 1489 87904 1501 87907
rect 1268 87876 1501 87904
rect 1268 87864 1274 87876
rect 1489 87873 1501 87876
rect 1535 87904 1547 87907
rect 1949 87907 2007 87913
rect 1949 87904 1961 87907
rect 1535 87876 1961 87904
rect 1535 87873 1547 87876
rect 1489 87867 1547 87873
rect 1949 87873 1961 87876
rect 1995 87873 2007 87907
rect 1949 87867 2007 87873
rect 1673 87771 1731 87777
rect 1673 87737 1685 87771
rect 1719 87768 1731 87771
rect 1857 87771 1915 87777
rect 1857 87768 1869 87771
rect 1719 87740 1869 87768
rect 1719 87737 1731 87740
rect 1673 87731 1731 87737
rect 1857 87737 1869 87740
rect 1903 87768 1915 87771
rect 8938 87768 8944 87780
rect 1903 87740 8944 87768
rect 1903 87737 1915 87740
rect 1857 87731 1915 87737
rect 8938 87728 8944 87740
rect 8996 87728 9002 87780
rect 1104 87610 7912 87632
rect 1104 87558 4214 87610
rect 4266 87558 4278 87610
rect 4330 87558 4342 87610
rect 4394 87558 4406 87610
rect 4458 87558 4470 87610
rect 4522 87558 7912 87610
rect 1104 87536 7912 87558
rect 104052 87610 108836 87632
rect 104052 87558 105922 87610
rect 105974 87558 105986 87610
rect 106038 87558 106050 87610
rect 106102 87558 106114 87610
rect 106166 87558 106178 87610
rect 106230 87558 108836 87610
rect 104052 87536 108836 87558
rect 1210 87184 1216 87236
rect 1268 87224 1274 87236
rect 1489 87227 1547 87233
rect 1489 87224 1501 87227
rect 1268 87196 1501 87224
rect 1268 87184 1274 87196
rect 1489 87193 1501 87196
rect 1535 87224 1547 87227
rect 1949 87227 2007 87233
rect 1949 87224 1961 87227
rect 1535 87196 1961 87224
rect 1535 87193 1547 87196
rect 1489 87187 1547 87193
rect 1949 87193 1961 87196
rect 1995 87193 2007 87227
rect 1949 87187 2007 87193
rect 1581 87159 1639 87165
rect 1581 87125 1593 87159
rect 1627 87156 1639 87159
rect 1854 87156 1860 87168
rect 1627 87128 1860 87156
rect 1627 87125 1639 87128
rect 1581 87119 1639 87125
rect 1854 87116 1860 87128
rect 1912 87116 1918 87168
rect 1104 87066 7912 87088
rect 1104 87014 4874 87066
rect 4926 87014 4938 87066
rect 4990 87014 5002 87066
rect 5054 87014 5066 87066
rect 5118 87014 5130 87066
rect 5182 87014 7912 87066
rect 1104 86992 7912 87014
rect 104052 87066 108836 87088
rect 104052 87014 106658 87066
rect 106710 87014 106722 87066
rect 106774 87014 106786 87066
rect 106838 87014 106850 87066
rect 106902 87014 106914 87066
rect 106966 87014 108836 87066
rect 104052 86992 108836 87014
rect 1302 86776 1308 86828
rect 1360 86816 1366 86828
rect 1489 86819 1547 86825
rect 1489 86816 1501 86819
rect 1360 86788 1501 86816
rect 1360 86776 1366 86788
rect 1489 86785 1501 86788
rect 1535 86816 1547 86819
rect 1949 86819 2007 86825
rect 1949 86816 1961 86819
rect 1535 86788 1961 86816
rect 1535 86785 1547 86788
rect 1489 86779 1547 86785
rect 1949 86785 1961 86788
rect 1995 86785 2007 86819
rect 1949 86779 2007 86785
rect 1673 86683 1731 86689
rect 1673 86649 1685 86683
rect 1719 86680 1731 86683
rect 1857 86683 1915 86689
rect 1857 86680 1869 86683
rect 1719 86652 1869 86680
rect 1719 86649 1731 86652
rect 1673 86643 1731 86649
rect 1857 86649 1869 86652
rect 1903 86680 1915 86683
rect 8662 86680 8668 86692
rect 1903 86652 8668 86680
rect 1903 86649 1915 86652
rect 1857 86643 1915 86649
rect 8662 86640 8668 86652
rect 8720 86640 8726 86692
rect 1104 86522 7912 86544
rect 1104 86470 4214 86522
rect 4266 86470 4278 86522
rect 4330 86470 4342 86522
rect 4394 86470 4406 86522
rect 4458 86470 4470 86522
rect 4522 86470 7912 86522
rect 1104 86448 7912 86470
rect 104052 86522 108836 86544
rect 104052 86470 105922 86522
rect 105974 86470 105986 86522
rect 106038 86470 106050 86522
rect 106102 86470 106114 86522
rect 106166 86470 106178 86522
rect 106230 86470 108836 86522
rect 104052 86448 108836 86470
rect 1302 86164 1308 86216
rect 1360 86204 1366 86216
rect 1397 86207 1455 86213
rect 1397 86204 1409 86207
rect 1360 86176 1409 86204
rect 1360 86164 1366 86176
rect 1397 86173 1409 86176
rect 1443 86204 1455 86207
rect 1673 86207 1731 86213
rect 1673 86204 1685 86207
rect 1443 86176 1685 86204
rect 1443 86173 1455 86176
rect 1397 86167 1455 86173
rect 1673 86173 1685 86176
rect 1719 86173 1731 86207
rect 1673 86167 1731 86173
rect 1854 86096 1860 86148
rect 1912 86136 1918 86148
rect 8570 86136 8576 86148
rect 1912 86108 8576 86136
rect 1912 86096 1918 86108
rect 8570 86096 8576 86108
rect 8628 86096 8634 86148
rect 1581 86071 1639 86077
rect 1581 86037 1593 86071
rect 1627 86068 1639 86071
rect 5994 86068 6000 86080
rect 1627 86040 6000 86068
rect 1627 86037 1639 86040
rect 1581 86031 1639 86037
rect 5994 86028 6000 86040
rect 6052 86028 6058 86080
rect 1104 85978 7912 86000
rect 1104 85926 4874 85978
rect 4926 85926 4938 85978
rect 4990 85926 5002 85978
rect 5054 85926 5066 85978
rect 5118 85926 5130 85978
rect 5182 85926 7912 85978
rect 1104 85904 7912 85926
rect 104052 85978 108836 86000
rect 104052 85926 106658 85978
rect 106710 85926 106722 85978
rect 106774 85926 106786 85978
rect 106838 85926 106850 85978
rect 106902 85926 106914 85978
rect 106966 85926 108836 85978
rect 104052 85904 108836 85926
rect 1104 85434 7912 85456
rect 1104 85382 4214 85434
rect 4266 85382 4278 85434
rect 4330 85382 4342 85434
rect 4394 85382 4406 85434
rect 4458 85382 4470 85434
rect 4522 85382 7912 85434
rect 1104 85360 7912 85382
rect 104052 85434 108836 85456
rect 104052 85382 105922 85434
rect 105974 85382 105986 85434
rect 106038 85382 106050 85434
rect 106102 85382 106114 85434
rect 106166 85382 106178 85434
rect 106230 85382 108836 85434
rect 104052 85360 108836 85382
rect 1210 85008 1216 85060
rect 1268 85048 1274 85060
rect 1489 85051 1547 85057
rect 1489 85048 1501 85051
rect 1268 85020 1501 85048
rect 1268 85008 1274 85020
rect 1489 85017 1501 85020
rect 1535 85048 1547 85051
rect 1949 85051 2007 85057
rect 1949 85048 1961 85051
rect 1535 85020 1961 85048
rect 1535 85017 1547 85020
rect 1489 85011 1547 85017
rect 1949 85017 1961 85020
rect 1995 85017 2007 85051
rect 1949 85011 2007 85017
rect 1581 84983 1639 84989
rect 1581 84949 1593 84983
rect 1627 84980 1639 84983
rect 1762 84980 1768 84992
rect 1627 84952 1768 84980
rect 1627 84949 1639 84952
rect 1581 84943 1639 84949
rect 1762 84940 1768 84952
rect 1820 84940 1826 84992
rect 1104 84890 7912 84912
rect 1104 84838 4874 84890
rect 4926 84838 4938 84890
rect 4990 84838 5002 84890
rect 5054 84838 5066 84890
rect 5118 84838 5130 84890
rect 5182 84838 7912 84890
rect 1104 84816 7912 84838
rect 104052 84890 108836 84912
rect 104052 84838 106658 84890
rect 106710 84838 106722 84890
rect 106774 84838 106786 84890
rect 106838 84838 106850 84890
rect 106902 84838 106914 84890
rect 106966 84838 108836 84890
rect 104052 84816 108836 84838
rect 1302 84600 1308 84652
rect 1360 84640 1366 84652
rect 1489 84643 1547 84649
rect 1489 84640 1501 84643
rect 1360 84612 1501 84640
rect 1360 84600 1366 84612
rect 1489 84609 1501 84612
rect 1535 84640 1547 84643
rect 1949 84643 2007 84649
rect 1949 84640 1961 84643
rect 1535 84612 1961 84640
rect 1535 84609 1547 84612
rect 1489 84603 1547 84609
rect 1949 84609 1961 84612
rect 1995 84609 2007 84643
rect 1949 84603 2007 84609
rect 1673 84507 1731 84513
rect 1673 84473 1685 84507
rect 1719 84504 1731 84507
rect 1765 84507 1823 84513
rect 1765 84504 1777 84507
rect 1719 84476 1777 84504
rect 1719 84473 1731 84476
rect 1673 84467 1731 84473
rect 1765 84473 1777 84476
rect 1811 84504 1823 84507
rect 1854 84504 1860 84516
rect 1811 84476 1860 84504
rect 1811 84473 1823 84476
rect 1765 84467 1823 84473
rect 1854 84464 1860 84476
rect 1912 84464 1918 84516
rect 1104 84346 7912 84368
rect 1104 84294 4214 84346
rect 4266 84294 4278 84346
rect 4330 84294 4342 84346
rect 4394 84294 4406 84346
rect 4458 84294 4470 84346
rect 4522 84294 7912 84346
rect 1104 84272 7912 84294
rect 104052 84346 108836 84368
rect 104052 84294 105922 84346
rect 105974 84294 105986 84346
rect 106038 84294 106050 84346
rect 106102 84294 106114 84346
rect 106166 84294 106178 84346
rect 106230 84294 108836 84346
rect 104052 84272 108836 84294
rect 1946 84124 1952 84176
rect 2004 84164 2010 84176
rect 9398 84164 9404 84176
rect 2004 84136 9404 84164
rect 2004 84124 2010 84136
rect 9398 84124 9404 84136
rect 9456 84124 9462 84176
rect 1302 83920 1308 83972
rect 1360 83960 1366 83972
rect 1489 83963 1547 83969
rect 1489 83960 1501 83963
rect 1360 83932 1501 83960
rect 1360 83920 1366 83932
rect 1489 83929 1501 83932
rect 1535 83929 1547 83963
rect 1489 83923 1547 83929
rect 1673 83963 1731 83969
rect 1673 83929 1685 83963
rect 1719 83960 1731 83963
rect 1857 83963 1915 83969
rect 1857 83960 1869 83963
rect 1719 83932 1869 83960
rect 1719 83929 1731 83932
rect 1673 83923 1731 83929
rect 1857 83929 1869 83932
rect 1903 83960 1915 83963
rect 8478 83960 8484 83972
rect 1903 83932 8484 83960
rect 1903 83929 1915 83932
rect 1857 83923 1915 83929
rect 1504 83892 1532 83923
rect 8478 83920 8484 83932
rect 8536 83920 8542 83972
rect 1949 83895 2007 83901
rect 1949 83892 1961 83895
rect 1504 83864 1961 83892
rect 1949 83861 1961 83864
rect 1995 83861 2007 83895
rect 1949 83855 2007 83861
rect 1104 83802 7912 83824
rect 1104 83750 4874 83802
rect 4926 83750 4938 83802
rect 4990 83750 5002 83802
rect 5054 83750 5066 83802
rect 5118 83750 5130 83802
rect 5182 83750 7912 83802
rect 1104 83728 7912 83750
rect 104052 83802 108836 83824
rect 104052 83750 106658 83802
rect 106710 83750 106722 83802
rect 106774 83750 106786 83802
rect 106838 83750 106850 83802
rect 106902 83750 106914 83802
rect 106966 83750 108836 83802
rect 104052 83728 108836 83750
rect 1302 83512 1308 83564
rect 1360 83552 1366 83564
rect 1489 83555 1547 83561
rect 1489 83552 1501 83555
rect 1360 83524 1501 83552
rect 1360 83512 1366 83524
rect 1489 83521 1501 83524
rect 1535 83552 1547 83555
rect 1949 83555 2007 83561
rect 1949 83552 1961 83555
rect 1535 83524 1961 83552
rect 1535 83521 1547 83524
rect 1489 83515 1547 83521
rect 1949 83521 1961 83524
rect 1995 83521 2007 83555
rect 1949 83515 2007 83521
rect 1581 83351 1639 83357
rect 1581 83317 1593 83351
rect 1627 83348 1639 83351
rect 1857 83351 1915 83357
rect 1857 83348 1869 83351
rect 1627 83320 1869 83348
rect 1627 83317 1639 83320
rect 1581 83311 1639 83317
rect 1857 83317 1869 83320
rect 1903 83348 1915 83351
rect 2498 83348 2504 83360
rect 1903 83320 2504 83348
rect 1903 83317 1915 83320
rect 1857 83311 1915 83317
rect 2498 83308 2504 83320
rect 2556 83308 2562 83360
rect 1104 83258 7912 83280
rect 1104 83206 4214 83258
rect 4266 83206 4278 83258
rect 4330 83206 4342 83258
rect 4394 83206 4406 83258
rect 4458 83206 4470 83258
rect 4522 83206 7912 83258
rect 1104 83184 7912 83206
rect 104052 83258 108836 83280
rect 104052 83206 105922 83258
rect 105974 83206 105986 83258
rect 106038 83206 106050 83258
rect 106102 83206 106114 83258
rect 106166 83206 106178 83258
rect 106230 83206 108836 83258
rect 104052 83184 108836 83206
rect 1854 82764 1860 82816
rect 1912 82804 1918 82816
rect 9214 82804 9220 82816
rect 1912 82776 9220 82804
rect 1912 82764 1918 82776
rect 9214 82764 9220 82776
rect 9272 82764 9278 82816
rect 1104 82714 7912 82736
rect 1104 82662 4874 82714
rect 4926 82662 4938 82714
rect 4990 82662 5002 82714
rect 5054 82662 5066 82714
rect 5118 82662 5130 82714
rect 5182 82662 7912 82714
rect 1104 82640 7912 82662
rect 104052 82714 108836 82736
rect 104052 82662 106658 82714
rect 106710 82662 106722 82714
rect 106774 82662 106786 82714
rect 106838 82662 106850 82714
rect 106902 82662 106914 82714
rect 106966 82662 108836 82714
rect 104052 82640 108836 82662
rect 1210 82424 1216 82476
rect 1268 82464 1274 82476
rect 1489 82467 1547 82473
rect 1489 82464 1501 82467
rect 1268 82436 1501 82464
rect 1268 82424 1274 82436
rect 1489 82433 1501 82436
rect 1535 82464 1547 82467
rect 1949 82467 2007 82473
rect 1949 82464 1961 82467
rect 1535 82436 1961 82464
rect 1535 82433 1547 82436
rect 1489 82427 1547 82433
rect 1949 82433 1961 82436
rect 1995 82433 2007 82467
rect 1949 82427 2007 82433
rect 1581 82263 1639 82269
rect 1581 82229 1593 82263
rect 1627 82260 1639 82263
rect 1857 82263 1915 82269
rect 1857 82260 1869 82263
rect 1627 82232 1869 82260
rect 1627 82229 1639 82232
rect 1581 82223 1639 82229
rect 1857 82229 1869 82232
rect 1903 82260 1915 82263
rect 2406 82260 2412 82272
rect 1903 82232 2412 82260
rect 1903 82229 1915 82232
rect 1857 82223 1915 82229
rect 2406 82220 2412 82232
rect 2464 82220 2470 82272
rect 1104 82170 7912 82192
rect 1104 82118 4214 82170
rect 4266 82118 4278 82170
rect 4330 82118 4342 82170
rect 4394 82118 4406 82170
rect 4458 82118 4470 82170
rect 4522 82118 7912 82170
rect 1104 82096 7912 82118
rect 104052 82170 108836 82192
rect 104052 82118 105922 82170
rect 105974 82118 105986 82170
rect 106038 82118 106050 82170
rect 106102 82118 106114 82170
rect 106166 82118 106178 82170
rect 106230 82118 108836 82170
rect 104052 82096 108836 82118
rect 1210 81744 1216 81796
rect 1268 81784 1274 81796
rect 1489 81787 1547 81793
rect 1489 81784 1501 81787
rect 1268 81756 1501 81784
rect 1268 81744 1274 81756
rect 1489 81753 1501 81756
rect 1535 81784 1547 81787
rect 1949 81787 2007 81793
rect 1949 81784 1961 81787
rect 1535 81756 1961 81784
rect 1535 81753 1547 81756
rect 1489 81747 1547 81753
rect 1949 81753 1961 81756
rect 1995 81753 2007 81787
rect 1949 81747 2007 81753
rect 1581 81719 1639 81725
rect 1581 81685 1593 81719
rect 1627 81716 1639 81719
rect 1854 81716 1860 81728
rect 1627 81688 1860 81716
rect 1627 81685 1639 81688
rect 1581 81679 1639 81685
rect 1854 81676 1860 81688
rect 1912 81676 1918 81728
rect 1104 81626 7912 81648
rect 1104 81574 4874 81626
rect 4926 81574 4938 81626
rect 4990 81574 5002 81626
rect 5054 81574 5066 81626
rect 5118 81574 5130 81626
rect 5182 81574 7912 81626
rect 1104 81552 7912 81574
rect 104052 81626 108836 81648
rect 104052 81574 106658 81626
rect 106710 81574 106722 81626
rect 106774 81574 106786 81626
rect 106838 81574 106850 81626
rect 106902 81574 106914 81626
rect 106966 81574 108836 81626
rect 104052 81552 108836 81574
rect 1302 81336 1308 81388
rect 1360 81376 1366 81388
rect 1489 81379 1547 81385
rect 1489 81376 1501 81379
rect 1360 81348 1501 81376
rect 1360 81336 1366 81348
rect 1489 81345 1501 81348
rect 1535 81376 1547 81379
rect 1949 81379 2007 81385
rect 1949 81376 1961 81379
rect 1535 81348 1961 81376
rect 1535 81345 1547 81348
rect 1489 81339 1547 81345
rect 1949 81345 1961 81348
rect 1995 81345 2007 81379
rect 1949 81339 2007 81345
rect 1854 81200 1860 81252
rect 1912 81240 1918 81252
rect 9766 81240 9772 81252
rect 1912 81212 9772 81240
rect 1912 81200 1918 81212
rect 9766 81200 9772 81212
rect 9824 81200 9830 81252
rect 1581 81175 1639 81181
rect 1581 81141 1593 81175
rect 1627 81172 1639 81175
rect 1765 81175 1823 81181
rect 1765 81172 1777 81175
rect 1627 81144 1777 81172
rect 1627 81141 1639 81144
rect 1581 81135 1639 81141
rect 1765 81141 1777 81144
rect 1811 81172 1823 81175
rect 5626 81172 5632 81184
rect 1811 81144 5632 81172
rect 1811 81141 1823 81144
rect 1765 81135 1823 81141
rect 5626 81132 5632 81144
rect 5684 81132 5690 81184
rect 1104 81082 7912 81104
rect 1104 81030 4214 81082
rect 4266 81030 4278 81082
rect 4330 81030 4342 81082
rect 4394 81030 4406 81082
rect 4458 81030 4470 81082
rect 4522 81030 7912 81082
rect 1104 81008 7912 81030
rect 104052 81082 108836 81104
rect 104052 81030 105922 81082
rect 105974 81030 105986 81082
rect 106038 81030 106050 81082
rect 106102 81030 106114 81082
rect 106166 81030 106178 81082
rect 106230 81030 108836 81082
rect 104052 81008 108836 81030
rect 2406 80792 2412 80844
rect 2464 80832 2470 80844
rect 9858 80832 9864 80844
rect 2464 80804 9864 80832
rect 2464 80792 2470 80804
rect 9858 80792 9864 80804
rect 9916 80792 9922 80844
rect 1302 80724 1308 80776
rect 1360 80764 1366 80776
rect 1397 80767 1455 80773
rect 1397 80764 1409 80767
rect 1360 80736 1409 80764
rect 1360 80724 1366 80736
rect 1397 80733 1409 80736
rect 1443 80733 1455 80767
rect 1397 80727 1455 80733
rect 1673 80767 1731 80773
rect 1673 80733 1685 80767
rect 1719 80764 1731 80767
rect 1719 80736 2452 80764
rect 1719 80733 1731 80736
rect 1673 80727 1731 80733
rect 2424 80637 2452 80736
rect 2498 80656 2504 80708
rect 2556 80696 2562 80708
rect 9950 80696 9956 80708
rect 2556 80668 9956 80696
rect 2556 80656 2562 80668
rect 9950 80656 9956 80668
rect 10008 80656 10014 80708
rect 2409 80631 2467 80637
rect 2409 80597 2421 80631
rect 2455 80628 2467 80631
rect 5534 80628 5540 80640
rect 2455 80600 5540 80628
rect 2455 80597 2467 80600
rect 2409 80591 2467 80597
rect 5534 80588 5540 80600
rect 5592 80588 5598 80640
rect 1104 80538 7912 80560
rect 1104 80486 4874 80538
rect 4926 80486 4938 80538
rect 4990 80486 5002 80538
rect 5054 80486 5066 80538
rect 5118 80486 5130 80538
rect 5182 80486 7912 80538
rect 1104 80464 7912 80486
rect 104052 80538 108836 80560
rect 104052 80486 106658 80538
rect 106710 80486 106722 80538
rect 106774 80486 106786 80538
rect 106838 80486 106850 80538
rect 106902 80486 106914 80538
rect 106966 80486 108836 80538
rect 104052 80464 108836 80486
rect 1302 80316 1308 80368
rect 1360 80356 1366 80368
rect 1397 80359 1455 80365
rect 1397 80356 1409 80359
rect 1360 80328 1409 80356
rect 1360 80316 1366 80328
rect 1397 80325 1409 80328
rect 1443 80325 1455 80359
rect 1397 80319 1455 80325
rect 1104 79994 7912 80016
rect 1104 79942 4214 79994
rect 4266 79942 4278 79994
rect 4330 79942 4342 79994
rect 4394 79942 4406 79994
rect 4458 79942 4470 79994
rect 4522 79942 7912 79994
rect 9950 79976 9956 80028
rect 10008 80016 10014 80028
rect 40954 80016 40960 80028
rect 10008 79988 40960 80016
rect 10008 79976 10014 79988
rect 40954 79976 40960 79988
rect 41012 79976 41018 80028
rect 104052 79994 108836 80016
rect 1104 79920 7912 79942
rect 9858 79908 9864 79960
rect 9916 79948 9922 79960
rect 39758 79948 39764 79960
rect 9916 79920 39764 79948
rect 9916 79908 9922 79920
rect 39758 79908 39764 79920
rect 39816 79908 39822 79960
rect 104052 79942 105922 79994
rect 105974 79942 105986 79994
rect 106038 79942 106050 79994
rect 106102 79942 106114 79994
rect 106166 79942 106178 79994
rect 106230 79942 108836 79994
rect 104052 79920 108836 79942
rect 9766 79840 9772 79892
rect 9824 79880 9830 79892
rect 38654 79880 38660 79892
rect 9824 79852 38660 79880
rect 9824 79840 9830 79852
rect 38654 79840 38660 79852
rect 38712 79840 38718 79892
rect 8938 79772 8944 79824
rect 8996 79812 9002 79824
rect 36262 79812 36268 79824
rect 8996 79784 36268 79812
rect 8996 79772 9002 79784
rect 36262 79772 36268 79784
rect 36320 79772 36326 79824
rect 8570 79704 8576 79756
rect 8628 79744 8634 79756
rect 34698 79744 34704 79756
rect 8628 79716 34704 79744
rect 8628 79704 8634 79716
rect 34698 79704 34704 79716
rect 34756 79704 34762 79756
rect 9214 79636 9220 79688
rect 9272 79676 9278 79688
rect 32306 79676 32312 79688
rect 9272 79648 32312 79676
rect 9272 79636 9278 79648
rect 32306 79636 32312 79648
rect 32364 79636 32370 79688
rect 1210 79568 1216 79620
rect 1268 79608 1274 79620
rect 1489 79611 1547 79617
rect 1489 79608 1501 79611
rect 1268 79580 1501 79608
rect 1268 79568 1274 79580
rect 1489 79577 1501 79580
rect 1535 79577 1547 79611
rect 1489 79571 1547 79577
rect 1673 79611 1731 79617
rect 1673 79577 1685 79611
rect 1719 79608 1731 79611
rect 1857 79611 1915 79617
rect 1857 79608 1869 79611
rect 1719 79580 1869 79608
rect 1719 79577 1731 79580
rect 1673 79571 1731 79577
rect 1857 79577 1869 79580
rect 1903 79608 1915 79611
rect 1903 79580 6914 79608
rect 1903 79577 1915 79580
rect 1857 79571 1915 79577
rect 1504 79540 1532 79571
rect 1949 79543 2007 79549
rect 1949 79540 1961 79543
rect 1504 79512 1961 79540
rect 1949 79509 1961 79512
rect 1995 79509 2007 79543
rect 6886 79540 6914 79580
rect 36998 79540 37004 79552
rect 6886 79512 37004 79540
rect 1949 79503 2007 79509
rect 36998 79500 37004 79512
rect 37056 79500 37062 79552
rect 1104 79450 7912 79472
rect 1104 79398 4874 79450
rect 4926 79398 4938 79450
rect 4990 79398 5002 79450
rect 5054 79398 5066 79450
rect 5118 79398 5130 79450
rect 5182 79398 7912 79450
rect 1104 79376 7912 79398
rect 104052 79450 108836 79472
rect 104052 79398 106658 79450
rect 106710 79398 106722 79450
rect 106774 79398 106786 79450
rect 106838 79398 106850 79450
rect 106902 79398 106914 79450
rect 106966 79398 108836 79450
rect 104052 79376 108836 79398
rect 61102 79296 61108 79348
rect 61160 79336 61166 79348
rect 101950 79336 101956 79348
rect 61160 79308 101956 79336
rect 61160 79296 61166 79308
rect 101950 79296 101956 79308
rect 102008 79296 102014 79348
rect 1302 79160 1308 79212
rect 1360 79200 1366 79212
rect 1489 79203 1547 79209
rect 1489 79200 1501 79203
rect 1360 79172 1501 79200
rect 1360 79160 1366 79172
rect 1489 79169 1501 79172
rect 1535 79200 1547 79203
rect 1949 79203 2007 79209
rect 1949 79200 1961 79203
rect 1535 79172 1961 79200
rect 1535 79169 1547 79172
rect 1489 79163 1547 79169
rect 1949 79169 1961 79172
rect 1995 79169 2007 79203
rect 108301 79203 108359 79209
rect 108301 79200 108313 79203
rect 1949 79163 2007 79169
rect 108132 79172 108313 79200
rect 1673 79067 1731 79073
rect 1673 79033 1685 79067
rect 1719 79064 1731 79067
rect 1857 79067 1915 79073
rect 1857 79064 1869 79067
rect 1719 79036 1869 79064
rect 1719 79033 1731 79036
rect 1673 79027 1731 79033
rect 1857 79033 1869 79036
rect 1903 79064 1915 79067
rect 1903 79036 6914 79064
rect 1903 79033 1915 79036
rect 1857 79027 1915 79033
rect 6886 78996 6914 79036
rect 42150 78996 42156 79008
rect 6886 78968 42156 78996
rect 42150 78956 42156 78968
rect 42208 78956 42214 79008
rect 88886 78956 88892 79008
rect 88944 78996 88950 79008
rect 108132 79005 108160 79172
rect 108301 79169 108313 79172
rect 108347 79169 108359 79203
rect 108301 79163 108359 79169
rect 108117 78999 108175 79005
rect 108117 78996 108129 78999
rect 88944 78968 108129 78996
rect 88944 78956 88950 78968
rect 108117 78965 108129 78968
rect 108163 78965 108175 78999
rect 108117 78959 108175 78965
rect 108482 78956 108488 79008
rect 108540 78956 108546 79008
rect 1104 78906 7912 78928
rect 1104 78854 4214 78906
rect 4266 78854 4278 78906
rect 4330 78854 4342 78906
rect 4394 78854 4406 78906
rect 4458 78854 4470 78906
rect 4522 78854 7912 78906
rect 1104 78832 7912 78854
rect 104052 78906 108836 78928
rect 104052 78854 105922 78906
rect 105974 78854 105986 78906
rect 106038 78854 106050 78906
rect 106102 78854 106114 78906
rect 106166 78854 106178 78906
rect 106230 78854 108836 78906
rect 104052 78832 108836 78854
rect 96522 78548 96528 78600
rect 96580 78588 96586 78600
rect 102134 78588 102140 78600
rect 96580 78560 102140 78588
rect 96580 78548 96586 78560
rect 102134 78548 102140 78560
rect 102192 78548 102198 78600
rect 108301 78591 108359 78597
rect 108301 78588 108313 78591
rect 108132 78560 108313 78588
rect 1302 78480 1308 78532
rect 1360 78520 1366 78532
rect 1489 78523 1547 78529
rect 1489 78520 1501 78523
rect 1360 78492 1501 78520
rect 1360 78480 1366 78492
rect 1489 78489 1501 78492
rect 1535 78489 1547 78523
rect 1489 78483 1547 78489
rect 1673 78523 1731 78529
rect 1673 78489 1685 78523
rect 1719 78520 1731 78523
rect 1857 78523 1915 78529
rect 1857 78520 1869 78523
rect 1719 78492 1869 78520
rect 1719 78489 1731 78492
rect 1673 78483 1731 78489
rect 1857 78489 1869 78492
rect 1903 78520 1915 78523
rect 1903 78492 6914 78520
rect 1903 78489 1915 78492
rect 1857 78483 1915 78489
rect 1504 78452 1532 78483
rect 1949 78455 2007 78461
rect 1949 78452 1961 78455
rect 1504 78424 1961 78452
rect 1949 78421 1961 78424
rect 1995 78421 2007 78455
rect 6886 78452 6914 78492
rect 79226 78480 79232 78532
rect 79284 78520 79290 78532
rect 91646 78520 91652 78532
rect 79284 78492 91652 78520
rect 79284 78480 79290 78492
rect 91646 78480 91652 78492
rect 91704 78480 91710 78532
rect 108132 78464 108160 78560
rect 108301 78557 108313 78560
rect 108347 78557 108359 78591
rect 108301 78551 108359 78557
rect 29546 78452 29552 78464
rect 6886 78424 29552 78452
rect 1949 78415 2007 78421
rect 29546 78412 29552 78424
rect 29604 78412 29610 78464
rect 76650 78412 76656 78464
rect 76708 78452 76714 78464
rect 89806 78452 89812 78464
rect 76708 78424 89812 78452
rect 76708 78412 76714 78424
rect 89806 78412 89812 78424
rect 89864 78412 89870 78464
rect 108114 78412 108120 78464
rect 108172 78412 108178 78464
rect 108482 78412 108488 78464
rect 108540 78412 108546 78464
rect 1104 78362 7912 78384
rect 1104 78310 4874 78362
rect 4926 78310 4938 78362
rect 4990 78310 5002 78362
rect 5054 78310 5066 78362
rect 5118 78310 5130 78362
rect 5182 78310 7912 78362
rect 71958 78344 71964 78396
rect 72016 78384 72022 78396
rect 85666 78384 85672 78396
rect 72016 78356 85672 78384
rect 72016 78344 72022 78356
rect 85666 78344 85672 78356
rect 85724 78344 85730 78396
rect 104052 78362 108836 78384
rect 1104 78288 7912 78310
rect 22738 78276 22744 78328
rect 22796 78316 22802 78328
rect 22796 78288 25268 78316
rect 22796 78276 22802 78288
rect 22094 78208 22100 78260
rect 22152 78248 22158 78260
rect 22152 78220 25176 78248
rect 22152 78208 22158 78220
rect 2314 78140 2320 78192
rect 2372 78180 2378 78192
rect 2372 78152 6914 78180
rect 2372 78140 2378 78152
rect 1302 78072 1308 78124
rect 1360 78112 1366 78124
rect 1489 78115 1547 78121
rect 1489 78112 1501 78115
rect 1360 78084 1501 78112
rect 1360 78072 1366 78084
rect 1489 78081 1501 78084
rect 1535 78112 1547 78115
rect 1949 78115 2007 78121
rect 1949 78112 1961 78115
rect 1535 78084 1961 78112
rect 1535 78081 1547 78084
rect 1489 78075 1547 78081
rect 1949 78081 1961 78084
rect 1995 78081 2007 78115
rect 6886 78112 6914 78152
rect 25038 78112 25044 78124
rect 6886 78084 25044 78112
rect 1949 78075 2007 78081
rect 25038 78072 25044 78084
rect 25096 78072 25102 78124
rect 25148 78112 25176 78220
rect 25240 78180 25268 78288
rect 73522 78276 73528 78328
rect 73580 78316 73586 78328
rect 80054 78316 80060 78328
rect 73580 78288 80060 78316
rect 73580 78276 73586 78288
rect 80054 78276 80060 78288
rect 80112 78276 80118 78328
rect 104052 78310 106658 78362
rect 106710 78310 106722 78362
rect 106774 78310 106786 78362
rect 106838 78310 106850 78362
rect 106902 78310 106914 78362
rect 106966 78310 108836 78362
rect 104052 78288 108836 78310
rect 26050 78208 26056 78260
rect 26108 78248 26114 78260
rect 30282 78248 30288 78260
rect 26108 78220 30288 78248
rect 26108 78208 26114 78220
rect 30282 78208 30288 78220
rect 30340 78208 30346 78260
rect 69750 78208 69756 78260
rect 69808 78248 69814 78260
rect 102410 78248 102416 78260
rect 69808 78220 102416 78248
rect 69808 78208 69814 78220
rect 102410 78208 102416 78220
rect 102468 78208 102474 78260
rect 34790 78180 34796 78192
rect 25240 78152 34796 78180
rect 34790 78140 34796 78152
rect 34848 78140 34854 78192
rect 63954 78140 63960 78192
rect 64012 78180 64018 78192
rect 81342 78180 81348 78192
rect 64012 78152 81348 78180
rect 64012 78140 64018 78152
rect 81342 78140 81348 78152
rect 81400 78140 81406 78192
rect 25148 78084 30696 78112
rect 20806 78004 20812 78056
rect 20864 78044 20870 78056
rect 27246 78044 27252 78056
rect 20864 78016 27252 78044
rect 20864 78004 20870 78016
rect 27246 78004 27252 78016
rect 27304 78004 27310 78056
rect 1673 77979 1731 77985
rect 1673 77945 1685 77979
rect 1719 77976 1731 77979
rect 1857 77979 1915 77985
rect 1857 77976 1869 77979
rect 1719 77948 1869 77976
rect 1719 77945 1731 77948
rect 1673 77939 1731 77945
rect 1857 77945 1869 77948
rect 1903 77976 1915 77979
rect 1903 77948 6914 77976
rect 1903 77945 1915 77948
rect 1857 77939 1915 77945
rect 6886 77908 6914 77948
rect 21266 77936 21272 77988
rect 21324 77976 21330 77988
rect 30558 77976 30564 77988
rect 21324 77948 30564 77976
rect 21324 77936 21330 77948
rect 30558 77936 30564 77948
rect 30616 77936 30622 77988
rect 30668 77976 30696 78084
rect 31478 78072 31484 78124
rect 31536 78112 31542 78124
rect 33962 78112 33968 78124
rect 31536 78084 33968 78112
rect 31536 78072 31542 78084
rect 33962 78072 33968 78084
rect 34020 78072 34026 78124
rect 63586 78072 63592 78124
rect 63644 78112 63650 78124
rect 71130 78112 71136 78124
rect 63644 78084 71136 78112
rect 63644 78072 63650 78084
rect 71130 78072 71136 78084
rect 71188 78072 71194 78124
rect 74442 78072 74448 78124
rect 74500 78112 74506 78124
rect 88978 78112 88984 78124
rect 74500 78084 88984 78112
rect 74500 78072 74506 78084
rect 88978 78072 88984 78084
rect 89036 78072 89042 78124
rect 102594 78112 102600 78124
rect 89088 78084 102600 78112
rect 30742 78004 30748 78056
rect 30800 78044 30806 78056
rect 39850 78044 39856 78056
rect 30800 78016 39856 78044
rect 30800 78004 30806 78016
rect 39850 78004 39856 78016
rect 39908 78004 39914 78056
rect 58618 78004 58624 78056
rect 58676 78044 58682 78056
rect 58676 78016 64368 78044
rect 58676 78004 58682 78016
rect 43254 77976 43260 77988
rect 30668 77948 43260 77976
rect 43254 77936 43260 77948
rect 43312 77976 43318 77988
rect 43806 77976 43812 77988
rect 43312 77948 43812 77976
rect 43312 77936 43318 77948
rect 43806 77936 43812 77948
rect 43864 77936 43870 77988
rect 53558 77936 53564 77988
rect 53616 77976 53622 77988
rect 62482 77976 62488 77988
rect 53616 77948 62488 77976
rect 53616 77936 53622 77948
rect 62482 77936 62488 77948
rect 62540 77936 62546 77988
rect 31478 77908 31484 77920
rect 6886 77880 31484 77908
rect 31478 77868 31484 77880
rect 31536 77868 31542 77920
rect 31662 77868 31668 77920
rect 31720 77908 31726 77920
rect 36078 77908 36084 77920
rect 31720 77880 36084 77908
rect 31720 77868 31726 77880
rect 36078 77868 36084 77880
rect 36136 77868 36142 77920
rect 56134 77868 56140 77920
rect 56192 77908 56198 77920
rect 64138 77908 64144 77920
rect 56192 77880 64144 77908
rect 56192 77868 56198 77880
rect 64138 77868 64144 77880
rect 64196 77868 64202 77920
rect 64340 77908 64368 78016
rect 69106 78004 69112 78056
rect 69164 78044 69170 78056
rect 85942 78044 85948 78056
rect 69164 78016 85948 78044
rect 69164 78004 69170 78016
rect 85942 78004 85948 78016
rect 86000 78004 86006 78056
rect 87322 78004 87328 78056
rect 87380 78044 87386 78056
rect 89088 78044 89116 78084
rect 102594 78072 102600 78084
rect 102652 78072 102658 78124
rect 108301 78115 108359 78121
rect 108301 78112 108313 78115
rect 108132 78084 108313 78112
rect 87380 78016 89116 78044
rect 87380 78004 87386 78016
rect 93118 78004 93124 78056
rect 93176 78044 93182 78056
rect 107654 78044 107660 78056
rect 93176 78016 107660 78044
rect 93176 78004 93182 78016
rect 107654 78004 107660 78016
rect 107712 78004 107718 78056
rect 66070 77936 66076 77988
rect 66128 77976 66134 77988
rect 73430 77976 73436 77988
rect 66128 77948 73436 77976
rect 66128 77936 66134 77948
rect 73430 77936 73436 77948
rect 73488 77936 73494 77988
rect 80882 77936 80888 77988
rect 80940 77976 80946 77988
rect 94222 77976 94228 77988
rect 80940 77948 94228 77976
rect 80940 77936 80946 77948
rect 94222 77936 94228 77948
rect 94280 77936 94286 77988
rect 67634 77908 67640 77920
rect 64340 77880 67640 77908
rect 67634 77868 67640 77880
rect 67692 77868 67698 77920
rect 70394 77868 70400 77920
rect 70452 77908 70458 77920
rect 87046 77908 87052 77920
rect 70452 77880 87052 77908
rect 70452 77868 70458 77880
rect 87046 77868 87052 77880
rect 87104 77868 87110 77920
rect 90726 77868 90732 77920
rect 90784 77908 90790 77920
rect 99650 77908 99656 77920
rect 90784 77880 99656 77908
rect 90784 77868 90790 77880
rect 99650 77868 99656 77880
rect 99708 77868 99714 77920
rect 105814 77868 105820 77920
rect 105872 77908 105878 77920
rect 108132 77917 108160 78084
rect 108301 78081 108313 78084
rect 108347 78081 108359 78115
rect 108301 78075 108359 78081
rect 108117 77911 108175 77917
rect 108117 77908 108129 77911
rect 105872 77880 108129 77908
rect 105872 77868 105878 77880
rect 108117 77877 108129 77880
rect 108163 77877 108175 77911
rect 108117 77871 108175 77877
rect 108482 77868 108488 77920
rect 108540 77868 108546 77920
rect 1104 77818 108836 77840
rect 1104 77766 4214 77818
rect 4266 77766 4278 77818
rect 4330 77766 4342 77818
rect 4394 77766 4406 77818
rect 4458 77766 4470 77818
rect 4522 77766 34934 77818
rect 34986 77766 34998 77818
rect 35050 77766 35062 77818
rect 35114 77766 35126 77818
rect 35178 77766 35190 77818
rect 35242 77766 65654 77818
rect 65706 77766 65718 77818
rect 65770 77766 65782 77818
rect 65834 77766 65846 77818
rect 65898 77766 65910 77818
rect 65962 77766 96374 77818
rect 96426 77766 96438 77818
rect 96490 77766 96502 77818
rect 96554 77766 96566 77818
rect 96618 77766 96630 77818
rect 96682 77766 105922 77818
rect 105974 77766 105986 77818
rect 106038 77766 106050 77818
rect 106102 77766 106114 77818
rect 106166 77766 106178 77818
rect 106230 77766 108836 77818
rect 1104 77744 108836 77766
rect 21821 77707 21879 77713
rect 21821 77704 21833 77707
rect 19812 77676 21833 77704
rect 17862 77596 17868 77648
rect 17920 77636 17926 77648
rect 19812 77645 19840 77676
rect 21821 77673 21833 77676
rect 21867 77673 21879 77707
rect 27522 77704 27528 77716
rect 21821 77667 21879 77673
rect 23860 77676 27528 77704
rect 19797 77639 19855 77645
rect 19797 77636 19809 77639
rect 17920 77608 19809 77636
rect 17920 77596 17926 77608
rect 19797 77605 19809 77608
rect 19843 77605 19855 77639
rect 19797 77599 19855 77605
rect 21542 77568 21548 77580
rect 19628 77540 21548 77568
rect 6822 77324 6828 77376
rect 6880 77364 6886 77376
rect 16022 77364 16028 77376
rect 6880 77336 16028 77364
rect 6880 77324 6886 77336
rect 16022 77324 16028 77336
rect 16080 77364 16086 77376
rect 19628 77373 19656 77540
rect 21542 77528 21548 77540
rect 21600 77568 21606 77580
rect 22281 77571 22339 77577
rect 22281 77568 22293 77571
rect 21600 77540 22293 77568
rect 21600 77528 21606 77540
rect 22281 77537 22293 77540
rect 22327 77568 22339 77571
rect 22465 77571 22523 77577
rect 22465 77568 22477 77571
rect 22327 77540 22477 77568
rect 22327 77537 22339 77540
rect 22281 77531 22339 77537
rect 22465 77537 22477 77540
rect 22511 77537 22523 77571
rect 22465 77531 22523 77537
rect 22738 77528 22744 77580
rect 22796 77528 22802 77580
rect 23860 77486 23888 77676
rect 27522 77664 27528 77676
rect 27580 77664 27586 77716
rect 27614 77664 27620 77716
rect 27672 77664 27678 77716
rect 28166 77664 28172 77716
rect 28224 77664 28230 77716
rect 29546 77664 29552 77716
rect 29604 77664 29610 77716
rect 30466 77664 30472 77716
rect 30524 77664 30530 77716
rect 30558 77664 30564 77716
rect 30616 77704 30622 77716
rect 30745 77707 30803 77713
rect 30745 77704 30757 77707
rect 30616 77676 30757 77704
rect 30616 77664 30622 77676
rect 30745 77673 30757 77676
rect 30791 77673 30803 77707
rect 30745 77667 30803 77673
rect 31662 77664 31668 77716
rect 31720 77664 31726 77716
rect 32306 77664 32312 77716
rect 32364 77704 32370 77716
rect 32493 77707 32551 77713
rect 32493 77704 32505 77707
rect 32364 77676 32505 77704
rect 32364 77664 32370 77676
rect 32493 77673 32505 77676
rect 32539 77673 32551 77707
rect 32493 77667 32551 77673
rect 32950 77664 32956 77716
rect 33008 77704 33014 77716
rect 33689 77707 33747 77713
rect 33689 77704 33701 77707
rect 33008 77676 33701 77704
rect 33008 77664 33014 77676
rect 33689 77673 33701 77676
rect 33735 77673 33747 77707
rect 33689 77667 33747 77673
rect 33962 77664 33968 77716
rect 34020 77664 34026 77716
rect 34698 77664 34704 77716
rect 34756 77664 34762 77716
rect 34790 77664 34796 77716
rect 34848 77704 34854 77716
rect 34885 77707 34943 77713
rect 34885 77704 34897 77707
rect 34848 77676 34897 77704
rect 34848 77664 34854 77676
rect 34885 77673 34897 77676
rect 34931 77673 34943 77707
rect 34885 77667 34943 77673
rect 35250 77664 35256 77716
rect 35308 77704 35314 77716
rect 35805 77707 35863 77713
rect 35805 77704 35817 77707
rect 35308 77676 35817 77704
rect 35308 77664 35314 77676
rect 35805 77673 35817 77676
rect 35851 77704 35863 77707
rect 40678 77704 40684 77716
rect 35851 77676 40684 77704
rect 35851 77673 35863 77676
rect 35805 77667 35863 77673
rect 40678 77664 40684 77676
rect 40736 77664 40742 77716
rect 70213 77707 70271 77713
rect 55186 77676 68876 77704
rect 24670 77596 24676 77648
rect 24728 77596 24734 77648
rect 24762 77596 24768 77648
rect 24820 77636 24826 77648
rect 24857 77639 24915 77645
rect 24857 77636 24869 77639
rect 24820 77608 24869 77636
rect 24820 77596 24826 77608
rect 24857 77605 24869 77608
rect 24903 77605 24915 77639
rect 24857 77599 24915 77605
rect 25038 77596 25044 77648
rect 25096 77596 25102 77648
rect 26786 77596 26792 77648
rect 26844 77636 26850 77648
rect 27249 77639 27307 77645
rect 27249 77636 27261 77639
rect 26844 77608 27261 77636
rect 26844 77596 26850 77608
rect 27249 77605 27261 77608
rect 27295 77605 27307 77639
rect 31680 77636 31708 77664
rect 27249 77599 27307 77605
rect 31128 77608 31708 77636
rect 32140 77608 33272 77636
rect 20806 77392 20812 77444
rect 20864 77392 20870 77444
rect 21266 77392 21272 77444
rect 21324 77392 21330 77444
rect 16117 77367 16175 77373
rect 16117 77364 16129 77367
rect 16080 77336 16129 77364
rect 16080 77324 16086 77336
rect 16117 77333 16129 77336
rect 16163 77364 16175 77367
rect 19613 77367 19671 77373
rect 19613 77364 19625 77367
rect 16163 77336 19625 77364
rect 16163 77333 16175 77336
rect 16117 77327 16175 77333
rect 19613 77333 19625 77336
rect 19659 77333 19671 77367
rect 19613 77327 19671 77333
rect 21358 77324 21364 77376
rect 21416 77364 21422 77376
rect 24213 77367 24271 77373
rect 24213 77364 24225 77367
rect 21416 77336 24225 77364
rect 21416 77324 21422 77336
rect 24213 77333 24225 77336
rect 24259 77364 24271 77367
rect 24397 77367 24455 77373
rect 24397 77364 24409 77367
rect 24259 77336 24409 77364
rect 24259 77333 24271 77336
rect 24213 77327 24271 77333
rect 24397 77333 24409 77336
rect 24443 77333 24455 77367
rect 25056 77364 25084 77596
rect 26786 77460 26792 77512
rect 26844 77500 26850 77512
rect 31128 77509 31156 77608
rect 31202 77528 31208 77580
rect 31260 77528 31266 77580
rect 32140 77577 32168 77608
rect 31389 77571 31447 77577
rect 31389 77537 31401 77571
rect 31435 77568 31447 77571
rect 32125 77571 32183 77577
rect 32125 77568 32137 77571
rect 31435 77540 32137 77568
rect 31435 77537 31447 77540
rect 31389 77531 31447 77537
rect 32125 77537 32137 77540
rect 32171 77537 32183 77571
rect 32125 77531 32183 77537
rect 32950 77528 32956 77580
rect 33008 77568 33014 77580
rect 33244 77577 33272 77608
rect 38654 77596 38660 77648
rect 38712 77596 38718 77648
rect 39669 77639 39727 77645
rect 39669 77605 39681 77639
rect 39715 77636 39727 77639
rect 39758 77636 39764 77648
rect 39715 77608 39764 77636
rect 39715 77605 39727 77608
rect 39669 77599 39727 77605
rect 39758 77596 39764 77608
rect 39816 77596 39822 77648
rect 39850 77596 39856 77648
rect 39908 77596 39914 77648
rect 40144 77608 40540 77636
rect 33137 77571 33195 77577
rect 33137 77568 33149 77571
rect 33008 77540 33149 77568
rect 33008 77528 33014 77540
rect 33137 77537 33149 77540
rect 33183 77537 33195 77571
rect 33137 77531 33195 77537
rect 33229 77571 33287 77577
rect 33229 77537 33241 77571
rect 33275 77568 33287 77571
rect 34149 77571 34207 77577
rect 34149 77568 34161 77571
rect 33275 77540 34161 77568
rect 33275 77537 33287 77540
rect 33229 77531 33287 77537
rect 34149 77537 34161 77540
rect 34195 77568 34207 77571
rect 35437 77571 35495 77577
rect 35437 77568 35449 77571
rect 34195 77540 35449 77568
rect 34195 77537 34207 77540
rect 34149 77531 34207 77537
rect 35437 77537 35449 77540
rect 35483 77568 35495 77571
rect 36081 77571 36139 77577
rect 36081 77568 36093 77571
rect 35483 77540 36093 77568
rect 35483 77537 35495 77540
rect 35437 77531 35495 77537
rect 36081 77537 36093 77540
rect 36127 77568 36139 77571
rect 37829 77571 37887 77577
rect 37829 77568 37841 77571
rect 36127 77540 37841 77568
rect 36127 77537 36139 77540
rect 36081 77531 36139 77537
rect 37829 77537 37841 77540
rect 37875 77568 37887 77571
rect 38473 77571 38531 77577
rect 38473 77568 38485 77571
rect 37875 77540 38485 77568
rect 37875 77537 37887 77540
rect 37829 77531 37887 77537
rect 38473 77537 38485 77540
rect 38519 77568 38531 77571
rect 40144 77568 40172 77608
rect 40512 77577 40540 77608
rect 40862 77596 40868 77648
rect 40920 77596 40926 77648
rect 40954 77596 40960 77648
rect 41012 77636 41018 77648
rect 41233 77639 41291 77645
rect 41233 77636 41245 77639
rect 41012 77608 41245 77636
rect 41012 77596 41018 77608
rect 41233 77605 41245 77608
rect 41279 77605 41291 77639
rect 41233 77599 41291 77605
rect 42150 77596 42156 77648
rect 42208 77596 42214 77648
rect 43717 77639 43775 77645
rect 43717 77636 43729 77639
rect 43088 77608 43729 77636
rect 43088 77577 43116 77608
rect 43717 77605 43729 77608
rect 43763 77636 43775 77639
rect 55186 77636 55214 77676
rect 43763 77608 55214 77636
rect 43763 77605 43775 77608
rect 43717 77599 43775 77605
rect 62482 77596 62488 77648
rect 62540 77596 62546 77648
rect 63773 77639 63831 77645
rect 63144 77608 63448 77636
rect 38519 77540 40172 77568
rect 40497 77571 40555 77577
rect 38519 77537 38531 77540
rect 38473 77531 38531 77537
rect 40497 77537 40509 77571
rect 40543 77568 40555 77571
rect 41141 77571 41199 77577
rect 41141 77568 41153 77571
rect 40543 77540 41153 77568
rect 40543 77537 40555 77540
rect 40497 77531 40555 77537
rect 41141 77537 41153 77540
rect 41187 77568 41199 77571
rect 43073 77571 43131 77577
rect 43073 77568 43085 77571
rect 41187 77540 43085 77568
rect 41187 77537 41199 77540
rect 41141 77531 41199 77537
rect 43073 77537 43085 77540
rect 43119 77537 43131 77571
rect 43073 77531 43131 77537
rect 43806 77528 43812 77580
rect 43864 77528 43870 77580
rect 63144 77577 63172 77608
rect 61013 77571 61071 77577
rect 61013 77537 61025 77571
rect 61059 77568 61071 77571
rect 61841 77571 61899 77577
rect 61841 77568 61853 77571
rect 61059 77540 61853 77568
rect 61059 77537 61071 77540
rect 61013 77531 61071 77537
rect 61841 77537 61853 77540
rect 61887 77568 61899 77571
rect 63129 77571 63187 77577
rect 63129 77568 63141 77571
rect 61887 77540 63141 77568
rect 61887 77537 61899 77540
rect 61841 77531 61899 77537
rect 63129 77537 63141 77540
rect 63175 77537 63187 77571
rect 63420 77568 63448 77608
rect 63773 77605 63785 77639
rect 63819 77636 63831 77639
rect 63954 77636 63960 77648
rect 63819 77608 63960 77636
rect 63819 77605 63831 77608
rect 63773 77599 63831 77605
rect 63954 77596 63960 77608
rect 64012 77596 64018 77648
rect 64966 77596 64972 77648
rect 65024 77636 65030 77648
rect 65024 77608 65748 77636
rect 65024 77596 65030 77608
rect 64046 77568 64052 77580
rect 63420 77540 64052 77568
rect 63129 77531 63187 77537
rect 64046 77528 64052 77540
rect 64104 77528 64110 77580
rect 64138 77528 64144 77580
rect 64196 77568 64202 77580
rect 65720 77577 65748 77608
rect 67634 77596 67640 77648
rect 67692 77636 67698 77648
rect 67692 77608 68600 77636
rect 67692 77596 67698 77608
rect 65705 77571 65763 77577
rect 64196 77540 65196 77568
rect 64196 77528 64202 77540
rect 27065 77503 27123 77509
rect 27065 77500 27077 77503
rect 26844 77472 27077 77500
rect 26844 77460 26850 77472
rect 27065 77469 27077 77472
rect 27111 77469 27123 77503
rect 27065 77463 27123 77469
rect 31113 77503 31171 77509
rect 31113 77469 31125 77503
rect 31159 77469 31171 77503
rect 31220 77500 31248 77528
rect 31757 77503 31815 77509
rect 31757 77500 31769 77503
rect 31220 77472 31769 77500
rect 31113 77463 31171 77469
rect 31757 77469 31769 77472
rect 31803 77469 31815 77503
rect 31757 77463 31815 77469
rect 35250 77460 35256 77512
rect 35308 77460 35314 77512
rect 35342 77460 35348 77512
rect 35400 77500 35406 77512
rect 35897 77503 35955 77509
rect 35897 77500 35909 77503
rect 35400 77472 35909 77500
rect 35400 77460 35406 77472
rect 35897 77469 35909 77472
rect 35943 77469 35955 77503
rect 35897 77463 35955 77469
rect 36262 77460 36268 77512
rect 36320 77500 36326 77512
rect 36357 77503 36415 77509
rect 36357 77500 36369 77503
rect 36320 77472 36369 77500
rect 36320 77460 36326 77472
rect 36357 77469 36369 77472
rect 36403 77469 36415 77503
rect 36357 77463 36415 77469
rect 36998 77460 37004 77512
rect 37056 77460 37062 77512
rect 37645 77503 37703 77509
rect 37645 77469 37657 77503
rect 37691 77500 37703 77503
rect 38197 77503 38255 77509
rect 38197 77500 38209 77503
rect 37691 77472 38209 77500
rect 37691 77469 37703 77472
rect 37645 77463 37703 77469
rect 38197 77469 38209 77472
rect 38243 77500 38255 77503
rect 40034 77500 40040 77512
rect 38243 77472 40040 77500
rect 38243 77469 38255 77472
rect 38197 77463 38255 77469
rect 40034 77460 40040 77472
rect 40092 77460 40098 77512
rect 40773 77503 40831 77509
rect 40773 77500 40785 77503
rect 40328 77472 40785 77500
rect 26050 77392 26056 77444
rect 26108 77392 26114 77444
rect 26513 77435 26571 77441
rect 26513 77401 26525 77435
rect 26559 77432 26571 77435
rect 39942 77432 39948 77444
rect 26559 77404 39948 77432
rect 26559 77401 26571 77404
rect 26513 77395 26571 77401
rect 39942 77392 39948 77404
rect 40000 77392 40006 77444
rect 40221 77435 40279 77441
rect 40221 77401 40233 77435
rect 40267 77432 40279 77435
rect 40328 77432 40356 77472
rect 40773 77469 40785 77472
rect 40819 77500 40831 77503
rect 46106 77500 46112 77512
rect 40819 77472 46112 77500
rect 40819 77469 40831 77472
rect 40773 77463 40831 77469
rect 46106 77460 46112 77472
rect 46164 77460 46170 77512
rect 60553 77503 60611 77509
rect 60553 77469 60565 77503
rect 60599 77500 60611 77503
rect 61102 77500 61108 77512
rect 60599 77472 61108 77500
rect 60599 77469 60611 77472
rect 60553 77463 60611 77469
rect 61102 77460 61108 77472
rect 61160 77460 61166 77512
rect 62761 77503 62819 77509
rect 62761 77469 62773 77503
rect 62807 77500 62819 77503
rect 63310 77500 63316 77512
rect 62807 77472 63316 77500
rect 62807 77469 62819 77472
rect 62761 77463 62819 77469
rect 63310 77460 63316 77472
rect 63368 77460 63374 77512
rect 63512 77472 65104 77500
rect 40267 77404 40356 77432
rect 42797 77435 42855 77441
rect 40267 77401 40279 77404
rect 40221 77395 40279 77401
rect 42797 77401 42809 77435
rect 42843 77432 42855 77435
rect 43349 77435 43407 77441
rect 43349 77432 43361 77435
rect 42843 77404 43361 77432
rect 42843 77401 42855 77404
rect 42797 77395 42855 77401
rect 43349 77401 43361 77404
rect 43395 77432 43407 77435
rect 48590 77432 48596 77444
rect 43395 77404 48596 77432
rect 43395 77401 43407 77404
rect 43349 77395 43407 77401
rect 48590 77392 48596 77404
rect 48648 77392 48654 77444
rect 51074 77392 51080 77444
rect 51132 77432 51138 77444
rect 60737 77435 60795 77441
rect 60737 77432 60749 77435
rect 51132 77404 60749 77432
rect 51132 77392 51138 77404
rect 60737 77401 60749 77404
rect 60783 77432 60795 77435
rect 61197 77435 61255 77441
rect 61197 77432 61209 77435
rect 60783 77404 61209 77432
rect 60783 77401 60795 77404
rect 60737 77395 60795 77401
rect 61197 77401 61209 77404
rect 61243 77401 61255 77435
rect 61197 77395 61255 77401
rect 62482 77392 62488 77444
rect 62540 77432 62546 77444
rect 63405 77435 63463 77441
rect 63405 77432 63417 77435
rect 62540 77404 63417 77432
rect 62540 77392 62546 77404
rect 63405 77401 63417 77404
rect 63451 77401 63463 77435
rect 63405 77395 63463 77401
rect 27433 77367 27491 77373
rect 27433 77364 27445 77367
rect 25056 77336 27445 77364
rect 24397 77327 24455 77333
rect 27433 77333 27445 77336
rect 27479 77333 27491 77367
rect 27433 77327 27491 77333
rect 31570 77324 31576 77376
rect 31628 77364 31634 77376
rect 32309 77367 32367 77373
rect 32309 77364 32321 77367
rect 31628 77336 32321 77364
rect 31628 77324 31634 77336
rect 32309 77333 32321 77336
rect 32355 77333 32367 77367
rect 32309 77327 32367 77333
rect 32674 77324 32680 77376
rect 32732 77324 32738 77376
rect 33045 77367 33103 77373
rect 33045 77333 33057 77367
rect 33091 77364 33103 77367
rect 33597 77367 33655 77373
rect 33597 77364 33609 77367
rect 33091 77336 33609 77364
rect 33091 77333 33103 77336
rect 33045 77327 33103 77333
rect 33597 77333 33609 77336
rect 33643 77364 33655 77367
rect 35986 77364 35992 77376
rect 33643 77336 35992 77364
rect 33643 77333 33655 77336
rect 33597 77327 33655 77333
rect 35986 77324 35992 77336
rect 36044 77324 36050 77376
rect 37274 77324 37280 77376
rect 37332 77324 37338 77376
rect 37734 77324 37740 77376
rect 37792 77364 37798 77376
rect 38289 77367 38347 77373
rect 38289 77364 38301 77367
rect 37792 77336 38301 77364
rect 37792 77324 37798 77336
rect 38289 77333 38301 77336
rect 38335 77333 38347 77367
rect 38289 77327 38347 77333
rect 40126 77324 40132 77376
rect 40184 77364 40190 77376
rect 40313 77367 40371 77373
rect 40313 77364 40325 77367
rect 40184 77336 40325 77364
rect 40184 77324 40190 77336
rect 40313 77333 40325 77336
rect 40359 77333 40371 77367
rect 40313 77327 40371 77333
rect 42426 77324 42432 77376
rect 42484 77324 42490 77376
rect 42886 77324 42892 77376
rect 42944 77364 42950 77376
rect 43441 77367 43499 77373
rect 43441 77364 43453 77367
rect 42944 77336 43453 77364
rect 42944 77324 42950 77336
rect 43441 77333 43453 77336
rect 43487 77333 43499 77367
rect 43441 77327 43499 77333
rect 61565 77367 61623 77373
rect 61565 77333 61577 77367
rect 61611 77364 61623 77367
rect 61749 77367 61807 77373
rect 61749 77364 61761 77367
rect 61611 77336 61761 77364
rect 61611 77333 61623 77336
rect 61565 77327 61623 77333
rect 61749 77333 61761 77336
rect 61795 77364 61807 77367
rect 63512 77364 63540 77472
rect 61795 77336 63540 77364
rect 61795 77333 61807 77336
rect 61749 77327 61807 77333
rect 64046 77324 64052 77376
rect 64104 77364 64110 77376
rect 64966 77364 64972 77376
rect 64104 77336 64972 77364
rect 64104 77324 64110 77336
rect 64966 77324 64972 77336
rect 65024 77324 65030 77376
rect 65076 77364 65104 77472
rect 65168 77441 65196 77540
rect 65705 77537 65717 77571
rect 65751 77568 65763 77571
rect 66625 77571 66683 77577
rect 66625 77568 66637 77571
rect 65751 77540 66637 77568
rect 65751 77537 65763 77540
rect 65705 77531 65763 77537
rect 66625 77537 66637 77540
rect 66671 77568 66683 77571
rect 68278 77568 68284 77580
rect 66671 77540 68284 77568
rect 66671 77537 66683 77540
rect 66625 77531 66683 77537
rect 68278 77528 68284 77540
rect 68336 77528 68342 77580
rect 68462 77528 68468 77580
rect 68520 77528 68526 77580
rect 65337 77503 65395 77509
rect 65337 77469 65349 77503
rect 65383 77500 65395 77503
rect 65886 77500 65892 77512
rect 65383 77472 65892 77500
rect 65383 77469 65395 77472
rect 65337 77463 65395 77469
rect 65886 77460 65892 77472
rect 65944 77460 65950 77512
rect 67358 77500 67364 77512
rect 66088 77472 67364 77500
rect 65153 77435 65211 77441
rect 65153 77401 65165 77435
rect 65199 77432 65211 77435
rect 65981 77435 66039 77441
rect 65981 77432 65993 77435
rect 65199 77404 65993 77432
rect 65199 77401 65211 77404
rect 65153 77395 65211 77401
rect 65981 77401 65993 77404
rect 66027 77401 66039 77435
rect 65981 77395 66039 77401
rect 66088 77364 66116 77472
rect 67358 77460 67364 77472
rect 67416 77460 67422 77512
rect 67913 77503 67971 77509
rect 67913 77469 67925 77503
rect 67959 77500 67971 77503
rect 68480 77500 68508 77528
rect 68572 77509 68600 77608
rect 67959 77472 68508 77500
rect 68557 77503 68615 77509
rect 67959 77469 67971 77472
rect 67913 77463 67971 77469
rect 68557 77469 68569 77503
rect 68603 77469 68615 77503
rect 68848 77500 68876 77676
rect 69584 77676 69796 77704
rect 68925 77639 68983 77645
rect 68925 77605 68937 77639
rect 68971 77636 68983 77639
rect 69106 77636 69112 77648
rect 68971 77608 69112 77636
rect 68971 77605 68983 77608
rect 68925 77599 68983 77605
rect 69106 77596 69112 77608
rect 69164 77596 69170 77648
rect 69198 77528 69204 77580
rect 69256 77568 69262 77580
rect 69584 77577 69612 77676
rect 69768 77636 69796 77676
rect 70213 77673 70225 77707
rect 70259 77704 70271 77707
rect 70394 77704 70400 77716
rect 70259 77676 70400 77704
rect 70259 77673 70271 77676
rect 70213 77667 70271 77673
rect 70394 77664 70400 77676
rect 70452 77664 70458 77716
rect 70946 77664 70952 77716
rect 71004 77664 71010 77716
rect 71038 77664 71044 77716
rect 71096 77704 71102 77716
rect 71096 77676 71728 77704
rect 71096 77664 71102 77676
rect 70489 77639 70547 77645
rect 70489 77636 70501 77639
rect 69768 77608 70501 77636
rect 70489 77605 70501 77608
rect 70535 77605 70547 77639
rect 70489 77599 70547 77605
rect 69569 77571 69627 77577
rect 69569 77568 69581 77571
rect 69256 77540 69581 77568
rect 69256 77528 69262 77540
rect 69569 77537 69581 77540
rect 69615 77537 69627 77571
rect 69569 77531 69627 77537
rect 69750 77528 69756 77580
rect 69808 77528 69814 77580
rect 70504 77568 70532 77599
rect 71130 77596 71136 77648
rect 71188 77596 71194 77648
rect 71700 77636 71728 77676
rect 71958 77664 71964 77716
rect 72016 77664 72022 77716
rect 72068 77676 74120 77704
rect 72068 77636 72096 77676
rect 73433 77639 73491 77645
rect 71700 77608 72096 77636
rect 73264 77608 73384 77636
rect 71317 77571 71375 77577
rect 71317 77568 71329 77571
rect 70504 77540 71329 77568
rect 71317 77537 71329 77540
rect 71363 77568 71375 77571
rect 72053 77571 72111 77577
rect 72053 77568 72065 77571
rect 71363 77540 72065 77568
rect 71363 77537 71375 77540
rect 71317 77531 71375 77537
rect 72053 77537 72065 77540
rect 72099 77568 72111 77571
rect 73264 77568 73292 77608
rect 72099 77540 73292 77568
rect 73356 77568 73384 77608
rect 73433 77605 73445 77639
rect 73479 77636 73491 77639
rect 74092 77636 74120 77676
rect 74442 77664 74448 77716
rect 74500 77664 74506 77716
rect 76650 77664 76656 77716
rect 76708 77664 76714 77716
rect 78217 77707 78275 77713
rect 78217 77673 78229 77707
rect 78263 77704 78275 77707
rect 78766 77704 78772 77716
rect 78263 77676 78772 77704
rect 78263 77673 78275 77676
rect 78217 77667 78275 77673
rect 78766 77664 78772 77676
rect 78824 77664 78830 77716
rect 79226 77664 79232 77716
rect 79284 77664 79290 77716
rect 80054 77664 80060 77716
rect 80112 77664 80118 77716
rect 103790 77704 103796 77716
rect 80440 77676 83320 77704
rect 77757 77639 77815 77645
rect 77757 77636 77769 77639
rect 73479 77608 74028 77636
rect 74092 77608 77769 77636
rect 73479 77605 73491 77608
rect 73433 77599 73491 77605
rect 74000 77580 74028 77608
rect 77757 77605 77769 77608
rect 77803 77636 77815 77639
rect 79873 77639 79931 77645
rect 77803 77608 78904 77636
rect 77803 77605 77815 77608
rect 77757 77599 77815 77605
rect 73798 77568 73804 77580
rect 73356 77540 73804 77568
rect 72099 77537 72111 77540
rect 72053 77531 72111 77537
rect 73798 77528 73804 77540
rect 73856 77528 73862 77580
rect 73982 77528 73988 77580
rect 74040 77528 74046 77580
rect 76101 77571 76159 77577
rect 76101 77537 76113 77571
rect 76147 77537 76159 77571
rect 76101 77531 76159 77537
rect 74626 77500 74632 77512
rect 68848 77472 74632 77500
rect 68557 77463 68615 77469
rect 74626 77460 74632 77472
rect 74684 77500 74690 77512
rect 75457 77503 75515 77509
rect 75457 77500 75469 77503
rect 74684 77472 75469 77500
rect 74684 77460 74690 77472
rect 75457 77469 75469 77472
rect 75503 77469 75515 77503
rect 75457 77463 75515 77469
rect 66533 77435 66591 77441
rect 66533 77432 66545 77435
rect 66364 77404 66545 77432
rect 66364 77373 66392 77404
rect 66533 77401 66545 77404
rect 66579 77432 66591 77435
rect 71314 77432 71320 77444
rect 66579 77404 71320 77432
rect 66579 77401 66591 77404
rect 66533 77395 66591 77401
rect 71314 77392 71320 77404
rect 71372 77392 71378 77444
rect 71593 77435 71651 77441
rect 71593 77432 71605 77435
rect 71424 77404 71605 77432
rect 65076 77336 66116 77364
rect 66349 77367 66407 77373
rect 66349 77333 66361 77367
rect 66395 77333 66407 77367
rect 66349 77327 66407 77333
rect 68278 77324 68284 77376
rect 68336 77364 68342 77376
rect 69198 77364 69204 77376
rect 68336 77336 69204 77364
rect 68336 77324 68342 77336
rect 69198 77324 69204 77336
rect 69256 77324 69262 77376
rect 69293 77367 69351 77373
rect 69293 77333 69305 77367
rect 69339 77364 69351 77367
rect 69750 77364 69756 77376
rect 69339 77336 69756 77364
rect 69339 77333 69351 77336
rect 69293 77327 69351 77333
rect 69750 77324 69756 77336
rect 69808 77324 69814 77376
rect 69842 77324 69848 77376
rect 69900 77324 69906 77376
rect 71130 77324 71136 77376
rect 71188 77364 71194 77376
rect 71424 77364 71452 77404
rect 71593 77401 71605 77404
rect 71639 77401 71651 77435
rect 71593 77395 71651 77401
rect 73430 77392 73436 77444
rect 73488 77432 73494 77444
rect 73525 77435 73583 77441
rect 73525 77432 73537 77435
rect 73488 77404 73537 77432
rect 73488 77392 73494 77404
rect 73525 77401 73537 77404
rect 73571 77432 73583 77435
rect 74077 77435 74135 77441
rect 74077 77432 74089 77435
rect 73571 77404 74089 77432
rect 73571 77401 73583 77404
rect 73525 77395 73583 77401
rect 74077 77401 74089 77404
rect 74123 77401 74135 77435
rect 74997 77435 75055 77441
rect 74997 77432 75009 77435
rect 74077 77395 74135 77401
rect 74506 77404 75009 77432
rect 71188 77336 71452 77364
rect 71501 77367 71559 77373
rect 71188 77324 71194 77336
rect 71501 77333 71513 77367
rect 71547 77364 71559 77367
rect 71682 77364 71688 77376
rect 71547 77336 71688 77364
rect 71547 77333 71559 77336
rect 71501 77327 71559 77333
rect 71682 77324 71688 77336
rect 71740 77324 71746 77376
rect 73798 77324 73804 77376
rect 73856 77364 73862 77376
rect 74506 77364 74534 77404
rect 74997 77401 75009 77404
rect 75043 77432 75055 77435
rect 75181 77435 75239 77441
rect 75181 77432 75193 77435
rect 75043 77404 75193 77432
rect 75043 77401 75055 77404
rect 74997 77395 75055 77401
rect 75181 77401 75193 77404
rect 75227 77432 75239 77435
rect 75365 77435 75423 77441
rect 75365 77432 75377 77435
rect 75227 77404 75377 77432
rect 75227 77401 75239 77404
rect 75181 77395 75239 77401
rect 75365 77401 75377 77404
rect 75411 77432 75423 77435
rect 75733 77435 75791 77441
rect 75733 77432 75745 77435
rect 75411 77404 75745 77432
rect 75411 77401 75423 77404
rect 75365 77395 75423 77401
rect 75733 77401 75745 77404
rect 75779 77432 75791 77435
rect 76116 77432 76144 77531
rect 76190 77528 76196 77580
rect 76248 77528 76254 77580
rect 78677 77571 78735 77577
rect 78677 77537 78689 77571
rect 78723 77537 78735 77571
rect 78677 77531 78735 77537
rect 78033 77435 78091 77441
rect 78033 77432 78045 77435
rect 75779 77404 78045 77432
rect 75779 77401 75791 77404
rect 75733 77395 75791 77401
rect 78033 77401 78045 77404
rect 78079 77432 78091 77435
rect 78692 77432 78720 77531
rect 78766 77528 78772 77580
rect 78824 77528 78830 77580
rect 78876 77509 78904 77608
rect 79873 77605 79885 77639
rect 79919 77636 79931 77639
rect 80440 77636 80468 77676
rect 79919 77608 80468 77636
rect 79919 77605 79931 77608
rect 79873 77599 79931 77605
rect 80440 77577 80468 77608
rect 80882 77596 80888 77648
rect 80940 77596 80946 77648
rect 83292 77636 83320 77676
rect 84166 77676 103796 77704
rect 84166 77636 84194 77676
rect 103790 77664 103796 77676
rect 103848 77664 103854 77716
rect 83292 77608 84194 77636
rect 86586 77596 86592 77648
rect 86644 77636 86650 77648
rect 87322 77636 87328 77648
rect 86644 77608 87328 77636
rect 86644 77596 86650 77608
rect 87322 77596 87328 77608
rect 87380 77596 87386 77648
rect 90545 77639 90603 77645
rect 90545 77605 90557 77639
rect 90591 77636 90603 77639
rect 90726 77636 90732 77648
rect 90591 77608 90732 77636
rect 90591 77605 90603 77608
rect 90545 77599 90603 77605
rect 90726 77596 90732 77608
rect 90784 77596 90790 77648
rect 93118 77596 93124 77648
rect 93176 77596 93182 77648
rect 95697 77639 95755 77645
rect 95697 77605 95709 77639
rect 95743 77636 95755 77639
rect 95743 77608 99604 77636
rect 95743 77605 95755 77608
rect 95697 77599 95755 77605
rect 79689 77571 79747 77577
rect 79689 77537 79701 77571
rect 79735 77568 79747 77571
rect 80241 77571 80299 77577
rect 80241 77568 80253 77571
rect 79735 77540 80253 77568
rect 79735 77537 79747 77540
rect 79689 77531 79747 77537
rect 80241 77537 80253 77540
rect 80287 77537 80299 77571
rect 80241 77531 80299 77537
rect 80425 77571 80483 77577
rect 80425 77537 80437 77571
rect 80471 77537 80483 77571
rect 80425 77531 80483 77537
rect 81621 77571 81679 77577
rect 81621 77537 81633 77571
rect 81667 77568 81679 77571
rect 85669 77571 85727 77577
rect 81667 77540 83872 77568
rect 81667 77537 81679 77540
rect 81621 77531 81679 77537
rect 78861 77503 78919 77509
rect 78861 77469 78873 77503
rect 78907 77469 78919 77503
rect 78861 77463 78919 77469
rect 79704 77432 79732 77531
rect 83844 77512 83872 77540
rect 85669 77537 85681 77571
rect 85715 77568 85727 77571
rect 86221 77571 86279 77577
rect 86221 77568 86233 77571
rect 85715 77540 86233 77568
rect 85715 77537 85727 77540
rect 85669 77531 85727 77537
rect 86221 77537 86233 77540
rect 86267 77537 86279 77571
rect 86221 77531 86279 77537
rect 86494 77528 86500 77580
rect 86552 77528 86558 77580
rect 89070 77528 89076 77580
rect 89128 77568 89134 77580
rect 93949 77571 94007 77577
rect 93949 77568 93961 77571
rect 89128 77540 93961 77568
rect 89128 77528 89134 77540
rect 93949 77537 93961 77540
rect 93995 77568 94007 77571
rect 95789 77571 95847 77577
rect 95789 77568 95801 77571
rect 93995 77540 95801 77568
rect 93995 77537 94007 77540
rect 93949 77531 94007 77537
rect 95789 77537 95801 77540
rect 95835 77537 95847 77571
rect 95789 77531 95847 77537
rect 80054 77460 80060 77512
rect 80112 77500 80118 77512
rect 80517 77503 80575 77509
rect 80517 77500 80529 77503
rect 80112 77472 80529 77500
rect 80112 77460 80118 77472
rect 80517 77469 80529 77472
rect 80563 77469 80575 77503
rect 80517 77463 80575 77469
rect 83369 77503 83427 77509
rect 83369 77469 83381 77503
rect 83415 77500 83427 77503
rect 83415 77472 83688 77500
rect 83415 77469 83427 77472
rect 83369 77463 83427 77469
rect 78079 77404 79732 77432
rect 78079 77401 78091 77404
rect 78033 77395 78091 77401
rect 81526 77392 81532 77444
rect 81584 77432 81590 77444
rect 81584 77404 81926 77432
rect 81584 77392 81590 77404
rect 83090 77392 83096 77444
rect 83148 77392 83154 77444
rect 83660 77376 83688 77472
rect 83826 77460 83832 77512
rect 83884 77460 83890 77512
rect 85945 77503 86003 77509
rect 85945 77469 85957 77503
rect 85991 77469 86003 77503
rect 85945 77463 86003 77469
rect 84286 77392 84292 77444
rect 84344 77432 84350 77444
rect 85960 77432 85988 77463
rect 86402 77460 86408 77512
rect 86460 77500 86466 77512
rect 86589 77503 86647 77509
rect 86589 77500 86601 77503
rect 86460 77472 86601 77500
rect 86460 77460 86466 77472
rect 86589 77469 86601 77472
rect 86635 77469 86647 77503
rect 86589 77463 86647 77469
rect 86862 77460 86868 77512
rect 86920 77500 86926 77512
rect 88797 77503 88855 77509
rect 88797 77500 88809 77503
rect 86920 77472 88809 77500
rect 86920 77460 86926 77472
rect 88797 77469 88809 77472
rect 88843 77469 88855 77503
rect 88797 77463 88855 77469
rect 91373 77503 91431 77509
rect 91373 77469 91385 77503
rect 91419 77469 91431 77503
rect 91373 77463 91431 77469
rect 86880 77432 86908 77460
rect 84344 77404 84502 77432
rect 85960 77404 86908 77432
rect 86957 77435 87015 77441
rect 84344 77392 84350 77404
rect 86957 77401 86969 77435
rect 87003 77401 87015 77435
rect 86957 77395 87015 77401
rect 87141 77435 87199 77441
rect 87141 77401 87153 77435
rect 87187 77432 87199 77435
rect 87230 77432 87236 77444
rect 87187 77404 87236 77432
rect 87187 77401 87199 77404
rect 87141 77395 87199 77401
rect 73856 77336 74534 77364
rect 73856 77324 73862 77336
rect 75638 77324 75644 77376
rect 75696 77364 75702 77376
rect 76190 77364 76196 77376
rect 75696 77336 76196 77364
rect 75696 77324 75702 77336
rect 76190 77324 76196 77336
rect 76248 77324 76254 77376
rect 76282 77324 76288 77376
rect 76340 77324 76346 77376
rect 83642 77324 83648 77376
rect 83700 77324 83706 77376
rect 84010 77324 84016 77376
rect 84068 77324 84074 77376
rect 84197 77367 84255 77373
rect 84197 77333 84209 77367
rect 84243 77364 84255 77367
rect 86494 77364 86500 77376
rect 84243 77336 86500 77364
rect 84243 77333 84255 77336
rect 84197 77327 84255 77333
rect 86494 77324 86500 77336
rect 86552 77364 86558 77376
rect 86972 77364 87000 77395
rect 87230 77392 87236 77404
rect 87288 77392 87294 77444
rect 86552 77336 87000 77364
rect 88812 77364 88840 77463
rect 88978 77392 88984 77444
rect 89036 77432 89042 77444
rect 89073 77435 89131 77441
rect 89073 77432 89085 77435
rect 89036 77404 89085 77432
rect 89036 77392 89042 77404
rect 89073 77401 89085 77404
rect 89119 77401 89131 77435
rect 89073 77395 89131 77401
rect 89714 77392 89720 77444
rect 89772 77392 89778 77444
rect 90376 77404 90956 77432
rect 89438 77364 89444 77376
rect 88812 77336 89444 77364
rect 86552 77324 86558 77336
rect 89438 77324 89444 77336
rect 89496 77364 89502 77376
rect 90376 77364 90404 77404
rect 90928 77373 90956 77404
rect 89496 77336 90404 77364
rect 90913 77367 90971 77373
rect 89496 77324 89502 77336
rect 90913 77333 90925 77367
rect 90959 77364 90971 77367
rect 91388 77364 91416 77463
rect 91646 77392 91652 77444
rect 91704 77392 91710 77444
rect 92658 77392 92664 77444
rect 92716 77392 92722 77444
rect 92952 77404 93348 77432
rect 92014 77364 92020 77376
rect 90959 77336 92020 77364
rect 90959 77333 90971 77336
rect 90913 77327 90971 77333
rect 92014 77324 92020 77336
rect 92072 77364 92078 77376
rect 92952 77364 92980 77404
rect 93320 77373 93348 77404
rect 94222 77392 94228 77444
rect 94280 77392 94286 77444
rect 95234 77392 95240 77444
rect 95292 77392 95298 77444
rect 99576 77432 99604 77608
rect 99650 77528 99656 77580
rect 99708 77568 99714 77580
rect 108114 77568 108120 77580
rect 99708 77540 108120 77568
rect 99708 77528 99714 77540
rect 108114 77528 108120 77540
rect 108172 77528 108178 77580
rect 106274 77432 106280 77444
rect 95620 77404 95924 77432
rect 99576 77404 106280 77432
rect 92072 77336 92980 77364
rect 93305 77367 93363 77373
rect 92072 77324 92078 77336
rect 93305 77333 93317 77367
rect 93351 77364 93363 77367
rect 95620 77364 95648 77404
rect 93351 77336 95648 77364
rect 95896 77364 95924 77404
rect 106274 77392 106280 77404
rect 106332 77392 106338 77444
rect 104158 77364 104164 77376
rect 95896 77336 104164 77364
rect 93351 77333 93363 77336
rect 93305 77327 93363 77333
rect 104158 77324 104164 77336
rect 104216 77324 104222 77376
rect 1104 77274 108836 77296
rect 1104 77222 4874 77274
rect 4926 77222 4938 77274
rect 4990 77222 5002 77274
rect 5054 77222 5066 77274
rect 5118 77222 5130 77274
rect 5182 77222 35594 77274
rect 35646 77222 35658 77274
rect 35710 77222 35722 77274
rect 35774 77222 35786 77274
rect 35838 77222 35850 77274
rect 35902 77222 66314 77274
rect 66366 77222 66378 77274
rect 66430 77222 66442 77274
rect 66494 77222 66506 77274
rect 66558 77222 66570 77274
rect 66622 77222 97034 77274
rect 97086 77222 97098 77274
rect 97150 77222 97162 77274
rect 97214 77222 97226 77274
rect 97278 77222 97290 77274
rect 97342 77222 106658 77274
rect 106710 77222 106722 77274
rect 106774 77222 106786 77274
rect 106838 77222 106850 77274
rect 106902 77222 106914 77274
rect 106966 77222 108836 77274
rect 1104 77200 108836 77222
rect 1762 77120 1768 77172
rect 1820 77160 1826 77172
rect 23474 77160 23480 77172
rect 1820 77132 23480 77160
rect 1820 77120 1826 77132
rect 23474 77120 23480 77132
rect 23532 77120 23538 77172
rect 27246 77120 27252 77172
rect 27304 77160 27310 77172
rect 27617 77163 27675 77169
rect 27617 77160 27629 77163
rect 27304 77132 27629 77160
rect 27304 77120 27310 77132
rect 27617 77129 27629 77132
rect 27663 77129 27675 77163
rect 27617 77123 27675 77129
rect 68554 77120 68560 77172
rect 68612 77160 68618 77172
rect 75825 77163 75883 77169
rect 75825 77160 75837 77163
rect 68612 77132 75837 77160
rect 68612 77120 68618 77132
rect 75825 77129 75837 77132
rect 75871 77160 75883 77163
rect 76282 77160 76288 77172
rect 75871 77132 76288 77160
rect 75871 77129 75883 77132
rect 75825 77123 75883 77129
rect 76282 77120 76288 77132
rect 76340 77120 76346 77172
rect 81526 77120 81532 77172
rect 81584 77120 81590 77172
rect 83090 77120 83096 77172
rect 83148 77160 83154 77172
rect 83921 77163 83979 77169
rect 83921 77160 83933 77163
rect 83148 77132 83933 77160
rect 83148 77120 83154 77132
rect 83921 77129 83933 77132
rect 83967 77129 83979 77163
rect 88426 77160 88432 77172
rect 83921 77123 83979 77129
rect 85408 77132 88432 77160
rect 24762 77092 24768 77104
rect 23874 77064 24768 77092
rect 24762 77052 24768 77064
rect 24820 77052 24826 77104
rect 27430 77092 27436 77104
rect 25714 77064 27436 77092
rect 27430 77052 27436 77064
rect 27488 77052 27494 77104
rect 27522 77052 27528 77104
rect 27580 77092 27586 77104
rect 30285 77095 30343 77101
rect 30285 77092 30297 77095
rect 27580 77064 30297 77092
rect 27580 77052 27586 77064
rect 30285 77061 30297 77064
rect 30331 77061 30343 77095
rect 30285 77055 30343 77061
rect 69198 77052 69204 77104
rect 69256 77052 69262 77104
rect 75638 77052 75644 77104
rect 75696 77052 75702 77104
rect 1210 76984 1216 77036
rect 1268 77024 1274 77036
rect 1489 77027 1547 77033
rect 1489 77024 1501 77027
rect 1268 76996 1501 77024
rect 1268 76984 1274 76996
rect 1489 76993 1501 76996
rect 1535 77024 1547 77027
rect 1949 77027 2007 77033
rect 1949 77024 1961 77027
rect 1535 76996 1961 77024
rect 1535 76993 1547 76996
rect 1489 76987 1547 76993
rect 1949 76993 1961 76996
rect 1995 76993 2007 77027
rect 1949 76987 2007 76993
rect 26421 77027 26479 77033
rect 26421 76993 26433 77027
rect 26467 77024 26479 77027
rect 26786 77024 26792 77036
rect 26467 76996 26792 77024
rect 26467 76993 26479 76996
rect 26421 76987 26479 76993
rect 26786 76984 26792 76996
rect 26844 76984 26850 77036
rect 27709 77027 27767 77033
rect 27709 76993 27721 77027
rect 27755 77024 27767 77027
rect 27893 77027 27951 77033
rect 27893 77024 27905 77027
rect 27755 76996 27905 77024
rect 27755 76993 27767 76996
rect 27709 76987 27767 76993
rect 27893 76993 27905 76996
rect 27939 77024 27951 77027
rect 30377 77027 30435 77033
rect 30377 77024 30389 77027
rect 27939 76996 30389 77024
rect 27939 76993 27951 76996
rect 27893 76987 27951 76993
rect 30377 76993 30389 76996
rect 30423 77024 30435 77027
rect 81621 77027 81679 77033
rect 30423 76996 30604 77024
rect 30423 76993 30435 76996
rect 30377 76987 30435 76993
rect 22741 76959 22799 76965
rect 22741 76925 22753 76959
rect 22787 76956 22799 76959
rect 24302 76956 24308 76968
rect 22787 76928 24308 76956
rect 22787 76925 22799 76928
rect 22741 76919 22799 76925
rect 24302 76916 24308 76928
rect 24360 76916 24366 76968
rect 24578 76916 24584 76968
rect 24636 76916 24642 76968
rect 26145 76959 26203 76965
rect 26145 76925 26157 76959
rect 26191 76956 26203 76959
rect 30466 76956 30472 76968
rect 26191 76928 30472 76956
rect 26191 76925 26203 76928
rect 26145 76919 26203 76925
rect 30466 76916 30472 76928
rect 30524 76916 30530 76968
rect 1673 76891 1731 76897
rect 1673 76857 1685 76891
rect 1719 76888 1731 76891
rect 1857 76891 1915 76897
rect 1857 76888 1869 76891
rect 1719 76860 1869 76888
rect 1719 76857 1731 76860
rect 1673 76851 1731 76857
rect 1857 76857 1869 76860
rect 1903 76888 1915 76891
rect 1903 76860 6914 76888
rect 1903 76857 1915 76860
rect 1857 76851 1915 76857
rect 6886 76820 6914 76860
rect 22002 76848 22008 76900
rect 22060 76888 22066 76900
rect 22060 76860 22968 76888
rect 22060 76848 22066 76860
rect 22094 76820 22100 76832
rect 6886 76792 22100 76820
rect 22094 76780 22100 76792
rect 22152 76780 22158 76832
rect 22830 76780 22836 76832
rect 22888 76780 22894 76832
rect 22940 76820 22968 76860
rect 30576 76832 30604 76996
rect 81621 76993 81633 77027
rect 81667 77024 81679 77027
rect 81667 76996 81848 77024
rect 81667 76993 81679 76996
rect 81621 76987 81679 76993
rect 69385 76891 69443 76897
rect 69385 76888 69397 76891
rect 64846 76860 69397 76888
rect 24673 76823 24731 76829
rect 24673 76820 24685 76823
rect 22940 76792 24685 76820
rect 24673 76789 24685 76792
rect 24719 76820 24731 76823
rect 26513 76823 26571 76829
rect 26513 76820 26525 76823
rect 24719 76792 26525 76820
rect 24719 76789 24731 76792
rect 24673 76783 24731 76789
rect 26513 76789 26525 76792
rect 26559 76789 26571 76823
rect 26513 76783 26571 76789
rect 26786 76780 26792 76832
rect 26844 76780 26850 76832
rect 30558 76780 30564 76832
rect 30616 76780 30622 76832
rect 61102 76780 61108 76832
rect 61160 76820 61166 76832
rect 64846 76820 64874 76860
rect 69385 76857 69397 76860
rect 69431 76888 69443 76891
rect 69842 76888 69848 76900
rect 69431 76860 69848 76888
rect 69431 76857 69443 76860
rect 69385 76851 69443 76857
rect 69842 76848 69848 76860
rect 69900 76848 69906 76900
rect 81820 76829 81848 76996
rect 83826 76984 83832 77036
rect 83884 77024 83890 77036
rect 84013 77027 84071 77033
rect 84013 77024 84025 77027
rect 83884 76996 84025 77024
rect 83884 76984 83890 76996
rect 84013 76993 84025 76996
rect 84059 77024 84071 77027
rect 84105 77027 84163 77033
rect 84105 77024 84117 77027
rect 84059 76996 84117 77024
rect 84059 76993 84071 76996
rect 84013 76987 84071 76993
rect 84105 76993 84117 76996
rect 84151 76993 84163 77027
rect 84105 76987 84163 76993
rect 83918 76916 83924 76968
rect 83976 76956 83982 76968
rect 85408 76956 85436 77132
rect 88426 77120 88432 77132
rect 88484 77120 88490 77172
rect 88613 77163 88671 77169
rect 88613 77129 88625 77163
rect 88659 77160 88671 77163
rect 88886 77160 88892 77172
rect 88659 77132 88892 77160
rect 88659 77129 88671 77132
rect 88613 77123 88671 77129
rect 88886 77120 88892 77132
rect 88944 77120 88950 77172
rect 92014 77120 92020 77172
rect 92072 77120 92078 77172
rect 85758 77052 85764 77104
rect 85816 77092 85822 77104
rect 85816 77064 87630 77092
rect 85816 77052 85822 77064
rect 88518 77052 88524 77104
rect 88576 77092 88582 77104
rect 91741 77095 91799 77101
rect 88576 77064 90206 77092
rect 88576 77052 88582 77064
rect 91741 77061 91753 77095
rect 91787 77092 91799 77095
rect 95234 77092 95240 77104
rect 91787 77064 95240 77092
rect 91787 77061 91799 77064
rect 91741 77055 91799 77061
rect 95234 77052 95240 77064
rect 95292 77052 95298 77104
rect 85574 76984 85580 77036
rect 85632 77024 85638 77036
rect 85945 77027 86003 77033
rect 85945 77024 85957 77027
rect 85632 76996 85957 77024
rect 85632 76984 85638 76996
rect 85945 76993 85957 76996
rect 85991 77024 86003 77027
rect 86402 77024 86408 77036
rect 85991 76996 86408 77024
rect 85991 76993 86003 76996
rect 85945 76987 86003 76993
rect 86402 76984 86408 76996
rect 86460 76984 86466 77036
rect 86494 76984 86500 77036
rect 86552 77024 86558 77036
rect 86589 77027 86647 77033
rect 86589 77024 86601 77027
rect 86552 76996 86601 77024
rect 86552 76984 86558 76996
rect 86589 76993 86601 76996
rect 86635 76993 86647 77027
rect 86589 76987 86647 76993
rect 86773 77027 86831 77033
rect 86773 76993 86785 77027
rect 86819 77024 86831 77027
rect 86862 77024 86868 77036
rect 86819 76996 86868 77024
rect 86819 76993 86831 76996
rect 86773 76987 86831 76993
rect 86862 76984 86868 76996
rect 86920 76984 86926 77036
rect 88978 76984 88984 77036
rect 89036 77024 89042 77036
rect 89073 77027 89131 77033
rect 89073 77024 89085 77027
rect 89036 76996 89085 77024
rect 89036 76984 89042 76996
rect 89073 76993 89085 76996
rect 89119 77024 89131 77027
rect 89438 77024 89444 77036
rect 89119 76996 89444 77024
rect 89119 76993 89131 76996
rect 89073 76987 89131 76993
rect 89438 76984 89444 76996
rect 89496 76984 89502 77036
rect 91462 76984 91468 77036
rect 91520 77024 91526 77036
rect 91649 77027 91707 77033
rect 91649 77024 91661 77027
rect 91520 76996 91661 77024
rect 91520 76984 91526 76996
rect 91649 76993 91661 76996
rect 91695 76993 91707 77027
rect 91649 76987 91707 76993
rect 106274 76984 106280 77036
rect 106332 77024 106338 77036
rect 108301 77027 108359 77033
rect 108301 77024 108313 77027
rect 106332 76996 108313 77024
rect 106332 76984 106338 76996
rect 108301 76993 108313 76996
rect 108347 76993 108359 77027
rect 108301 76987 108359 76993
rect 83976 76928 85436 76956
rect 83976 76916 83982 76928
rect 85666 76916 85672 76968
rect 85724 76956 85730 76968
rect 87141 76959 87199 76965
rect 87141 76956 87153 76959
rect 85724 76928 87153 76956
rect 85724 76916 85730 76928
rect 87141 76925 87153 76928
rect 87187 76925 87199 76959
rect 87141 76919 87199 76925
rect 89717 76959 89775 76965
rect 89717 76925 89729 76959
rect 89763 76956 89775 76959
rect 89806 76956 89812 76968
rect 89763 76928 89812 76956
rect 89763 76925 89775 76928
rect 89717 76919 89775 76925
rect 89806 76916 89812 76928
rect 89864 76916 89870 76968
rect 86770 76888 86776 76900
rect 84166 76860 86776 76888
rect 61160 76792 64874 76820
rect 81805 76823 81863 76829
rect 61160 76780 61166 76792
rect 81805 76789 81817 76823
rect 81851 76820 81863 76823
rect 82814 76820 82820 76832
rect 81851 76792 82820 76820
rect 81851 76789 81863 76792
rect 81805 76783 81863 76789
rect 82814 76780 82820 76792
rect 82872 76780 82878 76832
rect 84010 76780 84016 76832
rect 84068 76820 84074 76832
rect 84166 76820 84194 76860
rect 86770 76848 86776 76860
rect 86828 76848 86834 76900
rect 91189 76891 91247 76897
rect 91189 76857 91201 76891
rect 91235 76888 91247 76891
rect 91373 76891 91431 76897
rect 91373 76888 91385 76891
rect 91235 76860 91385 76888
rect 91235 76857 91247 76860
rect 91189 76851 91247 76857
rect 91373 76857 91385 76860
rect 91419 76888 91431 76891
rect 105814 76888 105820 76900
rect 91419 76860 105820 76888
rect 91419 76857 91431 76860
rect 91373 76851 91431 76857
rect 105814 76848 105820 76860
rect 105872 76848 105878 76900
rect 108482 76848 108488 76900
rect 108540 76848 108546 76900
rect 84068 76792 84194 76820
rect 84289 76823 84347 76829
rect 84068 76780 84074 76792
rect 84289 76789 84301 76823
rect 84335 76820 84347 76823
rect 85574 76820 85580 76832
rect 84335 76792 85580 76820
rect 84335 76789 84347 76792
rect 84289 76783 84347 76789
rect 85574 76780 85580 76792
rect 85632 76780 85638 76832
rect 85853 76823 85911 76829
rect 85853 76789 85865 76823
rect 85899 76820 85911 76823
rect 86126 76820 86132 76832
rect 85899 76792 86132 76820
rect 85899 76789 85911 76792
rect 85853 76783 85911 76789
rect 86126 76780 86132 76792
rect 86184 76780 86190 76832
rect 86405 76823 86463 76829
rect 86405 76789 86417 76823
rect 86451 76820 86463 76823
rect 86586 76820 86592 76832
rect 86451 76792 86592 76820
rect 86451 76789 86463 76792
rect 86405 76783 86463 76789
rect 86586 76780 86592 76792
rect 86644 76780 86650 76832
rect 87230 76780 87236 76832
rect 87288 76820 87294 76832
rect 89898 76820 89904 76832
rect 87288 76792 89904 76820
rect 87288 76780 87294 76792
rect 89898 76780 89904 76792
rect 89956 76780 89962 76832
rect 91462 76780 91468 76832
rect 91520 76780 91526 76832
rect 1104 76730 108836 76752
rect 1104 76678 4214 76730
rect 4266 76678 4278 76730
rect 4330 76678 4342 76730
rect 4394 76678 4406 76730
rect 4458 76678 4470 76730
rect 4522 76678 34934 76730
rect 34986 76678 34998 76730
rect 35050 76678 35062 76730
rect 35114 76678 35126 76730
rect 35178 76678 35190 76730
rect 35242 76678 65654 76730
rect 65706 76678 65718 76730
rect 65770 76678 65782 76730
rect 65834 76678 65846 76730
rect 65898 76678 65910 76730
rect 65962 76678 96374 76730
rect 96426 76678 96438 76730
rect 96490 76678 96502 76730
rect 96554 76678 96566 76730
rect 96618 76678 96630 76730
rect 96682 76678 108836 76730
rect 1104 76656 108836 76678
rect 21542 76576 21548 76628
rect 21600 76576 21606 76628
rect 23474 76576 23480 76628
rect 23532 76616 23538 76628
rect 23569 76619 23627 76625
rect 23569 76616 23581 76619
rect 23532 76588 23581 76616
rect 23532 76576 23538 76588
rect 23569 76585 23581 76588
rect 23615 76585 23627 76619
rect 23569 76579 23627 76585
rect 24578 76576 24584 76628
rect 24636 76616 24642 76628
rect 24949 76619 25007 76625
rect 24949 76616 24961 76619
rect 24636 76588 24961 76616
rect 24636 76576 24642 76588
rect 24949 76585 24961 76588
rect 24995 76616 25007 76619
rect 26786 76616 26792 76628
rect 24995 76588 26792 76616
rect 24995 76585 25007 76588
rect 24949 76579 25007 76585
rect 26786 76576 26792 76588
rect 26844 76576 26850 76628
rect 27430 76576 27436 76628
rect 27488 76616 27494 76628
rect 31573 76619 31631 76625
rect 31573 76616 31585 76619
rect 27488 76588 31585 76616
rect 27488 76576 27494 76588
rect 31573 76585 31585 76588
rect 31619 76585 31631 76619
rect 31573 76579 31631 76585
rect 82817 76619 82875 76625
rect 82817 76585 82829 76619
rect 82863 76616 82875 76619
rect 84286 76616 84292 76628
rect 82863 76588 84292 76616
rect 82863 76585 82875 76588
rect 82817 76579 82875 76585
rect 84286 76576 84292 76588
rect 84344 76576 84350 76628
rect 85758 76576 85764 76628
rect 85816 76576 85822 76628
rect 85942 76576 85948 76628
rect 86000 76576 86006 76628
rect 86126 76576 86132 76628
rect 86184 76616 86190 76628
rect 86184 76588 88104 76616
rect 86184 76576 86190 76588
rect 21560 76480 21588 76576
rect 23014 76508 23020 76560
rect 23072 76548 23078 76560
rect 24673 76551 24731 76557
rect 24673 76548 24685 76551
rect 23072 76520 24685 76548
rect 23072 76508 23078 76520
rect 24673 76517 24685 76520
rect 24719 76517 24731 76551
rect 24673 76511 24731 76517
rect 24762 76508 24768 76560
rect 24820 76548 24826 76560
rect 31021 76551 31079 76557
rect 31021 76548 31033 76551
rect 24820 76520 31033 76548
rect 24820 76508 24826 76520
rect 31021 76517 31033 76520
rect 31067 76517 31079 76551
rect 31021 76511 31079 76517
rect 21729 76483 21787 76489
rect 21729 76480 21741 76483
rect 21560 76452 21741 76480
rect 21729 76449 21741 76452
rect 21775 76449 21787 76483
rect 21729 76443 21787 76449
rect 22005 76483 22063 76489
rect 22005 76449 22017 76483
rect 22051 76480 22063 76483
rect 32674 76480 32680 76492
rect 22051 76452 32680 76480
rect 22051 76449 22063 76452
rect 22005 76443 22063 76449
rect 32674 76440 32680 76452
rect 32732 76440 32738 76492
rect 83001 76483 83059 76489
rect 83001 76449 83013 76483
rect 83047 76480 83059 76483
rect 83642 76480 83648 76492
rect 83047 76452 83648 76480
rect 83047 76449 83059 76452
rect 83001 76443 83059 76449
rect 83642 76440 83648 76452
rect 83700 76480 83706 76492
rect 85117 76483 85175 76489
rect 85117 76480 85129 76483
rect 83700 76452 85129 76480
rect 83700 76440 83706 76452
rect 85117 76449 85129 76452
rect 85163 76480 85175 76483
rect 86221 76483 86279 76489
rect 86221 76480 86233 76483
rect 85163 76452 86233 76480
rect 85163 76449 85175 76452
rect 85117 76443 85175 76449
rect 86221 76449 86233 76452
rect 86267 76480 86279 76483
rect 86862 76480 86868 76492
rect 86267 76452 86868 76480
rect 86267 76449 86279 76452
rect 86221 76443 86279 76449
rect 86862 76440 86868 76452
rect 86920 76440 86926 76492
rect 88076 76480 88104 76588
rect 88518 76576 88524 76628
rect 88576 76576 88582 76628
rect 88978 76576 88984 76628
rect 89036 76576 89042 76628
rect 89809 76619 89867 76625
rect 89809 76585 89821 76619
rect 89855 76616 89867 76619
rect 92658 76616 92664 76628
rect 89855 76588 92664 76616
rect 89855 76585 89867 76588
rect 89809 76579 89867 76585
rect 92658 76576 92664 76588
rect 92716 76576 92722 76628
rect 88153 76551 88211 76557
rect 88153 76517 88165 76551
rect 88199 76548 88211 76551
rect 89714 76548 89720 76560
rect 88199 76520 89720 76548
rect 88199 76517 88211 76520
rect 88153 76511 88211 76517
rect 89714 76508 89720 76520
rect 89772 76508 89778 76560
rect 102226 76480 102232 76492
rect 88076 76452 102232 76480
rect 102226 76440 102232 76452
rect 102284 76440 102290 76492
rect 1581 76415 1639 76421
rect 1581 76381 1593 76415
rect 1627 76412 1639 76415
rect 1765 76415 1823 76421
rect 1765 76412 1777 76415
rect 1627 76384 1777 76412
rect 1627 76381 1639 76384
rect 1581 76375 1639 76381
rect 1765 76381 1777 76384
rect 1811 76412 1823 76415
rect 17862 76412 17868 76424
rect 1811 76384 17868 76412
rect 1811 76381 1823 76384
rect 1765 76375 1823 76381
rect 17862 76372 17868 76384
rect 17920 76372 17926 76424
rect 29089 76415 29147 76421
rect 29089 76381 29101 76415
rect 29135 76412 29147 76415
rect 29273 76415 29331 76421
rect 29273 76412 29285 76415
rect 29135 76384 29285 76412
rect 29135 76381 29147 76384
rect 29089 76375 29147 76381
rect 29273 76381 29285 76384
rect 29319 76412 29331 76415
rect 30558 76412 30564 76424
rect 29319 76384 30564 76412
rect 29319 76381 29331 76384
rect 29273 76375 29331 76381
rect 30558 76372 30564 76384
rect 30616 76412 30622 76424
rect 31113 76415 31171 76421
rect 31113 76412 31125 76415
rect 30616 76384 31125 76412
rect 30616 76372 30622 76384
rect 31113 76381 31125 76384
rect 31159 76412 31171 76415
rect 31297 76415 31355 76421
rect 31297 76412 31309 76415
rect 31159 76384 31309 76412
rect 31159 76381 31171 76384
rect 31113 76375 31171 76381
rect 31297 76381 31309 76384
rect 31343 76412 31355 76415
rect 31665 76415 31723 76421
rect 31665 76412 31677 76415
rect 31343 76384 31677 76412
rect 31343 76381 31355 76384
rect 31297 76375 31355 76381
rect 31665 76381 31677 76384
rect 31711 76412 31723 76415
rect 31849 76415 31907 76421
rect 31849 76412 31861 76415
rect 31711 76384 31861 76412
rect 31711 76381 31723 76384
rect 31665 76375 31723 76381
rect 31849 76381 31861 76384
rect 31895 76412 31907 76415
rect 32401 76415 32459 76421
rect 32401 76412 32413 76415
rect 31895 76384 32413 76412
rect 31895 76381 31907 76384
rect 31849 76375 31907 76381
rect 32401 76381 32413 76384
rect 32447 76412 32459 76415
rect 82265 76415 82323 76421
rect 32447 76384 32628 76412
rect 32447 76381 32459 76384
rect 32401 76375 32459 76381
rect 28997 76347 29055 76353
rect 28997 76344 29009 76347
rect 23230 76316 29009 76344
rect 28997 76313 29009 76316
rect 29043 76313 29055 76347
rect 28997 76307 29055 76313
rect 30282 76304 30288 76356
rect 30340 76344 30346 76356
rect 32309 76347 32367 76353
rect 32309 76344 32321 76347
rect 30340 76316 32321 76344
rect 30340 76304 30346 76316
rect 32309 76313 32321 76316
rect 32355 76313 32367 76347
rect 32309 76307 32367 76313
rect 842 76236 848 76288
rect 900 76276 906 76288
rect 32600 76285 32628 76384
rect 82265 76381 82277 76415
rect 82311 76412 82323 76415
rect 82357 76415 82415 76421
rect 82357 76412 82369 76415
rect 82311 76384 82369 76412
rect 82311 76381 82323 76384
rect 82265 76375 82323 76381
rect 82357 76381 82369 76384
rect 82403 76412 82415 76415
rect 82725 76415 82783 76421
rect 82725 76412 82737 76415
rect 82403 76384 82737 76412
rect 82403 76381 82415 76384
rect 82357 76375 82415 76381
rect 82725 76381 82737 76384
rect 82771 76412 82783 76415
rect 82814 76412 82820 76424
rect 82771 76384 82820 76412
rect 82771 76381 82783 76384
rect 82725 76375 82783 76381
rect 82814 76372 82820 76384
rect 82872 76372 82878 76424
rect 85669 76415 85727 76421
rect 85669 76381 85681 76415
rect 85715 76412 85727 76415
rect 88061 76415 88119 76421
rect 88061 76412 88073 76415
rect 85715 76384 86264 76412
rect 85715 76381 85727 76384
rect 85669 76375 85727 76381
rect 82449 76347 82507 76353
rect 82449 76313 82461 76347
rect 82495 76344 82507 76347
rect 82495 76316 83136 76344
rect 82495 76313 82507 76316
rect 82449 76307 82507 76313
rect 1397 76279 1455 76285
rect 1397 76276 1409 76279
rect 900 76248 1409 76276
rect 900 76236 906 76248
rect 1397 76245 1409 76248
rect 1443 76245 1455 76279
rect 1397 76239 1455 76245
rect 32585 76279 32643 76285
rect 32585 76245 32597 76279
rect 32631 76276 32643 76279
rect 73982 76276 73988 76288
rect 32631 76248 73988 76276
rect 32631 76245 32643 76248
rect 32585 76239 32643 76245
rect 73982 76236 73988 76248
rect 74040 76236 74046 76288
rect 83108 76276 83136 76316
rect 83274 76304 83280 76356
rect 83332 76304 83338 76356
rect 83384 76316 83766 76344
rect 83384 76276 83412 76316
rect 83108 76248 83412 76276
rect 84749 76279 84807 76285
rect 84749 76245 84761 76279
rect 84795 76276 84807 76279
rect 84933 76279 84991 76285
rect 84933 76276 84945 76279
rect 84795 76248 84945 76276
rect 84795 76245 84807 76248
rect 84749 76239 84807 76245
rect 84933 76245 84945 76248
rect 84979 76276 84991 76279
rect 85574 76276 85580 76288
rect 84979 76248 85580 76276
rect 84979 76245 84991 76248
rect 84933 76239 84991 76245
rect 85574 76236 85580 76248
rect 85632 76236 85638 76288
rect 86236 76276 86264 76384
rect 87800 76384 88073 76412
rect 86402 76304 86408 76356
rect 86460 76344 86466 76356
rect 86497 76347 86555 76353
rect 86497 76344 86509 76347
rect 86460 76316 86509 76344
rect 86460 76304 86466 76316
rect 86497 76313 86509 76316
rect 86543 76313 86555 76347
rect 86497 76307 86555 76313
rect 86954 76304 86960 76356
rect 87012 76304 87018 76356
rect 87138 76276 87144 76288
rect 86236 76248 87144 76276
rect 87138 76236 87144 76248
rect 87196 76276 87202 76288
rect 87800 76276 87828 76384
rect 88061 76381 88073 76384
rect 88107 76381 88119 76415
rect 88061 76375 88119 76381
rect 88426 76372 88432 76424
rect 88484 76412 88490 76424
rect 89162 76412 89168 76424
rect 88484 76384 89168 76412
rect 88484 76372 88490 76384
rect 89162 76372 89168 76384
rect 89220 76372 89226 76424
rect 89714 76372 89720 76424
rect 89772 76372 89778 76424
rect 107654 76372 107660 76424
rect 107712 76412 107718 76424
rect 108301 76415 108359 76421
rect 108301 76412 108313 76415
rect 107712 76384 108313 76412
rect 107712 76372 107718 76384
rect 108301 76381 108313 76384
rect 108347 76381 108359 76415
rect 108301 76375 108359 76381
rect 88797 76347 88855 76353
rect 88797 76344 88809 76347
rect 87984 76316 88809 76344
rect 87984 76285 88012 76316
rect 88797 76313 88809 76316
rect 88843 76344 88855 76347
rect 108114 76344 108120 76356
rect 88843 76316 108120 76344
rect 88843 76313 88855 76316
rect 88797 76307 88855 76313
rect 108114 76304 108120 76316
rect 108172 76304 108178 76356
rect 87196 76248 87828 76276
rect 87969 76279 88027 76285
rect 87196 76236 87202 76248
rect 87969 76245 87981 76279
rect 88015 76245 88027 76279
rect 87969 76239 88027 76245
rect 89162 76236 89168 76288
rect 89220 76276 89226 76288
rect 89714 76276 89720 76288
rect 89220 76248 89720 76276
rect 89220 76236 89226 76248
rect 89714 76236 89720 76248
rect 89772 76276 89778 76288
rect 89993 76279 90051 76285
rect 89993 76276 90005 76279
rect 89772 76248 90005 76276
rect 89772 76236 89778 76248
rect 89993 76245 90005 76248
rect 90039 76276 90051 76279
rect 91462 76276 91468 76288
rect 90039 76248 91468 76276
rect 90039 76245 90051 76248
rect 89993 76239 90051 76245
rect 91462 76236 91468 76248
rect 91520 76236 91526 76288
rect 108482 76236 108488 76288
rect 108540 76236 108546 76288
rect 1104 76186 108836 76208
rect 1104 76134 4874 76186
rect 4926 76134 4938 76186
rect 4990 76134 5002 76186
rect 5054 76134 5066 76186
rect 5118 76134 5130 76186
rect 5182 76134 35594 76186
rect 35646 76134 35658 76186
rect 35710 76134 35722 76186
rect 35774 76134 35786 76186
rect 35838 76134 35850 76186
rect 35902 76134 66314 76186
rect 66366 76134 66378 76186
rect 66430 76134 66442 76186
rect 66494 76134 66506 76186
rect 66558 76134 66570 76186
rect 66622 76134 97034 76186
rect 97086 76134 97098 76186
rect 97150 76134 97162 76186
rect 97214 76134 97226 76186
rect 97278 76134 97290 76186
rect 97342 76134 108836 76186
rect 1104 76112 108836 76134
rect 1765 76075 1823 76081
rect 1765 76041 1777 76075
rect 1811 76072 1823 76075
rect 2314 76072 2320 76084
rect 1811 76044 2320 76072
rect 1811 76041 1823 76044
rect 1765 76035 1823 76041
rect 1581 75939 1639 75945
rect 1581 75905 1593 75939
rect 1627 75936 1639 75939
rect 1780 75936 1808 76035
rect 2314 76032 2320 76044
rect 2372 76032 2378 76084
rect 82814 76032 82820 76084
rect 82872 76072 82878 76084
rect 83093 76075 83151 76081
rect 83093 76072 83105 76075
rect 82872 76044 83105 76072
rect 82872 76032 82878 76044
rect 83093 76041 83105 76044
rect 83139 76072 83151 76075
rect 83918 76072 83924 76084
rect 83139 76044 83924 76072
rect 83139 76041 83151 76044
rect 83093 76035 83151 76041
rect 24302 75964 24308 76016
rect 24360 76004 24366 76016
rect 37274 76004 37280 76016
rect 24360 75976 37280 76004
rect 24360 75964 24366 75976
rect 37274 75964 37280 75976
rect 37332 75964 37338 76016
rect 81342 75964 81348 76016
rect 81400 76004 81406 76016
rect 82909 76007 82967 76013
rect 82909 76004 82921 76007
rect 81400 75976 82921 76004
rect 81400 75964 81406 75976
rect 82909 75973 82921 75976
rect 82955 76004 82967 76007
rect 83274 76004 83280 76016
rect 82955 75976 83280 76004
rect 82955 75973 82967 75976
rect 82909 75967 82967 75973
rect 83274 75964 83280 75976
rect 83332 75964 83338 76016
rect 83660 75945 83688 76044
rect 83918 76032 83924 76044
rect 83976 76032 83982 76084
rect 84286 76032 84292 76084
rect 84344 76072 84350 76084
rect 86678 76072 86684 76084
rect 84344 76044 86684 76072
rect 84344 76032 84350 76044
rect 86678 76032 86684 76044
rect 86736 76032 86742 76084
rect 86770 76032 86776 76084
rect 86828 76072 86834 76084
rect 90085 76075 90143 76081
rect 90085 76072 90097 76075
rect 86828 76044 90097 76072
rect 86828 76032 86834 76044
rect 90085 76041 90097 76044
rect 90131 76041 90143 76075
rect 90085 76035 90143 76041
rect 83737 76007 83795 76013
rect 83737 75973 83749 76007
rect 83783 76004 83795 76007
rect 86405 76007 86463 76013
rect 83783 75976 85054 76004
rect 83783 75973 83795 75976
rect 83737 75967 83795 75973
rect 86405 75973 86417 76007
rect 86451 76004 86463 76007
rect 87230 76004 87236 76016
rect 86451 75976 87236 76004
rect 86451 75973 86463 75976
rect 86405 75967 86463 75973
rect 87230 75964 87236 75976
rect 87288 75964 87294 76016
rect 87414 75964 87420 76016
rect 87472 75964 87478 76016
rect 1627 75908 1808 75936
rect 83645 75939 83703 75945
rect 1627 75905 1639 75908
rect 1581 75899 1639 75905
rect 83645 75905 83657 75939
rect 83691 75905 83703 75939
rect 83645 75899 83703 75905
rect 84286 75896 84292 75948
rect 84344 75896 84350 75948
rect 89898 75896 89904 75948
rect 89956 75936 89962 75948
rect 89993 75939 90051 75945
rect 89993 75936 90005 75939
rect 89956 75908 90005 75936
rect 89956 75896 89962 75908
rect 89993 75905 90005 75908
rect 90039 75905 90051 75939
rect 90100 75936 90128 76035
rect 108114 76032 108120 76084
rect 108172 76032 108178 76084
rect 108482 76032 108488 76084
rect 108540 76032 108546 76084
rect 90269 76007 90327 76013
rect 90269 75973 90281 76007
rect 90315 76004 90327 76007
rect 90315 75976 90772 76004
rect 90315 75973 90327 75976
rect 90269 75967 90327 75973
rect 90744 75948 90772 75976
rect 90361 75939 90419 75945
rect 90361 75936 90373 75939
rect 90100 75908 90373 75936
rect 89993 75899 90051 75905
rect 90361 75905 90373 75908
rect 90407 75905 90419 75939
rect 90361 75899 90419 75905
rect 90726 75896 90732 75948
rect 90784 75936 90790 75948
rect 90821 75939 90879 75945
rect 90821 75936 90833 75939
rect 90784 75908 90833 75936
rect 90784 75896 90790 75908
rect 90821 75905 90833 75908
rect 90867 75905 90879 75939
rect 108132 75936 108160 76032
rect 108301 75939 108359 75945
rect 108301 75936 108313 75939
rect 108132 75908 108313 75936
rect 90821 75899 90879 75905
rect 108301 75905 108313 75908
rect 108347 75905 108359 75939
rect 108301 75899 108359 75905
rect 71774 75828 71780 75880
rect 71832 75868 71838 75880
rect 84197 75871 84255 75877
rect 84197 75868 84209 75871
rect 71832 75840 84209 75868
rect 71832 75828 71838 75840
rect 84197 75837 84209 75840
rect 84243 75868 84255 75871
rect 84565 75871 84623 75877
rect 84565 75868 84577 75871
rect 84243 75840 84577 75868
rect 84243 75837 84255 75840
rect 84197 75831 84255 75837
rect 84565 75837 84577 75840
rect 84611 75837 84623 75871
rect 84565 75831 84623 75837
rect 86678 75828 86684 75880
rect 86736 75828 86742 75880
rect 86957 75871 87015 75877
rect 86957 75837 86969 75871
rect 87003 75868 87015 75871
rect 87046 75868 87052 75880
rect 87003 75840 87052 75868
rect 87003 75837 87015 75840
rect 86957 75831 87015 75837
rect 87046 75828 87052 75840
rect 87104 75828 87110 75880
rect 88702 75828 88708 75880
rect 88760 75868 88766 75880
rect 88889 75871 88947 75877
rect 88889 75868 88901 75871
rect 88760 75840 88901 75868
rect 88760 75828 88766 75840
rect 88889 75837 88901 75840
rect 88935 75868 88947 75871
rect 89070 75868 89076 75880
rect 88935 75840 89076 75868
rect 88935 75837 88947 75840
rect 88889 75831 88947 75837
rect 89070 75828 89076 75840
rect 89128 75828 89134 75880
rect 86037 75803 86095 75809
rect 86037 75769 86049 75803
rect 86083 75800 86095 75803
rect 86586 75800 86592 75812
rect 86083 75772 86592 75800
rect 86083 75769 86095 75772
rect 86037 75763 86095 75769
rect 86586 75760 86592 75772
rect 86644 75760 86650 75812
rect 88429 75803 88487 75809
rect 88429 75769 88441 75803
rect 88475 75800 88487 75803
rect 88613 75803 88671 75809
rect 88613 75800 88625 75803
rect 88475 75772 88625 75800
rect 88475 75769 88487 75772
rect 88429 75763 88487 75769
rect 88613 75769 88625 75772
rect 88659 75800 88671 75803
rect 91005 75803 91063 75809
rect 88659 75772 90680 75800
rect 88659 75769 88671 75772
rect 88613 75763 88671 75769
rect 1394 75692 1400 75744
rect 1452 75692 1458 75744
rect 86310 75692 86316 75744
rect 86368 75692 86374 75744
rect 90174 75692 90180 75744
rect 90232 75732 90238 75744
rect 90269 75735 90327 75741
rect 90269 75732 90281 75735
rect 90232 75704 90281 75732
rect 90232 75692 90238 75704
rect 90269 75701 90281 75704
rect 90315 75701 90327 75735
rect 90269 75695 90327 75701
rect 90450 75692 90456 75744
rect 90508 75732 90514 75744
rect 90545 75735 90603 75741
rect 90545 75732 90557 75735
rect 90508 75704 90557 75732
rect 90508 75692 90514 75704
rect 90545 75701 90557 75704
rect 90591 75701 90603 75735
rect 90652 75732 90680 75772
rect 91005 75769 91017 75803
rect 91051 75800 91063 75803
rect 91189 75803 91247 75809
rect 91189 75800 91201 75803
rect 91051 75772 91201 75800
rect 91051 75769 91063 75772
rect 91005 75763 91063 75769
rect 91189 75769 91201 75772
rect 91235 75800 91247 75803
rect 102686 75800 102692 75812
rect 91235 75772 102692 75800
rect 91235 75769 91247 75772
rect 91189 75763 91247 75769
rect 102686 75760 102692 75772
rect 102744 75760 102750 75812
rect 108114 75732 108120 75744
rect 90652 75704 108120 75732
rect 90545 75695 90603 75701
rect 108114 75692 108120 75704
rect 108172 75692 108178 75744
rect 1104 75642 108836 75664
rect 1104 75590 4214 75642
rect 4266 75590 4278 75642
rect 4330 75590 4342 75642
rect 4394 75590 4406 75642
rect 4458 75590 4470 75642
rect 4522 75590 34934 75642
rect 34986 75590 34998 75642
rect 35050 75590 35062 75642
rect 35114 75590 35126 75642
rect 35178 75590 35190 75642
rect 35242 75590 65654 75642
rect 65706 75590 65718 75642
rect 65770 75590 65782 75642
rect 65834 75590 65846 75642
rect 65898 75590 65910 75642
rect 65962 75590 96374 75642
rect 96426 75590 96438 75642
rect 96490 75590 96502 75642
rect 96554 75590 96566 75642
rect 96618 75590 96630 75642
rect 96682 75590 108836 75642
rect 1104 75568 108836 75590
rect 86678 75488 86684 75540
rect 86736 75528 86742 75540
rect 86773 75531 86831 75537
rect 86773 75528 86785 75531
rect 86736 75500 86785 75528
rect 86736 75488 86742 75500
rect 86773 75497 86785 75500
rect 86819 75528 86831 75531
rect 88702 75528 88708 75540
rect 86819 75500 88708 75528
rect 86819 75497 86831 75500
rect 86773 75491 86831 75497
rect 88702 75488 88708 75500
rect 88760 75488 88766 75540
rect 89898 75488 89904 75540
rect 89956 75528 89962 75540
rect 90358 75528 90364 75540
rect 89956 75500 90364 75528
rect 89956 75488 89962 75500
rect 90358 75488 90364 75500
rect 90416 75528 90422 75540
rect 90637 75531 90695 75537
rect 90637 75528 90649 75531
rect 90416 75500 90649 75528
rect 90416 75488 90422 75500
rect 90637 75497 90649 75500
rect 90683 75497 90695 75531
rect 90637 75491 90695 75497
rect 86313 75463 86371 75469
rect 86313 75429 86325 75463
rect 86359 75460 86371 75463
rect 87414 75460 87420 75472
rect 86359 75432 87420 75460
rect 86359 75429 86371 75432
rect 86313 75423 86371 75429
rect 87414 75420 87420 75432
rect 87472 75420 87478 75472
rect 82725 75395 82783 75401
rect 82725 75392 82737 75395
rect 81820 75364 82737 75392
rect 1581 75327 1639 75333
rect 1581 75293 1593 75327
rect 1627 75324 1639 75327
rect 1627 75296 1808 75324
rect 1627 75293 1639 75296
rect 1581 75287 1639 75293
rect 842 75148 848 75200
rect 900 75188 906 75200
rect 1780 75197 1808 75296
rect 67358 75216 67364 75268
rect 67416 75256 67422 75268
rect 81820 75265 81848 75364
rect 82725 75361 82737 75364
rect 82771 75361 82783 75395
rect 82725 75355 82783 75361
rect 85577 75395 85635 75401
rect 85577 75361 85589 75395
rect 85623 75392 85635 75395
rect 86954 75392 86960 75404
rect 85623 75364 86960 75392
rect 85623 75361 85635 75364
rect 85577 75355 85635 75361
rect 86954 75352 86960 75364
rect 87012 75352 87018 75404
rect 88812 75364 93854 75392
rect 82170 75284 82176 75336
rect 82228 75284 82234 75336
rect 82449 75327 82507 75333
rect 82449 75293 82461 75327
rect 82495 75293 82507 75327
rect 82449 75287 82507 75293
rect 85485 75327 85543 75333
rect 85485 75293 85497 75327
rect 85531 75324 85543 75327
rect 86221 75327 86279 75333
rect 86221 75324 86233 75327
rect 85531 75296 86233 75324
rect 85531 75293 85543 75296
rect 85485 75287 85543 75293
rect 86221 75293 86233 75296
rect 86267 75293 86279 75327
rect 86221 75287 86279 75293
rect 81805 75259 81863 75265
rect 81805 75256 81817 75259
rect 67416 75228 81817 75256
rect 67416 75216 67422 75228
rect 81805 75225 81817 75228
rect 81851 75225 81863 75259
rect 82464 75256 82492 75287
rect 86236 75256 86264 75287
rect 86586 75284 86592 75336
rect 86644 75324 86650 75336
rect 88812 75324 88840 75364
rect 86644 75296 88840 75324
rect 86644 75284 86650 75296
rect 90450 75284 90456 75336
rect 90508 75324 90514 75336
rect 90508 75296 90864 75324
rect 90508 75284 90514 75296
rect 90836 75268 90864 75296
rect 87138 75256 87144 75268
rect 81805 75219 81863 75225
rect 82096 75228 82492 75256
rect 82832 75228 83214 75256
rect 86236 75228 87144 75256
rect 82096 75200 82124 75228
rect 1397 75191 1455 75197
rect 1397 75188 1409 75191
rect 900 75160 1409 75188
rect 900 75148 906 75160
rect 1397 75157 1409 75160
rect 1443 75157 1455 75191
rect 1397 75151 1455 75157
rect 1765 75191 1823 75197
rect 1765 75157 1777 75191
rect 1811 75188 1823 75191
rect 22002 75188 22008 75200
rect 1811 75160 22008 75188
rect 1811 75157 1823 75160
rect 1765 75151 1823 75157
rect 22002 75148 22008 75160
rect 22060 75148 22066 75200
rect 82078 75148 82084 75200
rect 82136 75148 82142 75200
rect 82265 75191 82323 75197
rect 82265 75157 82277 75191
rect 82311 75188 82323 75191
rect 82832 75188 82860 75228
rect 87138 75216 87144 75228
rect 87196 75216 87202 75268
rect 90818 75216 90824 75268
rect 90876 75216 90882 75268
rect 93826 75256 93854 75364
rect 108301 75327 108359 75333
rect 108301 75293 108313 75327
rect 108347 75293 108359 75327
rect 108301 75287 108359 75293
rect 108117 75259 108175 75265
rect 108117 75256 108129 75259
rect 93826 75228 108129 75256
rect 108117 75225 108129 75228
rect 108163 75256 108175 75259
rect 108316 75256 108344 75287
rect 108163 75228 108344 75256
rect 108163 75225 108175 75228
rect 108117 75219 108175 75225
rect 82311 75160 82860 75188
rect 84197 75191 84255 75197
rect 82311 75157 82323 75160
rect 82265 75151 82323 75157
rect 84197 75157 84209 75191
rect 84243 75188 84255 75191
rect 84378 75188 84384 75200
rect 84243 75160 84384 75188
rect 84243 75157 84255 75160
rect 84197 75151 84255 75157
rect 84378 75148 84384 75160
rect 84436 75148 84442 75200
rect 86957 75191 87015 75197
rect 86957 75157 86969 75191
rect 87003 75188 87015 75191
rect 87046 75188 87052 75200
rect 87003 75160 87052 75188
rect 87003 75157 87015 75160
rect 86957 75151 87015 75157
rect 87046 75148 87052 75160
rect 87104 75148 87110 75200
rect 90450 75148 90456 75200
rect 90508 75148 90514 75200
rect 90621 75191 90679 75197
rect 90621 75157 90633 75191
rect 90667 75188 90679 75191
rect 90726 75188 90732 75200
rect 90667 75160 90732 75188
rect 90667 75157 90679 75160
rect 90621 75151 90679 75157
rect 90726 75148 90732 75160
rect 90784 75148 90790 75200
rect 108482 75148 108488 75200
rect 108540 75148 108546 75200
rect 1104 75098 108836 75120
rect 1104 75046 4874 75098
rect 4926 75046 4938 75098
rect 4990 75046 5002 75098
rect 5054 75046 5066 75098
rect 5118 75046 5130 75098
rect 5182 75046 35594 75098
rect 35646 75046 35658 75098
rect 35710 75046 35722 75098
rect 35774 75046 35786 75098
rect 35838 75046 35850 75098
rect 35902 75046 66314 75098
rect 66366 75046 66378 75098
rect 66430 75046 66442 75098
rect 66494 75046 66506 75098
rect 66558 75046 66570 75098
rect 66622 75046 97034 75098
rect 97086 75046 97098 75098
rect 97150 75046 97162 75098
rect 97214 75046 97226 75098
rect 97278 75046 97290 75098
rect 97342 75046 108836 75098
rect 1104 75024 108836 75046
rect 82170 74944 82176 74996
rect 82228 74984 82234 74996
rect 82541 74987 82599 74993
rect 82541 74984 82553 74987
rect 82228 74956 82553 74984
rect 82228 74944 82234 74956
rect 82541 74953 82553 74956
rect 82587 74984 82599 74987
rect 82814 74984 82820 74996
rect 82587 74956 82820 74984
rect 82587 74953 82599 74956
rect 82541 74947 82599 74953
rect 82814 74944 82820 74956
rect 82872 74944 82878 74996
rect 84378 74944 84384 74996
rect 84436 74984 84442 74996
rect 102134 74984 102140 74996
rect 84436 74956 102140 74984
rect 84436 74944 84442 74956
rect 102134 74944 102140 74956
rect 102192 74944 102198 74996
rect 1104 74554 108836 74576
rect 1104 74502 4214 74554
rect 4266 74502 4278 74554
rect 4330 74502 4342 74554
rect 4394 74502 4406 74554
rect 4458 74502 4470 74554
rect 4522 74502 34934 74554
rect 34986 74502 34998 74554
rect 35050 74502 35062 74554
rect 35114 74502 35126 74554
rect 35178 74502 35190 74554
rect 35242 74502 65654 74554
rect 65706 74502 65718 74554
rect 65770 74502 65782 74554
rect 65834 74502 65846 74554
rect 65898 74502 65910 74554
rect 65962 74502 96374 74554
rect 96426 74502 96438 74554
rect 96490 74502 96502 74554
rect 96554 74502 96566 74554
rect 96618 74502 96630 74554
rect 96682 74502 108836 74554
rect 1104 74480 108836 74502
rect 842 74332 848 74384
rect 900 74372 906 74384
rect 1397 74375 1455 74381
rect 1397 74372 1409 74375
rect 900 74344 1409 74372
rect 900 74332 906 74344
rect 1397 74341 1409 74344
rect 1443 74341 1455 74375
rect 1397 74335 1455 74341
rect 1581 74239 1639 74245
rect 1581 74205 1593 74239
rect 1627 74236 1639 74239
rect 1765 74239 1823 74245
rect 1765 74236 1777 74239
rect 1627 74208 1777 74236
rect 1627 74205 1639 74208
rect 1581 74199 1639 74205
rect 1765 74205 1777 74208
rect 1811 74236 1823 74239
rect 22830 74236 22836 74248
rect 1811 74208 22836 74236
rect 1811 74205 1823 74208
rect 1765 74199 1823 74205
rect 22830 74196 22836 74208
rect 22888 74196 22894 74248
rect 85574 74196 85580 74248
rect 85632 74236 85638 74248
rect 108117 74239 108175 74245
rect 108117 74236 108129 74239
rect 85632 74208 108129 74236
rect 85632 74196 85638 74208
rect 108117 74205 108129 74208
rect 108163 74236 108175 74239
rect 108301 74239 108359 74245
rect 108301 74236 108313 74239
rect 108163 74208 108313 74236
rect 108163 74205 108175 74208
rect 108117 74199 108175 74205
rect 108301 74205 108313 74208
rect 108347 74205 108359 74239
rect 108301 74199 108359 74205
rect 108482 74060 108488 74112
rect 108540 74060 108546 74112
rect 1104 74010 108836 74032
rect 1104 73958 4874 74010
rect 4926 73958 4938 74010
rect 4990 73958 5002 74010
rect 5054 73958 5066 74010
rect 5118 73958 5130 74010
rect 5182 73958 35594 74010
rect 35646 73958 35658 74010
rect 35710 73958 35722 74010
rect 35774 73958 35786 74010
rect 35838 73958 35850 74010
rect 35902 73958 66314 74010
rect 66366 73958 66378 74010
rect 66430 73958 66442 74010
rect 66494 73958 66506 74010
rect 66558 73958 66570 74010
rect 66622 73958 97034 74010
rect 97086 73958 97098 74010
rect 97150 73958 97162 74010
rect 97214 73958 97226 74010
rect 97278 73958 97290 74010
rect 97342 73958 108836 74010
rect 1104 73936 108836 73958
rect 1581 73763 1639 73769
rect 1581 73729 1593 73763
rect 1627 73760 1639 73763
rect 1765 73763 1823 73769
rect 1765 73760 1777 73763
rect 1627 73732 1777 73760
rect 1627 73729 1639 73732
rect 1581 73723 1639 73729
rect 1765 73729 1777 73732
rect 1811 73760 1823 73763
rect 21358 73760 21364 73772
rect 1811 73732 21364 73760
rect 1811 73729 1823 73732
rect 1765 73723 1823 73729
rect 21358 73720 21364 73732
rect 21416 73720 21422 73772
rect 108301 73763 108359 73769
rect 108301 73760 108313 73763
rect 108132 73732 108313 73760
rect 842 73584 848 73636
rect 900 73624 906 73636
rect 1397 73627 1455 73633
rect 1397 73624 1409 73627
rect 900 73596 1409 73624
rect 900 73584 906 73596
rect 1397 73593 1409 73596
rect 1443 73593 1455 73627
rect 1397 73587 1455 73593
rect 102134 73516 102140 73568
rect 102192 73556 102198 73568
rect 108132 73565 108160 73732
rect 108301 73729 108313 73732
rect 108347 73729 108359 73763
rect 108301 73723 108359 73729
rect 108117 73559 108175 73565
rect 108117 73556 108129 73559
rect 102192 73528 108129 73556
rect 102192 73516 102198 73528
rect 108117 73525 108129 73528
rect 108163 73525 108175 73559
rect 108117 73519 108175 73525
rect 108482 73516 108488 73568
rect 108540 73516 108546 73568
rect 1104 73466 108836 73488
rect 1104 73414 4214 73466
rect 4266 73414 4278 73466
rect 4330 73414 4342 73466
rect 4394 73414 4406 73466
rect 4458 73414 4470 73466
rect 4522 73414 34934 73466
rect 34986 73414 34998 73466
rect 35050 73414 35062 73466
rect 35114 73414 35126 73466
rect 35178 73414 35190 73466
rect 35242 73414 65654 73466
rect 65706 73414 65718 73466
rect 65770 73414 65782 73466
rect 65834 73414 65846 73466
rect 65898 73414 65910 73466
rect 65962 73414 96374 73466
rect 96426 73414 96438 73466
rect 96490 73414 96502 73466
rect 96554 73414 96566 73466
rect 96618 73414 96630 73466
rect 96682 73414 108836 73466
rect 1104 73392 108836 73414
rect 1762 73312 1768 73364
rect 1820 73312 1826 73364
rect 108114 73312 108120 73364
rect 108172 73312 108178 73364
rect 88978 73244 88984 73296
rect 89036 73284 89042 73296
rect 90085 73287 90143 73293
rect 90085 73284 90097 73287
rect 89036 73256 90097 73284
rect 89036 73244 89042 73256
rect 90085 73253 90097 73256
rect 90131 73253 90143 73287
rect 90085 73247 90143 73253
rect 90266 73244 90272 73296
rect 90324 73284 90330 73296
rect 90634 73284 90640 73296
rect 90324 73256 90640 73284
rect 90324 73244 90330 73256
rect 90634 73244 90640 73256
rect 90692 73244 90698 73296
rect 1581 73151 1639 73157
rect 1581 73117 1593 73151
rect 1627 73148 1639 73151
rect 1762 73148 1768 73160
rect 1627 73120 1768 73148
rect 1627 73117 1639 73120
rect 1581 73111 1639 73117
rect 1762 73108 1768 73120
rect 1820 73108 1826 73160
rect 90085 73151 90143 73157
rect 90085 73117 90097 73151
rect 90131 73148 90143 73151
rect 90174 73148 90180 73160
rect 90131 73120 90180 73148
rect 90131 73117 90143 73120
rect 90085 73111 90143 73117
rect 90174 73108 90180 73120
rect 90232 73108 90238 73160
rect 90269 73151 90327 73157
rect 90269 73117 90281 73151
rect 90315 73148 90327 73151
rect 90450 73148 90456 73160
rect 90315 73120 90456 73148
rect 90315 73117 90327 73120
rect 90269 73111 90327 73117
rect 90450 73108 90456 73120
rect 90508 73148 90514 73160
rect 90634 73148 90640 73160
rect 90508 73120 90640 73148
rect 90508 73108 90514 73120
rect 90634 73108 90640 73120
rect 90692 73108 90698 73160
rect 108114 73108 108120 73160
rect 108172 73148 108178 73160
rect 108301 73151 108359 73157
rect 108301 73148 108313 73151
rect 108172 73120 108313 73148
rect 108172 73108 108178 73120
rect 108301 73117 108313 73120
rect 108347 73117 108359 73151
rect 108301 73111 108359 73117
rect 842 72972 848 73024
rect 900 73012 906 73024
rect 1397 73015 1455 73021
rect 1397 73012 1409 73015
rect 900 72984 1409 73012
rect 900 72972 906 72984
rect 1397 72981 1409 72984
rect 1443 72981 1455 73015
rect 1397 72975 1455 72981
rect 108482 72972 108488 73024
rect 108540 72972 108546 73024
rect 1104 72922 108836 72944
rect 1104 72870 4874 72922
rect 4926 72870 4938 72922
rect 4990 72870 5002 72922
rect 5054 72870 5066 72922
rect 5118 72870 5130 72922
rect 5182 72870 35594 72922
rect 35646 72870 35658 72922
rect 35710 72870 35722 72922
rect 35774 72870 35786 72922
rect 35838 72870 35850 72922
rect 35902 72870 66314 72922
rect 66366 72870 66378 72922
rect 66430 72870 66442 72922
rect 66494 72870 66506 72922
rect 66558 72870 66570 72922
rect 66622 72870 97034 72922
rect 97086 72870 97098 72922
rect 97150 72870 97162 72922
rect 97214 72870 97226 72922
rect 97278 72870 97290 72922
rect 97342 72870 108836 72922
rect 1104 72848 108836 72870
rect 26206 72780 44680 72808
rect 1118 72632 1124 72684
rect 1176 72672 1182 72684
rect 1489 72675 1547 72681
rect 1489 72672 1501 72675
rect 1176 72644 1501 72672
rect 1176 72632 1182 72644
rect 1489 72641 1501 72644
rect 1535 72672 1547 72675
rect 1949 72675 2007 72681
rect 1949 72672 1961 72675
rect 1535 72644 1961 72672
rect 1535 72641 1547 72644
rect 1489 72635 1547 72641
rect 1949 72641 1961 72644
rect 1995 72641 2007 72675
rect 1949 72635 2007 72641
rect 7282 72632 7288 72684
rect 7340 72672 7346 72684
rect 26206 72672 26234 72780
rect 26786 72700 26792 72752
rect 26844 72740 26850 72752
rect 44652 72749 44680 72780
rect 44637 72743 44695 72749
rect 26844 72712 44220 72740
rect 26844 72700 26850 72712
rect 44192 72684 44220 72712
rect 44637 72709 44649 72743
rect 44683 72740 44695 72743
rect 44683 72712 46612 72740
rect 44683 72709 44695 72712
rect 44637 72703 44695 72709
rect 7340 72644 26234 72672
rect 7340 72632 7346 72644
rect 44174 72632 44180 72684
rect 44232 72672 44238 72684
rect 46584 72681 46612 72712
rect 74074 72700 74080 72752
rect 74132 72700 74138 72752
rect 75089 72743 75147 72749
rect 75089 72709 75101 72743
rect 75135 72740 75147 72743
rect 77202 72740 77208 72752
rect 75135 72712 77208 72740
rect 75135 72709 75147 72712
rect 75089 72703 75147 72709
rect 77202 72700 77208 72712
rect 77260 72700 77266 72752
rect 46569 72675 46627 72681
rect 44232 72644 45554 72672
rect 44232 72632 44238 72644
rect 45526 72604 45554 72644
rect 46569 72641 46581 72675
rect 46615 72672 46627 72675
rect 46615 72644 55214 72672
rect 46615 72641 46627 72644
rect 46569 72635 46627 72641
rect 46385 72607 46443 72613
rect 46385 72604 46397 72607
rect 45526 72576 46397 72604
rect 46385 72573 46397 72576
rect 46431 72604 46443 72607
rect 46431 72576 46796 72604
rect 46431 72573 46443 72576
rect 46385 72567 46443 72573
rect 1673 72539 1731 72545
rect 1673 72505 1685 72539
rect 1719 72536 1731 72539
rect 1857 72539 1915 72545
rect 1857 72536 1869 72539
rect 1719 72508 1869 72536
rect 1719 72505 1731 72508
rect 1673 72499 1731 72505
rect 1857 72505 1869 72508
rect 1903 72536 1915 72539
rect 1903 72508 6914 72536
rect 1903 72505 1915 72508
rect 1857 72499 1915 72505
rect 6886 72468 6914 72508
rect 28166 72468 28172 72480
rect 6886 72440 28172 72468
rect 28166 72428 28172 72440
rect 28224 72428 28230 72480
rect 46768 72477 46796 72576
rect 55186 72536 55214 72644
rect 73617 72607 73675 72613
rect 73617 72573 73629 72607
rect 73663 72604 73675 72607
rect 75086 72604 75092 72616
rect 73663 72576 75092 72604
rect 73663 72573 73675 72576
rect 73617 72567 73675 72573
rect 75086 72564 75092 72576
rect 75144 72564 75150 72616
rect 75365 72607 75423 72613
rect 75365 72573 75377 72607
rect 75411 72604 75423 72607
rect 82078 72604 82084 72616
rect 75411 72576 82084 72604
rect 75411 72573 75423 72576
rect 75365 72567 75423 72573
rect 57790 72536 57796 72548
rect 55186 72508 57796 72536
rect 57790 72496 57796 72508
rect 57848 72496 57854 72548
rect 73448 72508 73752 72536
rect 73448 72477 73476 72508
rect 46753 72471 46811 72477
rect 46753 72437 46765 72471
rect 46799 72468 46811 72471
rect 73433 72471 73491 72477
rect 73433 72468 73445 72471
rect 46799 72440 73445 72468
rect 46799 72437 46811 72440
rect 46753 72431 46811 72437
rect 73433 72437 73445 72440
rect 73479 72437 73491 72471
rect 73724 72468 73752 72508
rect 75380 72468 75408 72567
rect 82078 72564 82084 72576
rect 82136 72564 82142 72616
rect 73724 72440 75408 72468
rect 73433 72431 73491 72437
rect 95142 72428 95148 72480
rect 95200 72468 95206 72480
rect 104342 72468 104348 72480
rect 95200 72440 104348 72468
rect 95200 72428 95206 72440
rect 104342 72428 104348 72440
rect 104400 72428 104406 72480
rect 1104 72378 108836 72400
rect 1104 72326 4214 72378
rect 4266 72326 4278 72378
rect 4330 72326 4342 72378
rect 4394 72326 4406 72378
rect 4458 72326 4470 72378
rect 4522 72326 34934 72378
rect 34986 72326 34998 72378
rect 35050 72326 35062 72378
rect 35114 72326 35126 72378
rect 35178 72326 35190 72378
rect 35242 72326 65654 72378
rect 65706 72326 65718 72378
rect 65770 72326 65782 72378
rect 65834 72326 65846 72378
rect 65898 72326 65910 72378
rect 65962 72326 96374 72378
rect 96426 72326 96438 72378
rect 96490 72326 96502 72378
rect 96554 72326 96566 72378
rect 96618 72326 96630 72378
rect 96682 72326 108836 72378
rect 1104 72304 108836 72326
rect 44174 72224 44180 72276
rect 44232 72264 44238 72276
rect 44637 72267 44695 72273
rect 44637 72264 44649 72267
rect 44232 72236 44649 72264
rect 44232 72224 44238 72236
rect 44637 72233 44649 72236
rect 44683 72233 44695 72267
rect 44637 72227 44695 72233
rect 74074 72224 74080 72276
rect 74132 72264 74138 72276
rect 74169 72267 74227 72273
rect 74169 72264 74181 72267
rect 74132 72236 74181 72264
rect 74132 72224 74138 72236
rect 74169 72233 74181 72236
rect 74215 72233 74227 72267
rect 94314 72264 94320 72276
rect 74169 72227 74227 72233
rect 84166 72236 94320 72264
rect 73982 72020 73988 72072
rect 74040 72060 74046 72072
rect 74077 72063 74135 72069
rect 74077 72060 74089 72063
rect 74040 72032 74089 72060
rect 74040 72020 74046 72032
rect 74077 72029 74089 72032
rect 74123 72060 74135 72063
rect 74350 72060 74356 72072
rect 74123 72032 74356 72060
rect 74123 72029 74135 72032
rect 74077 72023 74135 72029
rect 74350 72020 74356 72032
rect 74408 72020 74414 72072
rect 9582 71952 9588 72004
rect 9640 71992 9646 72004
rect 55861 71995 55919 72001
rect 55861 71992 55873 71995
rect 9640 71964 55873 71992
rect 9640 71952 9646 71964
rect 55861 71961 55873 71964
rect 55907 71992 55919 71995
rect 56045 71995 56103 72001
rect 56045 71992 56057 71995
rect 55907 71964 56057 71992
rect 55907 71961 55919 71964
rect 55861 71955 55919 71961
rect 56045 71961 56057 71964
rect 56091 71961 56103 71995
rect 56045 71955 56103 71961
rect 57790 71952 57796 72004
rect 57848 71952 57854 72004
rect 64846 71964 74534 71992
rect 57808 71924 57836 71952
rect 57977 71927 58035 71933
rect 57977 71924 57989 71927
rect 57808 71896 57989 71924
rect 57977 71893 57989 71896
rect 58023 71924 58035 71927
rect 64846 71924 64874 71964
rect 58023 71896 64874 71924
rect 58023 71893 58035 71896
rect 57977 71887 58035 71893
rect 74350 71884 74356 71936
rect 74408 71884 74414 71936
rect 74506 71924 74534 71964
rect 84166 71924 84194 72236
rect 94314 72224 94320 72236
rect 94372 72264 94378 72276
rect 95142 72264 95148 72276
rect 94372 72236 95148 72264
rect 94372 72224 94378 72236
rect 95142 72224 95148 72236
rect 95200 72224 95206 72276
rect 90729 72063 90787 72069
rect 90729 72029 90741 72063
rect 90775 72060 90787 72063
rect 90818 72060 90824 72072
rect 90775 72032 90824 72060
rect 90775 72029 90787 72032
rect 90729 72023 90787 72029
rect 90818 72020 90824 72032
rect 90876 72060 90882 72072
rect 91557 72063 91615 72069
rect 91557 72060 91569 72063
rect 90876 72032 91569 72060
rect 90876 72020 90882 72032
rect 91557 72029 91569 72032
rect 91603 72029 91615 72063
rect 91557 72023 91615 72029
rect 90358 71952 90364 72004
rect 90416 71992 90422 72004
rect 91741 71995 91799 72001
rect 91741 71992 91753 71995
rect 90416 71964 91753 71992
rect 90416 71952 90422 71964
rect 91741 71961 91753 71964
rect 91787 71961 91799 71995
rect 91741 71955 91799 71961
rect 91925 71995 91983 72001
rect 91925 71961 91937 71995
rect 91971 71992 91983 71995
rect 92382 71992 92388 72004
rect 91971 71964 92388 71992
rect 91971 71961 91983 71964
rect 91925 71955 91983 71961
rect 92382 71952 92388 71964
rect 92440 71992 92446 72004
rect 92477 71995 92535 72001
rect 92477 71992 92489 71995
rect 92440 71964 92489 71992
rect 92440 71952 92446 71964
rect 92477 71961 92489 71964
rect 92523 71961 92535 71995
rect 92477 71955 92535 71961
rect 92661 71995 92719 72001
rect 92661 71961 92673 71995
rect 92707 71992 92719 71995
rect 92845 71995 92903 72001
rect 92845 71992 92857 71995
rect 92707 71964 92857 71992
rect 92707 71961 92719 71964
rect 92661 71955 92719 71961
rect 92845 71961 92857 71964
rect 92891 71992 92903 71995
rect 102870 71992 102876 72004
rect 92891 71964 102876 71992
rect 92891 71961 92903 71964
rect 92845 71955 92903 71961
rect 102870 71952 102876 71964
rect 102928 71952 102934 72004
rect 74506 71896 84194 71924
rect 87690 71884 87696 71936
rect 87748 71924 87754 71936
rect 90545 71927 90603 71933
rect 90545 71924 90557 71927
rect 87748 71896 90557 71924
rect 87748 71884 87754 71896
rect 90545 71893 90557 71896
rect 90591 71893 90603 71927
rect 90545 71887 90603 71893
rect 91830 71884 91836 71936
rect 91888 71884 91894 71936
rect 92106 71884 92112 71936
rect 92164 71884 92170 71936
rect 1104 71834 108836 71856
rect 1104 71782 4874 71834
rect 4926 71782 4938 71834
rect 4990 71782 5002 71834
rect 5054 71782 5066 71834
rect 5118 71782 5130 71834
rect 5182 71782 35594 71834
rect 35646 71782 35658 71834
rect 35710 71782 35722 71834
rect 35774 71782 35786 71834
rect 35838 71782 35850 71834
rect 35902 71782 66314 71834
rect 66366 71782 66378 71834
rect 66430 71782 66442 71834
rect 66494 71782 66506 71834
rect 66558 71782 66570 71834
rect 66622 71782 97034 71834
rect 97086 71782 97098 71834
rect 97150 71782 97162 71834
rect 97214 71782 97226 71834
rect 97278 71782 97290 71834
rect 97342 71782 108836 71834
rect 1104 71760 108836 71782
rect 90726 71680 90732 71732
rect 90784 71680 90790 71732
rect 90913 71587 90971 71593
rect 90913 71553 90925 71587
rect 90959 71584 90971 71587
rect 91094 71584 91100 71596
rect 90959 71556 91100 71584
rect 90959 71553 90971 71556
rect 90913 71547 90971 71553
rect 91094 71544 91100 71556
rect 91152 71584 91158 71596
rect 91830 71584 91836 71596
rect 91152 71556 91836 71584
rect 91152 71544 91158 71556
rect 91830 71544 91836 71556
rect 91888 71544 91894 71596
rect 92017 71383 92075 71389
rect 92017 71349 92029 71383
rect 92063 71380 92075 71383
rect 92293 71383 92351 71389
rect 92293 71380 92305 71383
rect 92063 71352 92305 71380
rect 92063 71349 92075 71352
rect 92017 71343 92075 71349
rect 92293 71349 92305 71352
rect 92339 71380 92351 71383
rect 102226 71380 102232 71392
rect 92339 71352 102232 71380
rect 92339 71349 92351 71352
rect 92293 71343 92351 71349
rect 102226 71340 102232 71352
rect 102284 71340 102290 71392
rect 1104 71290 108836 71312
rect 1104 71238 4214 71290
rect 4266 71238 4278 71290
rect 4330 71238 4342 71290
rect 4394 71238 4406 71290
rect 4458 71238 4470 71290
rect 4522 71238 34934 71290
rect 34986 71238 34998 71290
rect 35050 71238 35062 71290
rect 35114 71238 35126 71290
rect 35178 71238 35190 71290
rect 35242 71238 65654 71290
rect 65706 71238 65718 71290
rect 65770 71238 65782 71290
rect 65834 71238 65846 71290
rect 65898 71238 65910 71290
rect 65962 71238 96374 71290
rect 96426 71238 96438 71290
rect 96490 71238 96502 71290
rect 96554 71238 96566 71290
rect 96618 71238 96630 71290
rect 96682 71238 108836 71290
rect 1104 71216 108836 71238
rect 90453 71179 90511 71185
rect 90453 71145 90465 71179
rect 90499 71176 90511 71179
rect 91094 71176 91100 71188
rect 90499 71148 91100 71176
rect 90499 71145 90511 71148
rect 90453 71139 90511 71145
rect 91094 71136 91100 71148
rect 91152 71136 91158 71188
rect 74626 71000 74632 71052
rect 74684 71040 74690 71052
rect 77757 71043 77815 71049
rect 77757 71040 77769 71043
rect 74684 71012 77769 71040
rect 74684 71000 74690 71012
rect 77757 71009 77769 71012
rect 77803 71040 77815 71043
rect 78030 71040 78036 71052
rect 77803 71012 78036 71040
rect 77803 71009 77815 71012
rect 77757 71003 77815 71009
rect 78030 71000 78036 71012
rect 78088 71040 78094 71052
rect 78125 71043 78183 71049
rect 78125 71040 78137 71043
rect 78088 71012 78137 71040
rect 78088 71000 78094 71012
rect 78125 71009 78137 71012
rect 78171 71009 78183 71043
rect 78125 71003 78183 71009
rect 88702 71000 88708 71052
rect 88760 71040 88766 71052
rect 90545 71043 90603 71049
rect 90545 71040 90557 71043
rect 88760 71012 90557 71040
rect 88760 71000 88766 71012
rect 90545 71009 90557 71012
rect 90591 71009 90603 71043
rect 90545 71003 90603 71009
rect 75086 70932 75092 70984
rect 75144 70972 75150 70984
rect 77573 70975 77631 70981
rect 77573 70972 77585 70975
rect 75144 70944 77585 70972
rect 75144 70932 75150 70944
rect 77573 70941 77585 70944
rect 77619 70941 77631 70975
rect 77573 70935 77631 70941
rect 87138 70932 87144 70984
rect 87196 70972 87202 70984
rect 87874 70972 87880 70984
rect 87196 70944 87880 70972
rect 87196 70932 87202 70944
rect 87874 70932 87880 70944
rect 87932 70932 87938 70984
rect 88978 70864 88984 70916
rect 89036 70864 89042 70916
rect 89088 70876 89470 70904
rect 87969 70839 88027 70845
rect 87969 70805 87981 70839
rect 88015 70836 88027 70839
rect 89088 70836 89116 70876
rect 88015 70808 89116 70836
rect 88015 70805 88027 70808
rect 87969 70799 88027 70805
rect 1104 70746 108836 70768
rect 1104 70694 4874 70746
rect 4926 70694 4938 70746
rect 4990 70694 5002 70746
rect 5054 70694 5066 70746
rect 5118 70694 5130 70746
rect 5182 70694 35594 70746
rect 35646 70694 35658 70746
rect 35710 70694 35722 70746
rect 35774 70694 35786 70746
rect 35838 70694 35850 70746
rect 35902 70694 66314 70746
rect 66366 70694 66378 70746
rect 66430 70694 66442 70746
rect 66494 70694 66506 70746
rect 66558 70694 66570 70746
rect 66622 70694 97034 70746
rect 97086 70694 97098 70746
rect 97150 70694 97162 70746
rect 97214 70694 97226 70746
rect 97278 70694 97290 70746
rect 97342 70694 108836 70746
rect 1104 70672 108836 70694
rect 78030 70592 78036 70644
rect 78088 70592 78094 70644
rect 77757 70499 77815 70505
rect 77757 70465 77769 70499
rect 77803 70496 77815 70499
rect 78048 70496 78076 70592
rect 77803 70468 78076 70496
rect 77803 70465 77815 70468
rect 77757 70459 77815 70465
rect 77202 70388 77208 70440
rect 77260 70428 77266 70440
rect 77389 70431 77447 70437
rect 77389 70428 77401 70431
rect 77260 70400 77401 70428
rect 77260 70388 77266 70400
rect 77389 70397 77401 70400
rect 77435 70397 77447 70431
rect 77389 70391 77447 70397
rect 77849 70431 77907 70437
rect 77849 70397 77861 70431
rect 77895 70428 77907 70431
rect 85666 70428 85672 70440
rect 77895 70400 85672 70428
rect 77895 70397 77907 70400
rect 77849 70391 77907 70397
rect 85666 70388 85672 70400
rect 85724 70388 85730 70440
rect 1104 70202 108836 70224
rect 1104 70150 4214 70202
rect 4266 70150 4278 70202
rect 4330 70150 4342 70202
rect 4394 70150 4406 70202
rect 4458 70150 4470 70202
rect 4522 70150 34934 70202
rect 34986 70150 34998 70202
rect 35050 70150 35062 70202
rect 35114 70150 35126 70202
rect 35178 70150 35190 70202
rect 35242 70150 65654 70202
rect 65706 70150 65718 70202
rect 65770 70150 65782 70202
rect 65834 70150 65846 70202
rect 65898 70150 65910 70202
rect 65962 70150 96374 70202
rect 96426 70150 96438 70202
rect 96490 70150 96502 70202
rect 96554 70150 96566 70202
rect 96618 70150 96630 70202
rect 96682 70150 108836 70202
rect 1104 70128 108836 70150
rect 1104 69658 108836 69680
rect 1104 69606 4874 69658
rect 4926 69606 4938 69658
rect 4990 69606 5002 69658
rect 5054 69606 5066 69658
rect 5118 69606 5130 69658
rect 5182 69606 35594 69658
rect 35646 69606 35658 69658
rect 35710 69606 35722 69658
rect 35774 69606 35786 69658
rect 35838 69606 35850 69658
rect 35902 69606 66314 69658
rect 66366 69606 66378 69658
rect 66430 69606 66442 69658
rect 66494 69606 66506 69658
rect 66558 69606 66570 69658
rect 66622 69606 97034 69658
rect 97086 69606 97098 69658
rect 97150 69606 97162 69658
rect 97214 69606 97226 69658
rect 97278 69606 97290 69658
rect 97342 69606 108836 69658
rect 1104 69584 108836 69606
rect 88978 69164 88984 69216
rect 89036 69204 89042 69216
rect 89073 69207 89131 69213
rect 89073 69204 89085 69207
rect 89036 69176 89085 69204
rect 89036 69164 89042 69176
rect 89073 69173 89085 69176
rect 89119 69204 89131 69207
rect 89162 69204 89168 69216
rect 89119 69176 89168 69204
rect 89119 69173 89131 69176
rect 89073 69167 89131 69173
rect 89162 69164 89168 69176
rect 89220 69164 89226 69216
rect 1104 69114 108836 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 34934 69114
rect 34986 69062 34998 69114
rect 35050 69062 35062 69114
rect 35114 69062 35126 69114
rect 35178 69062 35190 69114
rect 35242 69062 65654 69114
rect 65706 69062 65718 69114
rect 65770 69062 65782 69114
rect 65834 69062 65846 69114
rect 65898 69062 65910 69114
rect 65962 69062 96374 69114
rect 96426 69062 96438 69114
rect 96490 69062 96502 69114
rect 96554 69062 96566 69114
rect 96618 69062 96630 69114
rect 96682 69062 108836 69114
rect 1104 69040 108836 69062
rect 88978 68892 88984 68944
rect 89036 68932 89042 68944
rect 89806 68932 89812 68944
rect 89036 68904 89812 68932
rect 89036 68892 89042 68904
rect 89806 68892 89812 68904
rect 89864 68932 89870 68944
rect 90729 68935 90787 68941
rect 90729 68932 90741 68935
rect 89864 68904 90741 68932
rect 89864 68892 89870 68904
rect 90729 68901 90741 68904
rect 90775 68901 90787 68935
rect 90729 68895 90787 68901
rect 89257 68867 89315 68873
rect 89257 68864 89269 68867
rect 80026 68836 89269 68864
rect 74350 68688 74356 68740
rect 74408 68728 74414 68740
rect 80026 68728 80054 68836
rect 89257 68833 89269 68836
rect 89303 68864 89315 68867
rect 89303 68836 89944 68864
rect 89303 68833 89315 68836
rect 89257 68827 89315 68833
rect 88978 68756 88984 68808
rect 89036 68756 89042 68808
rect 89533 68799 89591 68805
rect 89533 68765 89545 68799
rect 89579 68765 89591 68799
rect 89533 68759 89591 68765
rect 74408 68700 80054 68728
rect 74408 68688 74414 68700
rect 87874 68688 87880 68740
rect 87932 68728 87938 68740
rect 88242 68728 88248 68740
rect 87932 68700 88248 68728
rect 87932 68688 87938 68700
rect 88242 68688 88248 68700
rect 88300 68728 88306 68740
rect 88705 68731 88763 68737
rect 88705 68728 88717 68731
rect 88300 68700 88717 68728
rect 88300 68688 88306 68700
rect 88705 68697 88717 68700
rect 88751 68697 88763 68731
rect 88705 68691 88763 68697
rect 89548 68660 89576 68759
rect 89806 68756 89812 68808
rect 89864 68756 89870 68808
rect 89916 68796 89944 68836
rect 90085 68799 90143 68805
rect 90085 68796 90097 68799
rect 89916 68768 90097 68796
rect 90085 68765 90097 68768
rect 90131 68796 90143 68799
rect 90177 68799 90235 68805
rect 90177 68796 90189 68799
rect 90131 68768 90189 68796
rect 90131 68765 90143 68768
rect 90085 68759 90143 68765
rect 90177 68765 90189 68768
rect 90223 68796 90235 68799
rect 90545 68799 90603 68805
rect 90545 68796 90557 68799
rect 90223 68768 90557 68796
rect 90223 68765 90235 68768
rect 90177 68759 90235 68765
rect 90545 68765 90557 68768
rect 90591 68765 90603 68799
rect 90545 68759 90603 68765
rect 90634 68756 90640 68808
rect 90692 68796 90698 68808
rect 92201 68799 92259 68805
rect 92201 68796 92213 68799
rect 90692 68768 92213 68796
rect 90692 68756 90698 68768
rect 92201 68765 92213 68768
rect 92247 68765 92259 68799
rect 92201 68759 92259 68765
rect 92382 68756 92388 68808
rect 92440 68756 92446 68808
rect 90744 68700 99374 68728
rect 90453 68663 90511 68669
rect 90453 68660 90465 68663
rect 89548 68632 90465 68660
rect 90453 68629 90465 68632
rect 90499 68660 90511 68663
rect 90744 68660 90772 68700
rect 90499 68632 90772 68660
rect 90499 68629 90511 68632
rect 90453 68623 90511 68629
rect 91094 68620 91100 68672
rect 91152 68660 91158 68672
rect 92293 68663 92351 68669
rect 92293 68660 92305 68663
rect 91152 68632 92305 68660
rect 91152 68620 91158 68632
rect 92293 68629 92305 68632
rect 92339 68629 92351 68663
rect 99346 68660 99374 68700
rect 107930 68660 107936 68672
rect 99346 68632 107936 68660
rect 92293 68623 92351 68629
rect 107930 68620 107936 68632
rect 107988 68620 107994 68672
rect 1104 68570 108836 68592
rect 1104 68518 4874 68570
rect 4926 68518 4938 68570
rect 4990 68518 5002 68570
rect 5054 68518 5066 68570
rect 5118 68518 5130 68570
rect 5182 68518 35594 68570
rect 35646 68518 35658 68570
rect 35710 68518 35722 68570
rect 35774 68518 35786 68570
rect 35838 68518 35850 68570
rect 35902 68518 66314 68570
rect 66366 68518 66378 68570
rect 66430 68518 66442 68570
rect 66494 68518 66506 68570
rect 66558 68518 66570 68570
rect 66622 68518 97034 68570
rect 97086 68518 97098 68570
rect 97150 68518 97162 68570
rect 97214 68518 97226 68570
rect 97278 68518 97290 68570
rect 97342 68518 108836 68570
rect 1104 68496 108836 68518
rect 85482 68280 85488 68332
rect 85540 68320 85546 68332
rect 86589 68323 86647 68329
rect 86589 68320 86601 68323
rect 85540 68292 86601 68320
rect 85540 68280 85546 68292
rect 86589 68289 86601 68292
rect 86635 68320 86647 68323
rect 88242 68320 88248 68332
rect 86635 68292 88248 68320
rect 86635 68289 86647 68292
rect 86589 68283 86647 68289
rect 88242 68280 88248 68292
rect 88300 68320 88306 68332
rect 88981 68323 89039 68329
rect 88981 68320 88993 68323
rect 88300 68292 88993 68320
rect 88300 68280 88306 68292
rect 88981 68289 88993 68292
rect 89027 68289 89039 68323
rect 88981 68283 89039 68289
rect 86681 68119 86739 68125
rect 86681 68085 86693 68119
rect 86727 68116 86739 68119
rect 86954 68116 86960 68128
rect 86727 68088 86960 68116
rect 86727 68085 86739 68088
rect 86681 68079 86739 68085
rect 86954 68076 86960 68088
rect 87012 68076 87018 68128
rect 89073 68119 89131 68125
rect 89073 68085 89085 68119
rect 89119 68116 89131 68119
rect 90726 68116 90732 68128
rect 89119 68088 90732 68116
rect 89119 68085 89131 68088
rect 89073 68079 89131 68085
rect 90726 68076 90732 68088
rect 90784 68076 90790 68128
rect 1104 68026 108836 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 34934 68026
rect 34986 67974 34998 68026
rect 35050 67974 35062 68026
rect 35114 67974 35126 68026
rect 35178 67974 35190 68026
rect 35242 67974 65654 68026
rect 65706 67974 65718 68026
rect 65770 67974 65782 68026
rect 65834 67974 65846 68026
rect 65898 67974 65910 68026
rect 65962 67974 96374 68026
rect 96426 67974 96438 68026
rect 96490 67974 96502 68026
rect 96554 67974 96566 68026
rect 96618 67974 96630 68026
rect 96682 67974 108836 68026
rect 1104 67952 108836 67974
rect 90542 67872 90548 67924
rect 90600 67872 90606 67924
rect 107930 67872 107936 67924
rect 107988 67912 107994 67924
rect 108301 67915 108359 67921
rect 108301 67912 108313 67915
rect 107988 67884 108313 67912
rect 107988 67872 107994 67884
rect 108301 67881 108313 67884
rect 108347 67881 108359 67915
rect 108301 67875 108359 67881
rect 88797 67847 88855 67853
rect 88797 67813 88809 67847
rect 88843 67844 88855 67847
rect 92569 67847 92627 67853
rect 88843 67816 89714 67844
rect 88843 67813 88855 67816
rect 88797 67807 88855 67813
rect 89686 67776 89714 67816
rect 92569 67813 92581 67847
rect 92615 67844 92627 67847
rect 92845 67847 92903 67853
rect 92845 67844 92857 67847
rect 92615 67816 92857 67844
rect 92615 67813 92627 67816
rect 92569 67807 92627 67813
rect 92845 67813 92857 67816
rect 92891 67844 92903 67847
rect 101950 67844 101956 67856
rect 92891 67816 101956 67844
rect 92891 67813 92903 67816
rect 92845 67807 92903 67813
rect 101950 67804 101956 67816
rect 102008 67804 102014 67856
rect 91554 67776 91560 67788
rect 89686 67748 90404 67776
rect 84378 67668 84384 67720
rect 84436 67708 84442 67720
rect 85482 67708 85488 67720
rect 84436 67680 85488 67708
rect 84436 67668 84442 67680
rect 85482 67668 85488 67680
rect 85540 67708 85546 67720
rect 86221 67711 86279 67717
rect 86221 67708 86233 67711
rect 85540 67680 86233 67708
rect 85540 67668 85546 67680
rect 86221 67677 86233 67680
rect 86267 67677 86279 67711
rect 86221 67671 86279 67677
rect 88426 67668 88432 67720
rect 88484 67708 88490 67720
rect 88613 67711 88671 67717
rect 88613 67708 88625 67711
rect 88484 67680 88625 67708
rect 88484 67668 88490 67680
rect 88613 67677 88625 67680
rect 88659 67677 88671 67711
rect 89717 67711 89775 67717
rect 89717 67708 89729 67711
rect 88613 67671 88671 67677
rect 89456 67680 89729 67708
rect 86313 67643 86371 67649
rect 86313 67609 86325 67643
rect 86359 67640 86371 67643
rect 87046 67640 87052 67652
rect 86359 67612 87052 67640
rect 86359 67609 86371 67612
rect 86313 67603 86371 67609
rect 87046 67600 87052 67612
rect 87104 67600 87110 67652
rect 89346 67600 89352 67652
rect 89404 67640 89410 67652
rect 89456 67649 89484 67680
rect 89717 67677 89729 67680
rect 89763 67677 89775 67711
rect 89717 67671 89775 67677
rect 89806 67668 89812 67720
rect 89864 67708 89870 67720
rect 90376 67717 90404 67748
rect 90928 67748 91560 67776
rect 90177 67711 90235 67717
rect 90177 67708 90189 67711
rect 89864 67680 90189 67708
rect 89864 67668 89870 67680
rect 90177 67677 90189 67680
rect 90223 67677 90235 67711
rect 90177 67671 90235 67677
rect 90361 67711 90419 67717
rect 90361 67677 90373 67711
rect 90407 67708 90419 67711
rect 90542 67708 90548 67720
rect 90407 67680 90548 67708
rect 90407 67677 90419 67680
rect 90361 67671 90419 67677
rect 90542 67668 90548 67680
rect 90600 67668 90606 67720
rect 90928 67717 90956 67748
rect 91554 67736 91560 67748
rect 91612 67776 91618 67788
rect 92106 67776 92112 67788
rect 91612 67748 92112 67776
rect 91612 67736 91618 67748
rect 92106 67736 92112 67748
rect 92164 67736 92170 67788
rect 90913 67711 90971 67717
rect 90913 67677 90925 67711
rect 90959 67677 90971 67711
rect 90913 67671 90971 67677
rect 91094 67668 91100 67720
rect 91152 67668 91158 67720
rect 92382 67668 92388 67720
rect 92440 67668 92446 67720
rect 108209 67711 108267 67717
rect 108209 67677 108221 67711
rect 108255 67708 108267 67711
rect 108482 67708 108488 67720
rect 108255 67680 108488 67708
rect 108255 67677 108267 67680
rect 108209 67671 108267 67677
rect 108482 67668 108488 67680
rect 108540 67668 108546 67720
rect 89441 67643 89499 67649
rect 89441 67640 89453 67643
rect 89404 67612 89453 67640
rect 89404 67600 89410 67612
rect 89441 67609 89453 67612
rect 89487 67609 89499 67643
rect 89441 67603 89499 67609
rect 89625 67643 89683 67649
rect 89625 67609 89637 67643
rect 89671 67640 89683 67643
rect 90085 67643 90143 67649
rect 90085 67640 90097 67643
rect 89671 67612 90097 67640
rect 89671 67609 89683 67612
rect 89625 67603 89683 67609
rect 90085 67609 90097 67612
rect 90131 67640 90143 67643
rect 102962 67640 102968 67652
rect 90131 67612 102968 67640
rect 90131 67609 90143 67612
rect 90085 67603 90143 67609
rect 102962 67600 102968 67612
rect 103020 67600 103026 67652
rect 89901 67575 89959 67581
rect 89901 67541 89913 67575
rect 89947 67572 89959 67575
rect 89990 67572 89996 67584
rect 89947 67544 89996 67572
rect 89947 67541 89959 67544
rect 89901 67535 89959 67541
rect 89990 67532 89996 67544
rect 90048 67532 90054 67584
rect 91005 67575 91063 67581
rect 91005 67541 91017 67575
rect 91051 67572 91063 67575
rect 91094 67572 91100 67584
rect 91051 67544 91100 67572
rect 91051 67541 91063 67544
rect 91005 67535 91063 67541
rect 91094 67532 91100 67544
rect 91152 67532 91158 67584
rect 1104 67482 108836 67504
rect 1104 67430 4874 67482
rect 4926 67430 4938 67482
rect 4990 67430 5002 67482
rect 5054 67430 5066 67482
rect 5118 67430 5130 67482
rect 5182 67430 35594 67482
rect 35646 67430 35658 67482
rect 35710 67430 35722 67482
rect 35774 67430 35786 67482
rect 35838 67430 35850 67482
rect 35902 67430 66314 67482
rect 66366 67430 66378 67482
rect 66430 67430 66442 67482
rect 66494 67430 66506 67482
rect 66558 67430 66570 67482
rect 66622 67430 97034 67482
rect 97086 67430 97098 67482
rect 97150 67430 97162 67482
rect 97214 67430 97226 67482
rect 97278 67430 97290 67482
rect 97342 67430 108836 67482
rect 1104 67408 108836 67430
rect 88613 67371 88671 67377
rect 88613 67337 88625 67371
rect 88659 67368 88671 67371
rect 88702 67368 88708 67380
rect 88659 67340 88708 67368
rect 88659 67337 88671 67340
rect 88613 67331 88671 67337
rect 88628 67300 88656 67331
rect 88702 67328 88708 67340
rect 88760 67368 88766 67380
rect 88797 67371 88855 67377
rect 88797 67368 88809 67371
rect 88760 67340 88809 67368
rect 88760 67328 88766 67340
rect 88797 67337 88809 67340
rect 88843 67337 88855 67371
rect 88797 67331 88855 67337
rect 89714 67328 89720 67380
rect 89772 67368 89778 67380
rect 90174 67368 90180 67380
rect 89772 67340 90180 67368
rect 89772 67328 89778 67340
rect 90174 67328 90180 67340
rect 90232 67328 90238 67380
rect 91094 67368 91100 67380
rect 90284 67340 91100 67368
rect 89162 67300 89168 67312
rect 88628 67272 89168 67300
rect 83921 67235 83979 67241
rect 83921 67201 83933 67235
rect 83967 67232 83979 67235
rect 84378 67232 84384 67244
rect 83967 67204 84384 67232
rect 83967 67201 83979 67204
rect 83921 67195 83979 67201
rect 84378 67192 84384 67204
rect 84436 67192 84442 67244
rect 87046 67192 87052 67244
rect 87104 67192 87110 67244
rect 88429 67235 88487 67241
rect 88429 67201 88441 67235
rect 88475 67232 88487 67235
rect 88628 67232 88656 67272
rect 89162 67260 89168 67272
rect 89220 67300 89226 67312
rect 90284 67309 90312 67340
rect 91094 67328 91100 67340
rect 91152 67328 91158 67380
rect 91741 67371 91799 67377
rect 91741 67337 91753 67371
rect 91787 67368 91799 67371
rect 92382 67368 92388 67380
rect 91787 67340 92388 67368
rect 91787 67337 91799 67340
rect 91741 67331 91799 67337
rect 92382 67328 92388 67340
rect 92440 67328 92446 67380
rect 90269 67303 90327 67309
rect 89220 67272 90036 67300
rect 89220 67260 89226 67272
rect 88475 67204 88656 67232
rect 88475 67201 88487 67204
rect 88429 67195 88487 67201
rect 88702 67192 88708 67244
rect 88760 67232 88766 67244
rect 89346 67232 89352 67244
rect 88760 67204 89352 67232
rect 88760 67192 88766 67204
rect 89346 67192 89352 67204
rect 89404 67192 89410 67244
rect 89530 67192 89536 67244
rect 89588 67232 89594 67244
rect 90008 67241 90036 67272
rect 90269 67269 90281 67303
rect 90315 67269 90327 67303
rect 90269 67263 90327 67269
rect 90726 67260 90732 67312
rect 90784 67260 90790 67312
rect 89625 67235 89683 67241
rect 89625 67232 89637 67235
rect 89588 67204 89637 67232
rect 89588 67192 89594 67204
rect 89625 67201 89637 67204
rect 89671 67201 89683 67235
rect 89625 67195 89683 67201
rect 89993 67235 90051 67241
rect 89993 67201 90005 67235
rect 90039 67201 90051 67235
rect 89993 67195 90051 67201
rect 88153 67167 88211 67173
rect 88153 67133 88165 67167
rect 88199 67164 88211 67167
rect 89254 67164 89260 67176
rect 88199 67136 89260 67164
rect 88199 67133 88211 67136
rect 88153 67127 88211 67133
rect 89254 67124 89260 67136
rect 89312 67124 89318 67176
rect 89441 67167 89499 67173
rect 89441 67133 89453 67167
rect 89487 67164 89499 67167
rect 89487 67136 89852 67164
rect 89487 67133 89499 67136
rect 89441 67127 89499 67133
rect 89824 67096 89852 67136
rect 89898 67096 89904 67108
rect 89824 67068 89904 67096
rect 89898 67056 89904 67068
rect 89956 67056 89962 67108
rect 83829 67031 83887 67037
rect 83829 66997 83841 67031
rect 83875 67028 83887 67031
rect 84378 67028 84384 67040
rect 83875 67000 84384 67028
rect 83875 66997 83887 67000
rect 83829 66991 83887 66997
rect 84378 66988 84384 67000
rect 84436 66988 84442 67040
rect 84473 67031 84531 67037
rect 84473 66997 84485 67031
rect 84519 67028 84531 67031
rect 85574 67028 85580 67040
rect 84519 67000 85580 67028
rect 84519 66997 84531 67000
rect 84473 66991 84531 66997
rect 85574 66988 85580 67000
rect 85632 66988 85638 67040
rect 86681 67031 86739 67037
rect 86681 66997 86693 67031
rect 86727 67028 86739 67031
rect 88426 67028 88432 67040
rect 86727 67000 88432 67028
rect 86727 66997 86739 67000
rect 86681 66991 86739 66997
rect 88426 66988 88432 67000
rect 88484 66988 88490 67040
rect 88886 66988 88892 67040
rect 88944 67028 88950 67040
rect 88981 67031 89039 67037
rect 88981 67028 88993 67031
rect 88944 67000 88993 67028
rect 88944 66988 88950 67000
rect 88981 66997 88993 67000
rect 89027 66997 89039 67031
rect 88981 66991 89039 66997
rect 89806 66988 89812 67040
rect 89864 66988 89870 67040
rect 90008 67028 90036 67195
rect 90266 67124 90272 67176
rect 90324 67164 90330 67176
rect 91554 67164 91560 67176
rect 90324 67136 91560 67164
rect 90324 67124 90330 67136
rect 91554 67124 91560 67136
rect 91612 67124 91618 67176
rect 91925 67031 91983 67037
rect 91925 67028 91937 67031
rect 90008 67000 91937 67028
rect 91925 66997 91937 67000
rect 91971 67028 91983 67031
rect 95878 67028 95884 67040
rect 91971 67000 95884 67028
rect 91971 66997 91983 67000
rect 91925 66991 91983 66997
rect 95878 66988 95884 67000
rect 95936 66988 95942 67040
rect 1104 66938 108836 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 96374 66938
rect 96426 66886 96438 66938
rect 96490 66886 96502 66938
rect 96554 66886 96566 66938
rect 96618 66886 96630 66938
rect 96682 66886 108836 66938
rect 1104 66864 108836 66886
rect 82078 66784 82084 66836
rect 82136 66824 82142 66836
rect 83829 66827 83887 66833
rect 83829 66824 83841 66827
rect 82136 66796 83841 66824
rect 82136 66784 82142 66796
rect 83829 66793 83841 66796
rect 83875 66793 83887 66827
rect 83829 66787 83887 66793
rect 85761 66827 85819 66833
rect 85761 66793 85773 66827
rect 85807 66824 85819 66827
rect 85807 66796 89208 66824
rect 85807 66793 85819 66796
rect 85761 66787 85819 66793
rect 83844 66688 83872 66787
rect 89180 66756 89208 66796
rect 89254 66784 89260 66836
rect 89312 66824 89318 66836
rect 91005 66827 91063 66833
rect 91005 66824 91017 66827
rect 89312 66796 91017 66824
rect 89312 66784 89318 66796
rect 91005 66793 91017 66796
rect 91051 66793 91063 66827
rect 91005 66787 91063 66793
rect 89346 66756 89352 66768
rect 89180 66728 89352 66756
rect 89346 66716 89352 66728
rect 89404 66716 89410 66768
rect 89993 66759 90051 66765
rect 89993 66756 90005 66759
rect 89640 66728 90005 66756
rect 84013 66691 84071 66697
rect 84013 66688 84025 66691
rect 83844 66660 84025 66688
rect 84013 66657 84025 66660
rect 84059 66657 84071 66691
rect 84013 66651 84071 66657
rect 87325 66691 87383 66697
rect 87325 66657 87337 66691
rect 87371 66688 87383 66691
rect 88150 66688 88156 66700
rect 87371 66660 88156 66688
rect 87371 66657 87383 66660
rect 87325 66651 87383 66657
rect 88150 66648 88156 66660
rect 88208 66688 88214 66700
rect 89162 66688 89168 66700
rect 88208 66660 89168 66688
rect 88208 66648 88214 66660
rect 89162 66648 89168 66660
rect 89220 66648 89226 66700
rect 89254 66580 89260 66632
rect 89312 66620 89318 66632
rect 89640 66629 89668 66728
rect 89993 66725 90005 66728
rect 90039 66725 90051 66759
rect 89993 66719 90051 66725
rect 90545 66759 90603 66765
rect 90545 66725 90557 66759
rect 90591 66725 90603 66759
rect 90545 66719 90603 66725
rect 89898 66648 89904 66700
rect 89956 66688 89962 66700
rect 90560 66688 90588 66719
rect 90634 66716 90640 66768
rect 90692 66756 90698 66768
rect 90692 66728 91784 66756
rect 90692 66716 90698 66728
rect 89956 66660 90312 66688
rect 90560 66660 91054 66688
rect 89956 66648 89962 66660
rect 90284 66632 90312 66660
rect 89625 66623 89683 66629
rect 89625 66620 89637 66623
rect 89312 66592 89637 66620
rect 89312 66580 89318 66592
rect 89625 66589 89637 66592
rect 89671 66589 89683 66623
rect 89625 66583 89683 66589
rect 89990 66580 89996 66632
rect 90048 66620 90054 66632
rect 90177 66623 90235 66629
rect 90177 66620 90189 66623
rect 90048 66592 90189 66620
rect 90048 66580 90054 66592
rect 90177 66589 90189 66592
rect 90223 66589 90235 66623
rect 90177 66583 90235 66589
rect 90266 66580 90272 66632
rect 90324 66580 90330 66632
rect 90634 66620 90640 66632
rect 90468 66592 90640 66620
rect 84286 66512 84292 66564
rect 84344 66512 84350 66564
rect 84378 66512 84384 66564
rect 84436 66552 84442 66564
rect 84436 66524 84778 66552
rect 84436 66512 84442 66524
rect 86954 66512 86960 66564
rect 87012 66552 87018 66564
rect 87012 66524 87722 66552
rect 87012 66512 87018 66524
rect 88886 66512 88892 66564
rect 88944 66512 88950 66564
rect 88978 66512 88984 66564
rect 89036 66552 89042 66564
rect 89346 66552 89352 66564
rect 89036 66524 89352 66552
rect 89036 66512 89042 66524
rect 89346 66512 89352 66524
rect 89404 66512 89410 66564
rect 90468 66552 90496 66592
rect 90634 66580 90640 66592
rect 90692 66580 90698 66632
rect 91026 66629 91054 66660
rect 91005 66623 91063 66629
rect 91005 66589 91017 66623
rect 91051 66589 91063 66623
rect 91005 66583 91063 66589
rect 91189 66623 91247 66629
rect 91189 66589 91201 66623
rect 91235 66620 91247 66623
rect 91278 66620 91284 66632
rect 91235 66592 91284 66620
rect 91235 66589 91247 66592
rect 91189 66583 91247 66589
rect 91278 66580 91284 66592
rect 91336 66580 91342 66632
rect 91370 66580 91376 66632
rect 91428 66620 91434 66632
rect 91756 66629 91784 66728
rect 91557 66623 91615 66629
rect 91557 66620 91569 66623
rect 91428 66592 91569 66620
rect 91428 66580 91434 66592
rect 91557 66589 91569 66592
rect 91603 66589 91615 66623
rect 91557 66583 91615 66589
rect 91741 66623 91799 66629
rect 91741 66589 91753 66623
rect 91787 66620 91799 66623
rect 102318 66620 102324 66632
rect 91787 66592 102324 66620
rect 91787 66589 91799 66592
rect 91741 66583 91799 66589
rect 102318 66580 102324 66592
rect 102376 66580 102382 66632
rect 89824 66524 90496 66552
rect 87417 66487 87475 66493
rect 87417 66453 87429 66487
rect 87463 66484 87475 66487
rect 88702 66484 88708 66496
rect 87463 66456 88708 66484
rect 87463 66453 87475 66456
rect 87417 66447 87475 66453
rect 88702 66444 88708 66456
rect 88760 66444 88766 66496
rect 89441 66487 89499 66493
rect 89441 66453 89453 66487
rect 89487 66484 89499 66487
rect 89714 66484 89720 66496
rect 89487 66456 89720 66484
rect 89487 66453 89499 66456
rect 89441 66447 89499 66453
rect 89714 66444 89720 66456
rect 89772 66444 89778 66496
rect 89824 66493 89852 66524
rect 90542 66512 90548 66564
rect 90600 66512 90606 66564
rect 90729 66555 90787 66561
rect 90729 66521 90741 66555
rect 90775 66521 90787 66555
rect 90729 66515 90787 66521
rect 90913 66555 90971 66561
rect 90913 66521 90925 66555
rect 90959 66552 90971 66555
rect 90959 66524 91968 66552
rect 90959 66521 90971 66524
rect 90913 66515 90971 66521
rect 89809 66487 89867 66493
rect 89809 66453 89821 66487
rect 89855 66453 89867 66487
rect 89809 66447 89867 66453
rect 89990 66444 89996 66496
rect 90048 66484 90054 66496
rect 90361 66487 90419 66493
rect 90361 66484 90373 66487
rect 90048 66456 90373 66484
rect 90048 66444 90054 66456
rect 90361 66453 90373 66456
rect 90407 66453 90419 66487
rect 90361 66447 90419 66453
rect 90450 66444 90456 66496
rect 90508 66484 90514 66496
rect 90744 66484 90772 66515
rect 91940 66496 91968 66524
rect 91373 66487 91431 66493
rect 91373 66484 91385 66487
rect 90508 66456 91385 66484
rect 90508 66444 90514 66456
rect 91373 66453 91385 66456
rect 91419 66453 91431 66487
rect 91373 66447 91431 66453
rect 91922 66444 91928 66496
rect 91980 66444 91986 66496
rect 1104 66394 108836 66416
rect 1104 66342 4874 66394
rect 4926 66342 4938 66394
rect 4990 66342 5002 66394
rect 5054 66342 5066 66394
rect 5118 66342 5130 66394
rect 5182 66342 35594 66394
rect 35646 66342 35658 66394
rect 35710 66342 35722 66394
rect 35774 66342 35786 66394
rect 35838 66342 35850 66394
rect 35902 66342 66314 66394
rect 66366 66342 66378 66394
rect 66430 66342 66442 66394
rect 66494 66342 66506 66394
rect 66558 66342 66570 66394
rect 66622 66342 97034 66394
rect 97086 66342 97098 66394
rect 97150 66342 97162 66394
rect 97214 66342 97226 66394
rect 97278 66342 97290 66394
rect 97342 66342 106658 66394
rect 106710 66342 106722 66394
rect 106774 66342 106786 66394
rect 106838 66342 106850 66394
rect 106902 66342 106914 66394
rect 106966 66342 108836 66394
rect 1104 66320 108836 66342
rect 84286 66240 84292 66292
rect 84344 66280 84350 66292
rect 85209 66283 85267 66289
rect 85209 66280 85221 66283
rect 84344 66252 85221 66280
rect 84344 66240 84350 66252
rect 85209 66249 85221 66252
rect 85255 66249 85267 66283
rect 85209 66243 85267 66249
rect 88426 66240 88432 66292
rect 88484 66240 88490 66292
rect 89257 66283 89315 66289
rect 89257 66249 89269 66283
rect 89303 66280 89315 66283
rect 89438 66280 89444 66292
rect 89303 66252 89444 66280
rect 89303 66249 89315 66252
rect 89257 66243 89315 66249
rect 89438 66240 89444 66252
rect 89496 66240 89502 66292
rect 89714 66240 89720 66292
rect 89772 66280 89778 66292
rect 89898 66280 89904 66292
rect 89772 66252 89904 66280
rect 89772 66240 89778 66252
rect 89898 66240 89904 66252
rect 89956 66240 89962 66292
rect 89990 66240 89996 66292
rect 90048 66280 90054 66292
rect 90726 66280 90732 66292
rect 90048 66252 90732 66280
rect 90048 66240 90054 66252
rect 90726 66240 90732 66252
rect 90784 66240 90790 66292
rect 91002 66240 91008 66292
rect 91060 66240 91066 66292
rect 91370 66280 91376 66292
rect 91112 66252 91376 66280
rect 36078 66172 36084 66224
rect 36136 66172 36142 66224
rect 37918 66172 37924 66224
rect 37976 66212 37982 66224
rect 38470 66212 38476 66224
rect 37976 66184 38476 66212
rect 37976 66172 37982 66184
rect 38470 66172 38476 66184
rect 38528 66212 38534 66224
rect 38657 66215 38715 66221
rect 38657 66212 38669 66215
rect 38528 66184 38669 66212
rect 38528 66172 38534 66184
rect 38657 66181 38669 66184
rect 38703 66181 38715 66215
rect 38657 66175 38715 66181
rect 41138 66172 41144 66224
rect 41196 66172 41202 66224
rect 43622 66172 43628 66224
rect 43680 66172 43686 66224
rect 46106 66172 46112 66224
rect 46164 66172 46170 66224
rect 48590 66172 48596 66224
rect 48648 66172 48654 66224
rect 51074 66172 51080 66224
rect 51132 66172 51138 66224
rect 53558 66172 53564 66224
rect 53616 66172 53622 66224
rect 56134 66172 56140 66224
rect 56192 66172 56198 66224
rect 58618 66172 58624 66224
rect 58676 66172 58682 66224
rect 61102 66172 61108 66224
rect 61160 66172 61166 66224
rect 63586 66172 63592 66224
rect 63644 66172 63650 66224
rect 66070 66172 66076 66224
rect 66128 66172 66134 66224
rect 68554 66172 68560 66224
rect 68612 66172 68618 66224
rect 71038 66172 71044 66224
rect 71096 66172 71102 66224
rect 73522 66172 73528 66224
rect 73580 66172 73586 66224
rect 85574 66172 85580 66224
rect 85632 66212 85638 66224
rect 85632 66184 86526 66212
rect 85632 66172 85638 66184
rect 87598 66172 87604 66224
rect 87656 66212 87662 66224
rect 88061 66215 88119 66221
rect 88061 66212 88073 66215
rect 87656 66184 88073 66212
rect 87656 66172 87662 66184
rect 88061 66181 88073 66184
rect 88107 66181 88119 66215
rect 88061 66175 88119 66181
rect 88245 66215 88303 66221
rect 88245 66181 88257 66215
rect 88291 66212 88303 66215
rect 89533 66215 89591 66221
rect 89533 66212 89545 66215
rect 88291 66184 89545 66212
rect 88291 66181 88303 66184
rect 88245 66175 88303 66181
rect 89533 66181 89545 66184
rect 89579 66181 89591 66215
rect 90450 66212 90456 66224
rect 89533 66175 89591 66181
rect 89640 66184 90456 66212
rect 85666 66104 85672 66156
rect 85724 66104 85730 66156
rect 87969 66147 88027 66153
rect 87969 66113 87981 66147
rect 88015 66144 88027 66147
rect 88150 66144 88156 66156
rect 88015 66116 88156 66144
rect 88015 66113 88027 66116
rect 87969 66107 88027 66113
rect 88150 66104 88156 66116
rect 88208 66104 88214 66156
rect 88337 66147 88395 66153
rect 88337 66113 88349 66147
rect 88383 66144 88395 66147
rect 89349 66147 89407 66153
rect 88383 66116 89208 66144
rect 88383 66113 88395 66116
rect 88337 66107 88395 66113
rect 85684 66076 85712 66104
rect 87598 66076 87604 66088
rect 85684 66048 87604 66076
rect 87598 66036 87604 66048
rect 87656 66036 87662 66088
rect 87693 66079 87751 66085
rect 87693 66045 87705 66079
rect 87739 66076 87751 66079
rect 87739 66048 88012 66076
rect 87739 66045 87751 66048
rect 87693 66039 87751 66045
rect 85393 66011 85451 66017
rect 85393 65977 85405 66011
rect 85439 66008 85451 66011
rect 87984 66008 88012 66048
rect 88058 66036 88064 66088
rect 88116 66076 88122 66088
rect 88797 66079 88855 66085
rect 88797 66076 88809 66079
rect 88116 66048 88809 66076
rect 88116 66036 88122 66048
rect 88797 66045 88809 66048
rect 88843 66045 88855 66079
rect 88797 66039 88855 66045
rect 88978 66036 88984 66088
rect 89036 66036 89042 66088
rect 89073 66079 89131 66085
rect 89073 66045 89085 66079
rect 89119 66045 89131 66079
rect 89180 66076 89208 66116
rect 89349 66113 89361 66147
rect 89395 66144 89407 66147
rect 89640 66144 89668 66184
rect 89916 66153 89944 66184
rect 90450 66172 90456 66184
rect 90508 66172 90514 66224
rect 90637 66215 90695 66221
rect 90637 66181 90649 66215
rect 90683 66212 90695 66215
rect 90910 66212 90916 66224
rect 90683 66184 90916 66212
rect 90683 66181 90695 66184
rect 90637 66175 90695 66181
rect 90910 66172 90916 66184
rect 90968 66172 90974 66224
rect 89395 66116 89668 66144
rect 89717 66147 89775 66153
rect 89395 66113 89407 66116
rect 89349 66107 89407 66113
rect 89717 66113 89729 66147
rect 89763 66113 89775 66147
rect 89717 66107 89775 66113
rect 89901 66147 89959 66153
rect 89901 66113 89913 66147
rect 89947 66113 89959 66147
rect 89901 66107 89959 66113
rect 89438 66076 89444 66088
rect 89180 66048 89444 66076
rect 89073 66039 89131 66045
rect 88613 66011 88671 66017
rect 85439 65980 86724 66008
rect 87984 65980 88564 66008
rect 85439 65977 85451 65980
rect 85393 65971 85451 65977
rect 86218 65900 86224 65952
rect 86276 65900 86282 65952
rect 86696 65940 86724 65980
rect 87874 65940 87880 65952
rect 86696 65912 87880 65940
rect 87874 65900 87880 65912
rect 87932 65900 87938 65952
rect 88536 65940 88564 65980
rect 88613 65977 88625 66011
rect 88659 66008 88671 66011
rect 89088 66008 89116 66039
rect 89438 66036 89444 66048
rect 89496 66036 89502 66088
rect 89732 66076 89760 66107
rect 90358 66104 90364 66156
rect 90416 66142 90422 66156
rect 90821 66147 90879 66153
rect 90821 66144 90833 66147
rect 90468 66142 90833 66144
rect 90416 66116 90833 66142
rect 90416 66114 90496 66116
rect 90416 66104 90422 66114
rect 90821 66113 90833 66116
rect 90867 66144 90879 66147
rect 91112 66144 91140 66252
rect 91370 66240 91376 66252
rect 91428 66240 91434 66292
rect 91922 66240 91928 66292
rect 91980 66280 91986 66292
rect 102134 66280 102140 66292
rect 91980 66252 102140 66280
rect 91980 66240 91986 66252
rect 102134 66240 102140 66252
rect 102192 66240 102198 66292
rect 91554 66221 91560 66224
rect 91541 66215 91560 66221
rect 91541 66181 91553 66215
rect 91541 66175 91560 66181
rect 91554 66172 91560 66175
rect 91612 66172 91618 66224
rect 91741 66215 91799 66221
rect 91741 66181 91753 66215
rect 91787 66181 91799 66215
rect 91741 66175 91799 66181
rect 90867 66116 91140 66144
rect 90867 66113 90879 66116
rect 90821 66107 90879 66113
rect 91186 66104 91192 66156
rect 91244 66104 91250 66156
rect 89548 66048 89760 66076
rect 90453 66079 90511 66085
rect 89254 66008 89260 66020
rect 88659 65980 89260 66008
rect 88659 65977 88671 65980
rect 88613 65971 88671 65977
rect 89254 65968 89260 65980
rect 89312 65968 89318 66020
rect 89346 65968 89352 66020
rect 89404 66008 89410 66020
rect 89548 66008 89576 66048
rect 90453 66045 90465 66079
rect 90499 66076 90511 66079
rect 90634 66076 90640 66088
rect 90499 66048 90640 66076
rect 90499 66045 90511 66048
rect 90453 66039 90511 66045
rect 90634 66036 90640 66048
rect 90692 66036 90698 66088
rect 90726 66036 90732 66088
rect 90784 66076 90790 66088
rect 90784 66048 91140 66076
rect 90784 66036 90790 66048
rect 89404 65980 89576 66008
rect 91112 66008 91140 66048
rect 91756 66008 91784 66175
rect 94314 66172 94320 66224
rect 94372 66212 94378 66224
rect 94409 66215 94467 66221
rect 94409 66212 94421 66215
rect 94372 66184 94421 66212
rect 94372 66172 94378 66184
rect 94409 66181 94421 66184
rect 94455 66181 94467 66215
rect 94409 66175 94467 66181
rect 91922 66104 91928 66156
rect 91980 66104 91986 66156
rect 91112 65980 91784 66008
rect 89404 65968 89410 65980
rect 89993 65943 90051 65949
rect 89993 65940 90005 65943
rect 88536 65912 90005 65940
rect 89993 65909 90005 65912
rect 90039 65909 90051 65943
rect 89993 65903 90051 65909
rect 90634 65900 90640 65952
rect 90692 65940 90698 65952
rect 91278 65940 91284 65952
rect 90692 65912 91284 65940
rect 90692 65900 90698 65912
rect 91278 65900 91284 65912
rect 91336 65940 91342 65952
rect 91373 65943 91431 65949
rect 91373 65940 91385 65943
rect 91336 65912 91385 65940
rect 91336 65900 91342 65912
rect 91373 65909 91385 65912
rect 91419 65909 91431 65943
rect 91373 65903 91431 65909
rect 91554 65900 91560 65952
rect 91612 65900 91618 65952
rect 92017 65943 92075 65949
rect 92017 65909 92029 65943
rect 92063 65940 92075 65943
rect 92290 65940 92296 65952
rect 92063 65912 92296 65940
rect 92063 65909 92075 65912
rect 92017 65903 92075 65909
rect 92290 65900 92296 65912
rect 92348 65900 92354 65952
rect 95878 65900 95884 65952
rect 95936 65940 95942 65952
rect 96249 65943 96307 65949
rect 96249 65940 96261 65943
rect 95936 65912 96261 65940
rect 95936 65900 95942 65912
rect 96249 65909 96261 65912
rect 96295 65940 96307 65943
rect 96525 65943 96583 65949
rect 96525 65940 96537 65943
rect 96295 65912 96537 65940
rect 96295 65909 96307 65912
rect 96249 65903 96307 65909
rect 96525 65909 96537 65912
rect 96571 65909 96583 65943
rect 96525 65903 96583 65909
rect 1104 65850 108836 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 96374 65850
rect 96426 65798 96438 65850
rect 96490 65798 96502 65850
rect 96554 65798 96566 65850
rect 96618 65798 96630 65850
rect 96682 65798 105922 65850
rect 105974 65798 105986 65850
rect 106038 65798 106050 65850
rect 106102 65798 106114 65850
rect 106166 65798 106178 65850
rect 106230 65798 108836 65850
rect 1104 65776 108836 65798
rect 86218 65696 86224 65748
rect 86276 65736 86282 65748
rect 90358 65736 90364 65748
rect 86276 65708 90364 65736
rect 86276 65696 86282 65708
rect 90358 65696 90364 65708
rect 90416 65696 90422 65748
rect 90542 65696 90548 65748
rect 90600 65736 90606 65748
rect 91554 65736 91560 65748
rect 90600 65708 91560 65736
rect 90600 65696 90606 65708
rect 91554 65696 91560 65708
rect 91612 65696 91618 65748
rect 88426 65628 88432 65680
rect 88484 65668 88490 65680
rect 91186 65668 91192 65680
rect 88484 65640 91192 65668
rect 88484 65628 88490 65640
rect 91186 65628 91192 65640
rect 91244 65628 91250 65680
rect 92290 65628 92296 65680
rect 92348 65668 92354 65680
rect 103514 65668 103520 65680
rect 92348 65640 103520 65668
rect 92348 65628 92354 65640
rect 103514 65628 103520 65640
rect 103572 65628 103578 65680
rect 89806 65492 89812 65544
rect 89864 65532 89870 65544
rect 103606 65532 103612 65544
rect 89864 65504 103612 65532
rect 89864 65492 89870 65504
rect 103606 65492 103612 65504
rect 103664 65492 103670 65544
rect 1104 65306 7912 65328
rect 1104 65254 4874 65306
rect 4926 65254 4938 65306
rect 4990 65254 5002 65306
rect 5054 65254 5066 65306
rect 5118 65254 5130 65306
rect 5182 65254 7912 65306
rect 1104 65232 7912 65254
rect 104052 65306 108836 65328
rect 104052 65254 106658 65306
rect 106710 65254 106722 65306
rect 106774 65254 106786 65306
rect 106838 65254 106850 65306
rect 106902 65254 106914 65306
rect 106966 65254 108836 65306
rect 104052 65232 108836 65254
rect 1104 64762 7912 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 7912 64762
rect 1104 64688 7912 64710
rect 104052 64762 108836 64784
rect 104052 64710 105922 64762
rect 105974 64710 105986 64762
rect 106038 64710 106050 64762
rect 106102 64710 106114 64762
rect 106166 64710 106178 64762
rect 106230 64710 108836 64762
rect 104052 64688 108836 64710
rect 1104 64218 7912 64240
rect 1104 64166 4874 64218
rect 4926 64166 4938 64218
rect 4990 64166 5002 64218
rect 5054 64166 5066 64218
rect 5118 64166 5130 64218
rect 5182 64166 7912 64218
rect 1104 64144 7912 64166
rect 104052 64218 108836 64240
rect 104052 64166 106658 64218
rect 106710 64166 106722 64218
rect 106774 64166 106786 64218
rect 106838 64166 106850 64218
rect 106902 64166 106914 64218
rect 106966 64166 108836 64218
rect 104052 64144 108836 64166
rect 1104 63674 7912 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 7912 63674
rect 1104 63600 7912 63622
rect 104052 63674 108836 63696
rect 104052 63622 105922 63674
rect 105974 63622 105986 63674
rect 106038 63622 106050 63674
rect 106102 63622 106114 63674
rect 106166 63622 106178 63674
rect 106230 63622 108836 63674
rect 104052 63600 108836 63622
rect 1104 63130 7912 63152
rect 1104 63078 4874 63130
rect 4926 63078 4938 63130
rect 4990 63078 5002 63130
rect 5054 63078 5066 63130
rect 5118 63078 5130 63130
rect 5182 63078 7912 63130
rect 1104 63056 7912 63078
rect 104052 63130 108836 63152
rect 104052 63078 106658 63130
rect 106710 63078 106722 63130
rect 106774 63078 106786 63130
rect 106838 63078 106850 63130
rect 106902 63078 106914 63130
rect 106966 63078 108836 63130
rect 104052 63056 108836 63078
rect 1104 62586 7912 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 7912 62586
rect 1104 62512 7912 62534
rect 104052 62586 108836 62608
rect 104052 62534 105922 62586
rect 105974 62534 105986 62586
rect 106038 62534 106050 62586
rect 106102 62534 106114 62586
rect 106166 62534 106178 62586
rect 106230 62534 108836 62586
rect 104052 62512 108836 62534
rect 1104 62042 7912 62064
rect 1104 61990 4874 62042
rect 4926 61990 4938 62042
rect 4990 61990 5002 62042
rect 5054 61990 5066 62042
rect 5118 61990 5130 62042
rect 5182 61990 7912 62042
rect 1104 61968 7912 61990
rect 104052 62042 108836 62064
rect 104052 61990 106658 62042
rect 106710 61990 106722 62042
rect 106774 61990 106786 62042
rect 106838 61990 106850 62042
rect 106902 61990 106914 62042
rect 106966 61990 108836 62042
rect 104052 61968 108836 61990
rect 1104 61498 7912 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 7912 61498
rect 1104 61424 7912 61446
rect 104052 61498 108836 61520
rect 104052 61446 105922 61498
rect 105974 61446 105986 61498
rect 106038 61446 106050 61498
rect 106102 61446 106114 61498
rect 106166 61446 106178 61498
rect 106230 61446 108836 61498
rect 104052 61424 108836 61446
rect 1104 60954 7912 60976
rect 1104 60902 4874 60954
rect 4926 60902 4938 60954
rect 4990 60902 5002 60954
rect 5054 60902 5066 60954
rect 5118 60902 5130 60954
rect 5182 60902 7912 60954
rect 1104 60880 7912 60902
rect 104052 60954 108836 60976
rect 104052 60902 106658 60954
rect 106710 60902 106722 60954
rect 106774 60902 106786 60954
rect 106838 60902 106850 60954
rect 106902 60902 106914 60954
rect 106966 60902 108836 60954
rect 104052 60880 108836 60902
rect 7282 60664 7288 60716
rect 7340 60664 7346 60716
rect 6822 60596 6828 60648
rect 6880 60636 6886 60648
rect 7469 60639 7527 60645
rect 7469 60636 7481 60639
rect 6880 60608 7481 60636
rect 6880 60596 6886 60608
rect 7469 60605 7481 60608
rect 7515 60605 7527 60639
rect 7469 60599 7527 60605
rect 1104 60410 7912 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 7912 60410
rect 1104 60336 7912 60358
rect 104052 60410 108836 60432
rect 104052 60358 105922 60410
rect 105974 60358 105986 60410
rect 106038 60358 106050 60410
rect 106102 60358 106114 60410
rect 106166 60358 106178 60410
rect 106230 60358 108836 60410
rect 104052 60336 108836 60358
rect 6273 60299 6331 60305
rect 6273 60265 6285 60299
rect 6319 60296 6331 60299
rect 6822 60296 6828 60308
rect 6319 60268 6828 60296
rect 6319 60265 6331 60268
rect 6273 60259 6331 60265
rect 6822 60256 6828 60268
rect 6880 60256 6886 60308
rect 7282 60052 7288 60104
rect 7340 60092 7346 60104
rect 7561 60095 7619 60101
rect 7561 60092 7573 60095
rect 7340 60064 7573 60092
rect 7340 60052 7346 60064
rect 7561 60061 7573 60064
rect 7607 60061 7619 60095
rect 7561 60055 7619 60061
rect 104342 60052 104348 60104
rect 104400 60052 104406 60104
rect 1104 59866 7912 59888
rect 1104 59814 4874 59866
rect 4926 59814 4938 59866
rect 4990 59814 5002 59866
rect 5054 59814 5066 59866
rect 5118 59814 5130 59866
rect 5182 59814 7912 59866
rect 1104 59792 7912 59814
rect 104052 59866 108836 59888
rect 104052 59814 106658 59866
rect 106710 59814 106722 59866
rect 106774 59814 106786 59866
rect 106838 59814 106850 59866
rect 106902 59814 106914 59866
rect 106966 59814 108836 59866
rect 104052 59792 108836 59814
rect 6822 59712 6828 59764
rect 6880 59752 6886 59764
rect 6917 59755 6975 59761
rect 6917 59752 6929 59755
rect 6880 59724 6929 59752
rect 6880 59712 6886 59724
rect 6917 59721 6929 59724
rect 6963 59752 6975 59755
rect 6963 59724 7236 59752
rect 6963 59721 6975 59724
rect 6917 59715 6975 59721
rect 7208 59693 7236 59724
rect 7193 59687 7251 59693
rect 7193 59653 7205 59687
rect 7239 59653 7251 59687
rect 7193 59647 7251 59653
rect 1104 59322 7912 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 7912 59322
rect 1104 59248 7912 59270
rect 104052 59322 108836 59344
rect 104052 59270 105922 59322
rect 105974 59270 105986 59322
rect 106038 59270 106050 59322
rect 106102 59270 106114 59322
rect 106166 59270 106178 59322
rect 106230 59270 108836 59322
rect 104052 59248 108836 59270
rect 1104 58778 7912 58800
rect 1104 58726 4874 58778
rect 4926 58726 4938 58778
rect 4990 58726 5002 58778
rect 5054 58726 5066 58778
rect 5118 58726 5130 58778
rect 5182 58726 7912 58778
rect 1104 58704 7912 58726
rect 104052 58778 108836 58800
rect 104052 58726 106658 58778
rect 106710 58726 106722 58778
rect 106774 58726 106786 58778
rect 106838 58726 106850 58778
rect 106902 58726 106914 58778
rect 106966 58726 108836 58778
rect 104052 58704 108836 58726
rect 1104 58234 7912 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 7912 58234
rect 1104 58160 7912 58182
rect 104052 58234 108836 58256
rect 104052 58182 105922 58234
rect 105974 58182 105986 58234
rect 106038 58182 106050 58234
rect 106102 58182 106114 58234
rect 106166 58182 106178 58234
rect 106230 58182 108836 58234
rect 104052 58160 108836 58182
rect 1104 57690 7912 57712
rect 1104 57638 4874 57690
rect 4926 57638 4938 57690
rect 4990 57638 5002 57690
rect 5054 57638 5066 57690
rect 5118 57638 5130 57690
rect 5182 57638 7912 57690
rect 1104 57616 7912 57638
rect 104052 57690 108836 57712
rect 104052 57638 106658 57690
rect 106710 57638 106722 57690
rect 106774 57638 106786 57690
rect 106838 57638 106850 57690
rect 106902 57638 106914 57690
rect 106966 57638 108836 57690
rect 104052 57616 108836 57638
rect 1104 57146 7912 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 7912 57146
rect 1104 57072 7912 57094
rect 104052 57146 108836 57168
rect 104052 57094 105922 57146
rect 105974 57094 105986 57146
rect 106038 57094 106050 57146
rect 106102 57094 106114 57146
rect 106166 57094 106178 57146
rect 106230 57094 108836 57146
rect 104052 57072 108836 57094
rect 1104 56602 7912 56624
rect 1104 56550 4874 56602
rect 4926 56550 4938 56602
rect 4990 56550 5002 56602
rect 5054 56550 5066 56602
rect 5118 56550 5130 56602
rect 5182 56550 7912 56602
rect 1104 56528 7912 56550
rect 104052 56602 108836 56624
rect 104052 56550 106658 56602
rect 106710 56550 106722 56602
rect 106774 56550 106786 56602
rect 106838 56550 106850 56602
rect 106902 56550 106914 56602
rect 106966 56550 108836 56602
rect 104052 56528 108836 56550
rect 1104 56058 7912 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 7912 56058
rect 1104 55984 7912 56006
rect 104052 56058 108836 56080
rect 104052 56006 105922 56058
rect 105974 56006 105986 56058
rect 106038 56006 106050 56058
rect 106102 56006 106114 56058
rect 106166 56006 106178 56058
rect 106230 56006 108836 56058
rect 104052 55984 108836 56006
rect 1104 55514 7912 55536
rect 1104 55462 4874 55514
rect 4926 55462 4938 55514
rect 4990 55462 5002 55514
rect 5054 55462 5066 55514
rect 5118 55462 5130 55514
rect 5182 55462 7912 55514
rect 1104 55440 7912 55462
rect 104052 55514 108836 55536
rect 104052 55462 106658 55514
rect 106710 55462 106722 55514
rect 106774 55462 106786 55514
rect 106838 55462 106850 55514
rect 106902 55462 106914 55514
rect 106966 55462 108836 55514
rect 104052 55440 108836 55462
rect 1104 54970 7912 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 7912 54970
rect 1104 54896 7912 54918
rect 104052 54970 108836 54992
rect 104052 54918 105922 54970
rect 105974 54918 105986 54970
rect 106038 54918 106050 54970
rect 106102 54918 106114 54970
rect 106166 54918 106178 54970
rect 106230 54918 108836 54970
rect 104052 54896 108836 54918
rect 1104 54426 7912 54448
rect 1104 54374 4874 54426
rect 4926 54374 4938 54426
rect 4990 54374 5002 54426
rect 5054 54374 5066 54426
rect 5118 54374 5130 54426
rect 5182 54374 7912 54426
rect 1104 54352 7912 54374
rect 104052 54426 108836 54448
rect 104052 54374 106658 54426
rect 106710 54374 106722 54426
rect 106774 54374 106786 54426
rect 106838 54374 106850 54426
rect 106902 54374 106914 54426
rect 106966 54374 108836 54426
rect 104052 54352 108836 54374
rect 1104 53882 7912 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 7912 53882
rect 1104 53808 7912 53830
rect 104052 53882 108836 53904
rect 104052 53830 105922 53882
rect 105974 53830 105986 53882
rect 106038 53830 106050 53882
rect 106102 53830 106114 53882
rect 106166 53830 106178 53882
rect 106230 53830 108836 53882
rect 104052 53808 108836 53830
rect 1104 53338 7912 53360
rect 1104 53286 4874 53338
rect 4926 53286 4938 53338
rect 4990 53286 5002 53338
rect 5054 53286 5066 53338
rect 5118 53286 5130 53338
rect 5182 53286 7912 53338
rect 1104 53264 7912 53286
rect 104052 53338 108836 53360
rect 104052 53286 106658 53338
rect 106710 53286 106722 53338
rect 106774 53286 106786 53338
rect 106838 53286 106850 53338
rect 106902 53286 106914 53338
rect 106966 53286 108836 53338
rect 104052 53264 108836 53286
rect 1104 52794 7912 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 7912 52794
rect 1104 52720 7912 52742
rect 104052 52794 108836 52816
rect 104052 52742 105922 52794
rect 105974 52742 105986 52794
rect 106038 52742 106050 52794
rect 106102 52742 106114 52794
rect 106166 52742 106178 52794
rect 106230 52742 108836 52794
rect 104052 52720 108836 52742
rect 1104 52250 7912 52272
rect 1104 52198 4874 52250
rect 4926 52198 4938 52250
rect 4990 52198 5002 52250
rect 5054 52198 5066 52250
rect 5118 52198 5130 52250
rect 5182 52198 7912 52250
rect 1104 52176 7912 52198
rect 104052 52250 108836 52272
rect 104052 52198 106658 52250
rect 106710 52198 106722 52250
rect 106774 52198 106786 52250
rect 106838 52198 106850 52250
rect 106902 52198 106914 52250
rect 106966 52198 108836 52250
rect 104052 52176 108836 52198
rect 1104 51706 7912 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 7912 51706
rect 1104 51632 7912 51654
rect 104052 51706 108836 51728
rect 104052 51654 105922 51706
rect 105974 51654 105986 51706
rect 106038 51654 106050 51706
rect 106102 51654 106114 51706
rect 106166 51654 106178 51706
rect 106230 51654 108836 51706
rect 104052 51632 108836 51654
rect 1104 51162 7912 51184
rect 1104 51110 4874 51162
rect 4926 51110 4938 51162
rect 4990 51110 5002 51162
rect 5054 51110 5066 51162
rect 5118 51110 5130 51162
rect 5182 51110 7912 51162
rect 1104 51088 7912 51110
rect 104052 51162 108836 51184
rect 104052 51110 106658 51162
rect 106710 51110 106722 51162
rect 106774 51110 106786 51162
rect 106838 51110 106850 51162
rect 106902 51110 106914 51162
rect 106966 51110 108836 51162
rect 104052 51088 108836 51110
rect 1104 50618 7912 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 7912 50618
rect 1104 50544 7912 50566
rect 104052 50618 108836 50640
rect 104052 50566 105922 50618
rect 105974 50566 105986 50618
rect 106038 50566 106050 50618
rect 106102 50566 106114 50618
rect 106166 50566 106178 50618
rect 106230 50566 108836 50618
rect 104052 50544 108836 50566
rect 1104 50074 7912 50096
rect 1104 50022 4874 50074
rect 4926 50022 4938 50074
rect 4990 50022 5002 50074
rect 5054 50022 5066 50074
rect 5118 50022 5130 50074
rect 5182 50022 7912 50074
rect 1104 50000 7912 50022
rect 104052 50074 108836 50096
rect 104052 50022 106658 50074
rect 106710 50022 106722 50074
rect 106774 50022 106786 50074
rect 106838 50022 106850 50074
rect 106902 50022 106914 50074
rect 106966 50022 108836 50074
rect 104052 50000 108836 50022
rect 1104 49530 7912 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 7912 49530
rect 1104 49456 7912 49478
rect 104052 49530 108836 49552
rect 104052 49478 105922 49530
rect 105974 49478 105986 49530
rect 106038 49478 106050 49530
rect 106102 49478 106114 49530
rect 106166 49478 106178 49530
rect 106230 49478 108836 49530
rect 104052 49456 108836 49478
rect 1104 48986 7912 49008
rect 1104 48934 4874 48986
rect 4926 48934 4938 48986
rect 4990 48934 5002 48986
rect 5054 48934 5066 48986
rect 5118 48934 5130 48986
rect 5182 48934 7912 48986
rect 1104 48912 7912 48934
rect 104052 48986 108836 49008
rect 104052 48934 106658 48986
rect 106710 48934 106722 48986
rect 106774 48934 106786 48986
rect 106838 48934 106850 48986
rect 106902 48934 106914 48986
rect 106966 48934 108836 48986
rect 104052 48912 108836 48934
rect 1104 48442 7912 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 7912 48442
rect 1104 48368 7912 48390
rect 104052 48442 108836 48464
rect 104052 48390 105922 48442
rect 105974 48390 105986 48442
rect 106038 48390 106050 48442
rect 106102 48390 106114 48442
rect 106166 48390 106178 48442
rect 106230 48390 108836 48442
rect 104052 48368 108836 48390
rect 1104 47898 7912 47920
rect 1104 47846 4874 47898
rect 4926 47846 4938 47898
rect 4990 47846 5002 47898
rect 5054 47846 5066 47898
rect 5118 47846 5130 47898
rect 5182 47846 7912 47898
rect 1104 47824 7912 47846
rect 104052 47898 108836 47920
rect 104052 47846 106658 47898
rect 106710 47846 106722 47898
rect 106774 47846 106786 47898
rect 106838 47846 106850 47898
rect 106902 47846 106914 47898
rect 106966 47846 108836 47898
rect 104052 47824 108836 47846
rect 1104 47354 7912 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 7912 47354
rect 1104 47280 7912 47302
rect 104052 47354 108836 47376
rect 104052 47302 105922 47354
rect 105974 47302 105986 47354
rect 106038 47302 106050 47354
rect 106102 47302 106114 47354
rect 106166 47302 106178 47354
rect 106230 47302 108836 47354
rect 104052 47280 108836 47302
rect 1104 46810 7912 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 7912 46810
rect 1104 46736 7912 46758
rect 104052 46810 108836 46832
rect 104052 46758 106658 46810
rect 106710 46758 106722 46810
rect 106774 46758 106786 46810
rect 106838 46758 106850 46810
rect 106902 46758 106914 46810
rect 106966 46758 108836 46810
rect 104052 46736 108836 46758
rect 1104 46266 7912 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 7912 46266
rect 1104 46192 7912 46214
rect 104052 46266 108836 46288
rect 104052 46214 105922 46266
rect 105974 46214 105986 46266
rect 106038 46214 106050 46266
rect 106102 46214 106114 46266
rect 106166 46214 106178 46266
rect 106230 46214 108836 46266
rect 104052 46192 108836 46214
rect 1104 45722 7912 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 7912 45722
rect 1104 45648 7912 45670
rect 104052 45722 108836 45744
rect 104052 45670 106658 45722
rect 106710 45670 106722 45722
rect 106774 45670 106786 45722
rect 106838 45670 106850 45722
rect 106902 45670 106914 45722
rect 106966 45670 108836 45722
rect 104052 45648 108836 45670
rect 1104 45178 7912 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 7912 45178
rect 1104 45104 7912 45126
rect 104052 45178 108836 45200
rect 104052 45126 105922 45178
rect 105974 45126 105986 45178
rect 106038 45126 106050 45178
rect 106102 45126 106114 45178
rect 106166 45126 106178 45178
rect 106230 45126 108836 45178
rect 104052 45104 108836 45126
rect 1104 44634 7912 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 7912 44634
rect 1104 44560 7912 44582
rect 104052 44634 108836 44656
rect 104052 44582 106658 44634
rect 106710 44582 106722 44634
rect 106774 44582 106786 44634
rect 106838 44582 106850 44634
rect 106902 44582 106914 44634
rect 106966 44582 108836 44634
rect 104052 44560 108836 44582
rect 1104 44090 7912 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 7912 44090
rect 1104 44016 7912 44038
rect 104052 44090 108836 44112
rect 104052 44038 105922 44090
rect 105974 44038 105986 44090
rect 106038 44038 106050 44090
rect 106102 44038 106114 44090
rect 106166 44038 106178 44090
rect 106230 44038 108836 44090
rect 104052 44016 108836 44038
rect 1104 43546 7912 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 7912 43546
rect 1104 43472 7912 43494
rect 104052 43546 108836 43568
rect 104052 43494 106658 43546
rect 106710 43494 106722 43546
rect 106774 43494 106786 43546
rect 106838 43494 106850 43546
rect 106902 43494 106914 43546
rect 106966 43494 108836 43546
rect 104052 43472 108836 43494
rect 1104 43002 7912 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 7912 43002
rect 1104 42928 7912 42950
rect 104052 43002 108836 43024
rect 104052 42950 105922 43002
rect 105974 42950 105986 43002
rect 106038 42950 106050 43002
rect 106102 42950 106114 43002
rect 106166 42950 106178 43002
rect 106230 42950 108836 43002
rect 104052 42928 108836 42950
rect 1104 42458 7912 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 7912 42458
rect 1104 42384 7912 42406
rect 104052 42458 108836 42480
rect 104052 42406 106658 42458
rect 106710 42406 106722 42458
rect 106774 42406 106786 42458
rect 106838 42406 106850 42458
rect 106902 42406 106914 42458
rect 106966 42406 108836 42458
rect 104052 42384 108836 42406
rect 1104 41914 7912 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 7912 41914
rect 1104 41840 7912 41862
rect 104052 41914 108836 41936
rect 104052 41862 105922 41914
rect 105974 41862 105986 41914
rect 106038 41862 106050 41914
rect 106102 41862 106114 41914
rect 106166 41862 106178 41914
rect 106230 41862 108836 41914
rect 104052 41840 108836 41862
rect 7558 41420 7564 41472
rect 7616 41420 7622 41472
rect 1104 41370 7912 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 7912 41370
rect 1104 41296 7912 41318
rect 104052 41370 108836 41392
rect 104052 41318 106658 41370
rect 106710 41318 106722 41370
rect 106774 41318 106786 41370
rect 106838 41318 106850 41370
rect 106902 41318 106914 41370
rect 106966 41318 108836 41370
rect 104052 41296 108836 41318
rect 1104 40826 7912 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 7912 40826
rect 1104 40752 7912 40774
rect 104052 40826 108836 40848
rect 104052 40774 105922 40826
rect 105974 40774 105986 40826
rect 106038 40774 106050 40826
rect 106102 40774 106114 40826
rect 106166 40774 106178 40826
rect 106230 40774 108836 40826
rect 104052 40752 108836 40774
rect 1104 40282 7912 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 7912 40282
rect 1104 40208 7912 40230
rect 104052 40282 108836 40304
rect 104052 40230 106658 40282
rect 106710 40230 106722 40282
rect 106774 40230 106786 40282
rect 106838 40230 106850 40282
rect 106902 40230 106914 40282
rect 106966 40230 108836 40282
rect 104052 40208 108836 40230
rect 3418 39992 3424 40044
rect 3476 40032 3482 40044
rect 7558 40032 7564 40044
rect 3476 40004 7564 40032
rect 3476 39992 3482 40004
rect 7558 39992 7564 40004
rect 7616 39992 7622 40044
rect 7282 39788 7288 39840
rect 7340 39828 7346 39840
rect 7469 39831 7527 39837
rect 7469 39828 7481 39831
rect 7340 39800 7481 39828
rect 7340 39788 7346 39800
rect 7469 39797 7481 39800
rect 7515 39797 7527 39831
rect 7469 39791 7527 39797
rect 1104 39738 7912 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 7912 39738
rect 1104 39664 7912 39686
rect 104052 39738 108836 39760
rect 104052 39686 105922 39738
rect 105974 39686 105986 39738
rect 106038 39686 106050 39738
rect 106102 39686 106114 39738
rect 106166 39686 106178 39738
rect 106230 39686 108836 39738
rect 104052 39664 108836 39686
rect 1104 39194 7912 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 7912 39194
rect 1104 39120 7912 39142
rect 104052 39194 108836 39216
rect 104052 39142 106658 39194
rect 106710 39142 106722 39194
rect 106774 39142 106786 39194
rect 106838 39142 106850 39194
rect 106902 39142 106914 39194
rect 106966 39142 108836 39194
rect 104052 39120 108836 39142
rect 7558 38700 7564 38752
rect 7616 38700 7622 38752
rect 1104 38650 7912 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 7912 38650
rect 1104 38576 7912 38598
rect 104052 38650 108836 38672
rect 104052 38598 105922 38650
rect 105974 38598 105986 38650
rect 106038 38598 106050 38650
rect 106102 38598 106114 38650
rect 106166 38598 106178 38650
rect 106230 38598 108836 38650
rect 104052 38576 108836 38598
rect 1104 38106 7912 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 7912 38106
rect 1104 38032 7912 38054
rect 104052 38106 108836 38128
rect 104052 38054 106658 38106
rect 106710 38054 106722 38106
rect 106774 38054 106786 38106
rect 106838 38054 106850 38106
rect 106902 38054 106914 38106
rect 106966 38054 108836 38106
rect 104052 38032 108836 38054
rect 1104 37562 7912 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 7912 37562
rect 1104 37488 7912 37510
rect 104052 37562 108836 37584
rect 104052 37510 105922 37562
rect 105974 37510 105986 37562
rect 106038 37510 106050 37562
rect 106102 37510 106114 37562
rect 106166 37510 106178 37562
rect 106230 37510 108836 37562
rect 104052 37488 108836 37510
rect 1104 37018 7912 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 7912 37018
rect 1104 36944 7912 36966
rect 104052 37018 108836 37040
rect 104052 36966 106658 37018
rect 106710 36966 106722 37018
rect 106774 36966 106786 37018
rect 106838 36966 106850 37018
rect 106902 36966 106914 37018
rect 106966 36966 108836 37018
rect 104052 36944 108836 36966
rect 7558 36592 7564 36644
rect 7616 36592 7622 36644
rect 1104 36474 7912 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 7912 36474
rect 1104 36400 7912 36422
rect 104052 36474 108836 36496
rect 104052 36422 105922 36474
rect 105974 36422 105986 36474
rect 106038 36422 106050 36474
rect 106102 36422 106114 36474
rect 106166 36422 106178 36474
rect 106230 36422 108836 36474
rect 104052 36400 108836 36422
rect 1104 35930 7912 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 7912 35930
rect 1104 35856 7912 35878
rect 104052 35930 108836 35952
rect 104052 35878 106658 35930
rect 106710 35878 106722 35930
rect 106774 35878 106786 35930
rect 106838 35878 106850 35930
rect 106902 35878 106914 35930
rect 106966 35878 108836 35930
rect 104052 35856 108836 35878
rect 7466 35436 7472 35488
rect 7524 35436 7530 35488
rect 1104 35386 7912 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 7912 35386
rect 1104 35312 7912 35334
rect 104052 35386 108836 35408
rect 104052 35334 105922 35386
rect 105974 35334 105986 35386
rect 106038 35334 106050 35386
rect 106102 35334 106114 35386
rect 106166 35334 106178 35386
rect 106230 35334 108836 35386
rect 104052 35312 108836 35334
rect 1104 34842 7912 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 7912 34842
rect 1104 34768 7912 34790
rect 104052 34842 108836 34864
rect 104052 34790 106658 34842
rect 106710 34790 106722 34842
rect 106774 34790 106786 34842
rect 106838 34790 106850 34842
rect 106902 34790 106914 34842
rect 106966 34790 108836 34842
rect 104052 34768 108836 34790
rect 1104 34298 7912 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 7912 34298
rect 1104 34224 7912 34246
rect 104052 34298 108836 34320
rect 104052 34246 105922 34298
rect 105974 34246 105986 34298
rect 106038 34246 106050 34298
rect 106102 34246 106114 34298
rect 106166 34246 106178 34298
rect 106230 34246 108836 34298
rect 104052 34224 108836 34246
rect 7558 33872 7564 33924
rect 7616 33872 7622 33924
rect 1104 33754 7912 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 7912 33754
rect 1104 33680 7912 33702
rect 104052 33754 108836 33776
rect 104052 33702 106658 33754
rect 106710 33702 106722 33754
rect 106774 33702 106786 33754
rect 106838 33702 106850 33754
rect 106902 33702 106914 33754
rect 106966 33702 108836 33754
rect 104052 33680 108836 33702
rect 1104 33210 7912 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 7912 33210
rect 1104 33136 7912 33158
rect 104052 33210 108836 33232
rect 104052 33158 105922 33210
rect 105974 33158 105986 33210
rect 106038 33158 106050 33210
rect 106102 33158 106114 33210
rect 106166 33158 106178 33210
rect 106230 33158 108836 33210
rect 104052 33136 108836 33158
rect 1762 33056 1768 33108
rect 1820 33096 1826 33108
rect 7558 33096 7564 33108
rect 1820 33068 7564 33096
rect 1820 33056 1826 33068
rect 7558 33056 7564 33068
rect 7616 33056 7622 33108
rect 1104 32666 7912 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 7912 32666
rect 1104 32592 7912 32614
rect 104052 32666 108836 32688
rect 104052 32614 106658 32666
rect 106710 32614 106722 32666
rect 106774 32614 106786 32666
rect 106838 32614 106850 32666
rect 106902 32614 106914 32666
rect 106966 32614 108836 32666
rect 104052 32592 108836 32614
rect 1104 32122 7912 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 7912 32122
rect 1104 32048 7912 32070
rect 104052 32122 108836 32144
rect 104052 32070 105922 32122
rect 105974 32070 105986 32122
rect 106038 32070 106050 32122
rect 106102 32070 106114 32122
rect 106166 32070 106178 32122
rect 106230 32070 108836 32122
rect 104052 32048 108836 32070
rect 1104 31578 7912 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 7912 31578
rect 1104 31504 7912 31526
rect 104052 31578 108836 31600
rect 104052 31526 106658 31578
rect 106710 31526 106722 31578
rect 106774 31526 106786 31578
rect 106838 31526 106850 31578
rect 106902 31526 106914 31578
rect 106966 31526 108836 31578
rect 104052 31504 108836 31526
rect 1104 31034 7912 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 7912 31034
rect 1104 30960 7912 30982
rect 104052 31034 108836 31056
rect 104052 30982 105922 31034
rect 105974 30982 105986 31034
rect 106038 30982 106050 31034
rect 106102 30982 106114 31034
rect 106166 30982 106178 31034
rect 106230 30982 108836 31034
rect 104052 30960 108836 30982
rect 1104 30490 7912 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 7912 30490
rect 1104 30416 7912 30438
rect 104052 30490 108836 30512
rect 104052 30438 106658 30490
rect 106710 30438 106722 30490
rect 106774 30438 106786 30490
rect 106838 30438 106850 30490
rect 106902 30438 106914 30490
rect 106966 30438 108836 30490
rect 104052 30416 108836 30438
rect 1578 30268 1584 30320
rect 1636 30308 1642 30320
rect 7466 30308 7472 30320
rect 1636 30280 7472 30308
rect 1636 30268 1642 30280
rect 7466 30268 7472 30280
rect 7524 30268 7530 30320
rect 1104 29946 7912 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 7912 29946
rect 1104 29872 7912 29894
rect 104052 29946 108836 29968
rect 104052 29894 105922 29946
rect 105974 29894 105986 29946
rect 106038 29894 106050 29946
rect 106102 29894 106114 29946
rect 106166 29894 106178 29946
rect 106230 29894 108836 29946
rect 104052 29872 108836 29894
rect 1104 29402 7912 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 7912 29402
rect 1104 29328 7912 29350
rect 104052 29402 108836 29424
rect 104052 29350 106658 29402
rect 106710 29350 106722 29402
rect 106774 29350 106786 29402
rect 106838 29350 106850 29402
rect 106902 29350 106914 29402
rect 106966 29350 108836 29402
rect 104052 29328 108836 29350
rect 1104 28858 7912 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 7912 28858
rect 1104 28784 7912 28806
rect 104052 28858 108836 28880
rect 104052 28806 105922 28858
rect 105974 28806 105986 28858
rect 106038 28806 106050 28858
rect 106102 28806 106114 28858
rect 106166 28806 106178 28858
rect 106230 28806 108836 28858
rect 104052 28784 108836 28806
rect 1104 28314 7912 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 7912 28314
rect 1104 28240 7912 28262
rect 104052 28314 108836 28336
rect 104052 28262 106658 28314
rect 106710 28262 106722 28314
rect 106774 28262 106786 28314
rect 106838 28262 106850 28314
rect 106902 28262 106914 28314
rect 106966 28262 108836 28314
rect 104052 28240 108836 28262
rect 1104 27770 7912 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 7912 27770
rect 1104 27696 7912 27718
rect 104052 27770 108836 27792
rect 104052 27718 105922 27770
rect 105974 27718 105986 27770
rect 106038 27718 106050 27770
rect 106102 27718 106114 27770
rect 106166 27718 106178 27770
rect 106230 27718 108836 27770
rect 104052 27696 108836 27718
rect 1104 27226 7912 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 7912 27226
rect 1104 27152 7912 27174
rect 104052 27226 108836 27248
rect 104052 27174 106658 27226
rect 106710 27174 106722 27226
rect 106774 27174 106786 27226
rect 106838 27174 106850 27226
rect 106902 27174 106914 27226
rect 106966 27174 108836 27226
rect 104052 27152 108836 27174
rect 1104 26682 7912 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 7912 26682
rect 1104 26608 7912 26630
rect 104052 26682 108836 26704
rect 104052 26630 105922 26682
rect 105974 26630 105986 26682
rect 106038 26630 106050 26682
rect 106102 26630 106114 26682
rect 106166 26630 106178 26682
rect 106230 26630 108836 26682
rect 104052 26608 108836 26630
rect 1670 26256 1676 26308
rect 1728 26296 1734 26308
rect 7374 26296 7380 26308
rect 1728 26268 7380 26296
rect 1728 26256 1734 26268
rect 7374 26256 7380 26268
rect 7432 26256 7438 26308
rect 1104 26138 7912 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 7912 26138
rect 1104 26064 7912 26086
rect 104052 26138 108836 26160
rect 104052 26086 106658 26138
rect 106710 26086 106722 26138
rect 106774 26086 106786 26138
rect 106838 26086 106850 26138
rect 106902 26086 106914 26138
rect 106966 26086 108836 26138
rect 104052 26064 108836 26086
rect 1104 25594 7912 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 7912 25594
rect 1104 25520 7912 25542
rect 104052 25594 108836 25616
rect 104052 25542 105922 25594
rect 105974 25542 105986 25594
rect 106038 25542 106050 25594
rect 106102 25542 106114 25594
rect 106166 25542 106178 25594
rect 106230 25542 108836 25594
rect 104052 25520 108836 25542
rect 102594 25100 102600 25152
rect 102652 25140 102658 25152
rect 104345 25143 104403 25149
rect 104345 25140 104357 25143
rect 102652 25112 104357 25140
rect 102652 25100 102658 25112
rect 104345 25109 104357 25112
rect 104391 25109 104403 25143
rect 104345 25103 104403 25109
rect 1104 25050 7912 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 7912 25050
rect 1104 24976 7912 24998
rect 104052 25050 108836 25072
rect 104052 24998 106658 25050
rect 106710 24998 106722 25050
rect 106774 24998 106786 25050
rect 106838 24998 106850 25050
rect 106902 24998 106914 25050
rect 106966 24998 108836 25050
rect 104052 24976 108836 24998
rect 1104 24506 7912 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 7912 24506
rect 1104 24432 7912 24454
rect 104052 24506 108836 24528
rect 104052 24454 105922 24506
rect 105974 24454 105986 24506
rect 106038 24454 106050 24506
rect 106102 24454 106114 24506
rect 106166 24454 106178 24506
rect 106230 24454 108836 24506
rect 104052 24432 108836 24454
rect 1104 23962 7912 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 7912 23962
rect 1104 23888 7912 23910
rect 104052 23962 108836 23984
rect 104052 23910 106658 23962
rect 106710 23910 106722 23962
rect 106774 23910 106786 23962
rect 106838 23910 106850 23962
rect 106902 23910 106914 23962
rect 106966 23910 108836 23962
rect 104052 23888 108836 23910
rect 101950 23808 101956 23860
rect 102008 23848 102014 23860
rect 104345 23851 104403 23857
rect 104345 23848 104357 23851
rect 102008 23820 104357 23848
rect 102008 23808 102014 23820
rect 104345 23817 104357 23820
rect 104391 23817 104403 23851
rect 104345 23811 104403 23817
rect 1854 23604 1860 23656
rect 1912 23644 1918 23656
rect 7558 23644 7564 23656
rect 1912 23616 7564 23644
rect 1912 23604 1918 23616
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 1104 23418 7912 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 7912 23418
rect 1104 23344 7912 23366
rect 104052 23418 108836 23440
rect 104052 23366 105922 23418
rect 105974 23366 105986 23418
rect 106038 23366 106050 23418
rect 106102 23366 106114 23418
rect 106166 23366 106178 23418
rect 106230 23366 108836 23418
rect 104052 23344 108836 23366
rect 1104 22874 7912 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 7912 22874
rect 1104 22800 7912 22822
rect 104052 22874 108836 22896
rect 104052 22822 106658 22874
rect 106710 22822 106722 22874
rect 106774 22822 106786 22874
rect 106838 22822 106850 22874
rect 106902 22822 106914 22874
rect 106966 22822 108836 22874
rect 104052 22800 108836 22822
rect 102318 22720 102324 22772
rect 102376 22760 102382 22772
rect 104345 22763 104403 22769
rect 104345 22760 104357 22763
rect 102376 22732 104357 22760
rect 102376 22720 102382 22732
rect 104345 22729 104357 22732
rect 104391 22729 104403 22763
rect 104345 22723 104403 22729
rect 1104 22330 7912 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 7912 22330
rect 1104 22256 7912 22278
rect 104052 22330 108836 22352
rect 104052 22278 105922 22330
rect 105974 22278 105986 22330
rect 106038 22278 106050 22330
rect 106102 22278 106114 22330
rect 106166 22278 106178 22330
rect 106230 22278 108836 22330
rect 104052 22256 108836 22278
rect 1104 21786 7912 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 7912 21786
rect 1104 21712 7912 21734
rect 104052 21786 108836 21808
rect 104052 21734 106658 21786
rect 106710 21734 106722 21786
rect 106774 21734 106786 21786
rect 106838 21734 106850 21786
rect 106902 21734 106914 21786
rect 106966 21734 108836 21786
rect 104052 21712 108836 21734
rect 1104 21242 7912 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 7912 21242
rect 1104 21168 7912 21190
rect 104052 21242 108836 21264
rect 104052 21190 105922 21242
rect 105974 21190 105986 21242
rect 106038 21190 106050 21242
rect 106102 21190 106114 21242
rect 106166 21190 106178 21242
rect 106230 21190 108836 21242
rect 104052 21168 108836 21190
rect 1104 20698 7912 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 7912 20698
rect 1104 20624 7912 20646
rect 104052 20698 108836 20720
rect 104052 20646 106658 20698
rect 106710 20646 106722 20698
rect 106774 20646 106786 20698
rect 106838 20646 106850 20698
rect 106902 20646 106914 20698
rect 106966 20646 108836 20698
rect 104052 20624 108836 20646
rect 1104 20154 7912 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 7912 20154
rect 1104 20080 7912 20102
rect 104052 20154 108836 20176
rect 104052 20102 105922 20154
rect 105974 20102 105986 20154
rect 106038 20102 106050 20154
rect 106102 20102 106114 20154
rect 106166 20102 106178 20154
rect 106230 20102 108836 20154
rect 104052 20080 108836 20102
rect 1104 19610 7912 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 7912 19610
rect 1104 19536 7912 19558
rect 104052 19610 108836 19632
rect 104052 19558 106658 19610
rect 106710 19558 106722 19610
rect 106774 19558 106786 19610
rect 106838 19558 106850 19610
rect 106902 19558 106914 19610
rect 106966 19558 108836 19610
rect 104052 19536 108836 19558
rect 1104 19066 7912 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 7912 19066
rect 1104 18992 7912 19014
rect 104052 19066 108836 19088
rect 104052 19014 105922 19066
rect 105974 19014 105986 19066
rect 106038 19014 106050 19066
rect 106102 19014 106114 19066
rect 106166 19014 106178 19066
rect 106230 19014 108836 19066
rect 104052 18992 108836 19014
rect 1104 18522 7912 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 7912 18522
rect 1104 18448 7912 18470
rect 104052 18522 108836 18544
rect 104052 18470 106658 18522
rect 106710 18470 106722 18522
rect 106774 18470 106786 18522
rect 106838 18470 106850 18522
rect 106902 18470 106914 18522
rect 106966 18470 108836 18522
rect 104052 18448 108836 18470
rect 1104 17978 7912 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 7912 17978
rect 1104 17904 7912 17926
rect 104052 17978 108836 18000
rect 104052 17926 105922 17978
rect 105974 17926 105986 17978
rect 106038 17926 106050 17978
rect 106102 17926 106114 17978
rect 106166 17926 106178 17978
rect 106230 17926 108836 17978
rect 104052 17904 108836 17926
rect 1104 17434 7912 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 7912 17434
rect 1104 17360 7912 17382
rect 104052 17434 108836 17456
rect 104052 17382 106658 17434
rect 106710 17382 106722 17434
rect 106774 17382 106786 17434
rect 106838 17382 106850 17434
rect 106902 17382 106914 17434
rect 106966 17382 108836 17434
rect 104052 17360 108836 17382
rect 1104 16890 7912 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 7912 16890
rect 1104 16816 7912 16838
rect 104052 16890 108836 16912
rect 104052 16838 105922 16890
rect 105974 16838 105986 16890
rect 106038 16838 106050 16890
rect 106102 16838 106114 16890
rect 106166 16838 106178 16890
rect 106230 16838 108836 16890
rect 104052 16816 108836 16838
rect 1104 16346 7912 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 7912 16346
rect 1104 16272 7912 16294
rect 104052 16346 108836 16368
rect 104052 16294 106658 16346
rect 106710 16294 106722 16346
rect 106774 16294 106786 16346
rect 106838 16294 106850 16346
rect 106902 16294 106914 16346
rect 106966 16294 108836 16346
rect 104052 16272 108836 16294
rect 1104 15802 7912 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 7912 15802
rect 1104 15728 7912 15750
rect 104052 15802 108836 15824
rect 104052 15750 105922 15802
rect 105974 15750 105986 15802
rect 106038 15750 106050 15802
rect 106102 15750 106114 15802
rect 106166 15750 106178 15802
rect 106230 15750 108836 15802
rect 104052 15728 108836 15750
rect 7466 15308 7472 15360
rect 7524 15308 7530 15360
rect 1104 15258 7912 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 7912 15258
rect 1104 15184 7912 15206
rect 104052 15258 108836 15280
rect 104052 15206 106658 15258
rect 106710 15206 106722 15258
rect 106774 15206 106786 15258
rect 106838 15206 106850 15258
rect 106902 15206 106914 15258
rect 106966 15206 108836 15258
rect 104052 15184 108836 15206
rect 1104 14714 7912 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 7912 14714
rect 1104 14640 7912 14662
rect 104052 14714 108836 14736
rect 104052 14662 105922 14714
rect 105974 14662 105986 14714
rect 106038 14662 106050 14714
rect 106102 14662 106114 14714
rect 106166 14662 106178 14714
rect 106230 14662 108836 14714
rect 104052 14640 108836 14662
rect 1104 14170 7912 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 7912 14170
rect 1104 14096 7912 14118
rect 104052 14170 108836 14192
rect 104052 14118 106658 14170
rect 106710 14118 106722 14170
rect 106774 14118 106786 14170
rect 106838 14118 106850 14170
rect 106902 14118 106914 14170
rect 106966 14118 108836 14170
rect 104052 14096 108836 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1857 14059 1915 14065
rect 1857 14056 1869 14059
rect 1627 14028 1869 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1857 14025 1869 14028
rect 1903 14056 1915 14059
rect 3418 14056 3424 14068
rect 1903 14028 3424 14056
rect 1903 14025 1915 14028
rect 1857 14019 1915 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1949 13923 2007 13929
rect 1949 13920 1961 13923
rect 1544 13892 1961 13920
rect 1544 13880 1550 13892
rect 1949 13889 1961 13892
rect 1995 13889 2007 13923
rect 1949 13883 2007 13889
rect 1104 13626 7912 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 7912 13626
rect 1104 13552 7912 13574
rect 104052 13626 108836 13648
rect 104052 13574 105922 13626
rect 105974 13574 105986 13626
rect 106038 13574 106050 13626
rect 106102 13574 106114 13626
rect 106166 13574 106178 13626
rect 106230 13574 108836 13626
rect 104052 13552 108836 13574
rect 1581 13515 1639 13521
rect 1581 13481 1593 13515
rect 1627 13512 1639 13515
rect 1854 13512 1860 13524
rect 1627 13484 1860 13512
rect 1627 13481 1639 13484
rect 1581 13475 1639 13481
rect 1854 13472 1860 13484
rect 1912 13472 1918 13524
rect 1302 13200 1308 13252
rect 1360 13240 1366 13252
rect 1489 13243 1547 13249
rect 1489 13240 1501 13243
rect 1360 13212 1501 13240
rect 1360 13200 1366 13212
rect 1489 13209 1501 13212
rect 1535 13240 1547 13243
rect 1949 13243 2007 13249
rect 1949 13240 1961 13243
rect 1535 13212 1961 13240
rect 1535 13209 1547 13212
rect 1489 13203 1547 13209
rect 1949 13209 1961 13212
rect 1995 13209 2007 13243
rect 1949 13203 2007 13209
rect 1104 13082 7912 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 7912 13082
rect 1104 13008 7912 13030
rect 104052 13082 108836 13104
rect 104052 13030 106658 13082
rect 106710 13030 106722 13082
rect 106774 13030 106786 13082
rect 106838 13030 106850 13082
rect 106902 13030 106914 13082
rect 106966 13030 108836 13082
rect 104052 13008 108836 13030
rect 1670 12860 1676 12912
rect 1728 12900 1734 12912
rect 1765 12903 1823 12909
rect 1765 12900 1777 12903
rect 1728 12872 1777 12900
rect 1728 12860 1734 12872
rect 1765 12869 1777 12872
rect 1811 12869 1823 12903
rect 1765 12863 1823 12869
rect 1486 12792 1492 12844
rect 1544 12832 1550 12844
rect 1949 12835 2007 12841
rect 1949 12832 1961 12835
rect 1544 12804 1961 12832
rect 1544 12792 1550 12804
rect 1949 12801 1961 12804
rect 1995 12801 2007 12835
rect 1949 12795 2007 12801
rect 1104 12538 7912 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 7912 12538
rect 1104 12464 7912 12486
rect 104052 12538 108836 12560
rect 104052 12486 105922 12538
rect 105974 12486 105986 12538
rect 106038 12486 106050 12538
rect 106102 12486 106114 12538
rect 106166 12486 106178 12538
rect 106230 12486 108836 12538
rect 104052 12464 108836 12486
rect 1104 11994 7912 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 7912 11994
rect 1104 11920 7912 11942
rect 104052 11994 108836 12016
rect 104052 11942 106658 11994
rect 106710 11942 106722 11994
rect 106774 11942 106786 11994
rect 106838 11942 106850 11994
rect 106902 11942 106914 11994
rect 106966 11942 108836 11994
rect 104052 11920 108836 11942
rect 1578 11840 1584 11892
rect 1636 11880 1642 11892
rect 1765 11883 1823 11889
rect 1765 11880 1777 11883
rect 1636 11852 1777 11880
rect 1636 11840 1642 11852
rect 1765 11849 1777 11852
rect 1811 11849 1823 11883
rect 1765 11843 1823 11849
rect 1210 11704 1216 11756
rect 1268 11744 1274 11756
rect 1489 11747 1547 11753
rect 1489 11744 1501 11747
rect 1268 11716 1501 11744
rect 1268 11704 1274 11716
rect 1489 11713 1501 11716
rect 1535 11744 1547 11747
rect 1949 11747 2007 11753
rect 1949 11744 1961 11747
rect 1535 11716 1961 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1949 11713 1961 11716
rect 1995 11713 2007 11747
rect 1949 11707 2007 11713
rect 1104 11450 7912 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 7912 11450
rect 1104 11376 7912 11398
rect 104052 11450 108836 11472
rect 104052 11398 105922 11450
rect 105974 11398 105986 11450
rect 106038 11398 106050 11450
rect 106102 11398 106114 11450
rect 106166 11398 106178 11450
rect 106230 11398 108836 11450
rect 104052 11376 108836 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 1857 11339 1915 11345
rect 1857 11336 1869 11339
rect 1627 11308 1869 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 1857 11305 1869 11308
rect 1903 11336 1915 11339
rect 7282 11336 7288 11348
rect 1903 11308 7288 11336
rect 1903 11305 1915 11308
rect 1857 11299 1915 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 1486 11024 1492 11076
rect 1544 11064 1550 11076
rect 1949 11067 2007 11073
rect 1949 11064 1961 11067
rect 1544 11036 1961 11064
rect 1544 11024 1550 11036
rect 1949 11033 1961 11036
rect 1995 11033 2007 11067
rect 1949 11027 2007 11033
rect 1104 10906 7912 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 7912 10906
rect 1104 10832 7912 10854
rect 104052 10906 108836 10928
rect 104052 10854 106658 10906
rect 106710 10854 106722 10906
rect 106774 10854 106786 10906
rect 106838 10854 106850 10906
rect 106902 10854 106914 10906
rect 106966 10854 108836 10906
rect 104052 10832 108836 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 1762 10792 1768 10804
rect 1627 10764 1768 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 1489 10659 1547 10665
rect 1489 10656 1501 10659
rect 1360 10628 1501 10656
rect 1360 10616 1366 10628
rect 1489 10625 1501 10628
rect 1535 10656 1547 10659
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1535 10628 1961 10656
rect 1535 10625 1547 10628
rect 1489 10619 1547 10625
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 1949 10619 2007 10625
rect 1104 10362 7912 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 7912 10362
rect 1104 10288 7912 10310
rect 104052 10362 108836 10384
rect 104052 10310 105922 10362
rect 105974 10310 105986 10362
rect 106038 10310 106050 10362
rect 106102 10310 106114 10362
rect 106166 10310 106178 10362
rect 106230 10310 108836 10362
rect 104052 10288 108836 10310
rect 1486 9936 1492 9988
rect 1544 9936 1550 9988
rect 1673 9979 1731 9985
rect 1673 9945 1685 9979
rect 1719 9976 1731 9979
rect 1857 9979 1915 9985
rect 1857 9976 1869 9979
rect 1719 9948 1869 9976
rect 1719 9945 1731 9948
rect 1673 9939 1731 9945
rect 1857 9945 1869 9948
rect 1903 9976 1915 9979
rect 1903 9948 6914 9976
rect 1903 9945 1915 9948
rect 1857 9939 1915 9945
rect 1504 9908 1532 9936
rect 1949 9911 2007 9917
rect 1949 9908 1961 9911
rect 1504 9880 1961 9908
rect 1949 9877 1961 9880
rect 1995 9877 2007 9911
rect 6886 9908 6914 9948
rect 29546 9908 29552 9920
rect 6886 9880 29552 9908
rect 1949 9871 2007 9877
rect 29546 9868 29552 9880
rect 29604 9868 29610 9920
rect 1104 9818 7912 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 7912 9818
rect 1104 9744 7912 9766
rect 104052 9818 108836 9840
rect 104052 9766 106658 9818
rect 106710 9766 106722 9818
rect 106774 9766 106786 9818
rect 106838 9766 106850 9818
rect 106902 9766 106914 9818
rect 106966 9766 108836 9818
rect 104052 9744 108836 9766
rect 9582 9596 9588 9648
rect 9640 9636 9646 9648
rect 16114 9636 16120 9648
rect 9640 9608 16120 9636
rect 9640 9596 9646 9608
rect 16114 9596 16120 9608
rect 16172 9596 16178 9648
rect 90542 9596 90548 9648
rect 90600 9636 90606 9648
rect 103606 9636 103612 9648
rect 90600 9608 103612 9636
rect 90600 9596 90606 9608
rect 103606 9596 103612 9608
rect 103664 9596 103670 9648
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 16022 9568 16028 9580
rect 6972 9540 16028 9568
rect 6972 9528 6978 9540
rect 16022 9528 16028 9540
rect 16080 9528 16086 9580
rect 90910 9528 90916 9580
rect 90968 9568 90974 9580
rect 103514 9568 103520 9580
rect 90968 9540 103520 9568
rect 90968 9528 90974 9540
rect 103514 9528 103520 9540
rect 103572 9528 103578 9580
rect 90726 9460 90732 9512
rect 90784 9500 90790 9512
rect 102134 9500 102140 9512
rect 90784 9472 102140 9500
rect 90784 9460 90790 9472
rect 102134 9460 102140 9472
rect 102192 9460 102198 9512
rect 1104 9274 7912 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 7912 9274
rect 1104 9200 7912 9222
rect 104052 9274 108836 9296
rect 104052 9222 105922 9274
rect 105974 9222 105986 9274
rect 106038 9222 106050 9274
rect 106102 9222 106114 9274
rect 106166 9222 106178 9274
rect 106230 9222 108836 9274
rect 104052 9200 108836 9222
rect 1302 8848 1308 8900
rect 1360 8888 1366 8900
rect 1489 8891 1547 8897
rect 1489 8888 1501 8891
rect 1360 8860 1501 8888
rect 1360 8848 1366 8860
rect 1489 8857 1501 8860
rect 1535 8857 1547 8891
rect 1489 8851 1547 8857
rect 1673 8891 1731 8897
rect 1673 8857 1685 8891
rect 1719 8888 1731 8891
rect 1857 8891 1915 8897
rect 1857 8888 1869 8891
rect 1719 8860 1869 8888
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 1857 8857 1869 8860
rect 1903 8888 1915 8891
rect 1903 8860 6914 8888
rect 1903 8857 1915 8860
rect 1857 8851 1915 8857
rect 1504 8820 1532 8851
rect 1949 8823 2007 8829
rect 1949 8820 1961 8823
rect 1504 8792 1961 8820
rect 1949 8789 1961 8792
rect 1995 8789 2007 8823
rect 6886 8820 6914 8860
rect 26694 8820 26700 8832
rect 6886 8792 26700 8820
rect 1949 8783 2007 8789
rect 26694 8780 26700 8792
rect 26752 8780 26758 8832
rect 1104 8730 7912 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 7912 8730
rect 1104 8656 7912 8678
rect 104052 8730 108836 8752
rect 104052 8678 106658 8730
rect 106710 8678 106722 8730
rect 106774 8678 106786 8730
rect 106838 8678 106850 8730
rect 106902 8678 106914 8730
rect 106966 8678 108836 8730
rect 104052 8656 108836 8678
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8381 2007 8415
rect 1949 8375 2007 8381
rect 1964 8344 1992 8375
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 2096 8384 2237 8412
rect 2096 8372 2102 8384
rect 2225 8381 2237 8384
rect 2271 8381 2283 8415
rect 2225 8375 2283 8381
rect 2409 8347 2467 8353
rect 2409 8344 2421 8347
rect 1964 8316 2421 8344
rect 2409 8313 2421 8316
rect 2455 8344 2467 8347
rect 24670 8344 24676 8356
rect 2455 8316 24676 8344
rect 2455 8313 2467 8316
rect 2409 8307 2467 8313
rect 24670 8304 24676 8316
rect 24728 8304 24734 8356
rect 1104 8186 7912 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 7912 8186
rect 1104 8112 7912 8134
rect 104052 8186 108836 8208
rect 104052 8134 105922 8186
rect 105974 8134 105986 8186
rect 106038 8134 106050 8186
rect 106102 8134 106114 8186
rect 106166 8134 106178 8186
rect 106230 8134 108836 8186
rect 104052 8112 108836 8134
rect 1946 8032 1952 8084
rect 2004 8032 2010 8084
rect 2133 7871 2191 7877
rect 2133 7868 2145 7871
rect 1504 7840 2145 7868
rect 1302 7760 1308 7812
rect 1360 7800 1366 7812
rect 1504 7809 1532 7840
rect 2133 7837 2145 7840
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 1489 7803 1547 7809
rect 1489 7800 1501 7803
rect 1360 7772 1501 7800
rect 1360 7760 1366 7772
rect 1489 7769 1501 7772
rect 1535 7769 1547 7803
rect 1489 7763 1547 7769
rect 1673 7803 1731 7809
rect 1673 7769 1685 7803
rect 1719 7800 1731 7803
rect 1857 7803 1915 7809
rect 1857 7800 1869 7803
rect 1719 7772 1869 7800
rect 1719 7769 1731 7772
rect 1673 7763 1731 7769
rect 1857 7769 1869 7772
rect 1903 7800 1915 7803
rect 1903 7772 6914 7800
rect 1903 7769 1915 7772
rect 1857 7763 1915 7769
rect 6886 7732 6914 7772
rect 30466 7732 30472 7744
rect 6886 7704 30472 7732
rect 30466 7692 30472 7704
rect 30524 7692 30530 7744
rect 1104 7642 108836 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 66314 7642
rect 66366 7590 66378 7642
rect 66430 7590 66442 7642
rect 66494 7590 66506 7642
rect 66558 7590 66570 7642
rect 66622 7590 97034 7642
rect 97086 7590 97098 7642
rect 97150 7590 97162 7642
rect 97214 7590 97226 7642
rect 97278 7590 97290 7642
rect 97342 7590 106658 7642
rect 106710 7590 106722 7642
rect 106774 7590 106786 7642
rect 106838 7590 106850 7642
rect 106902 7590 106914 7642
rect 106966 7590 108836 7642
rect 1104 7568 108836 7590
rect 16022 7488 16028 7540
rect 16080 7528 16086 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 16080 7500 16129 7528
rect 16080 7488 16086 7500
rect 16117 7497 16129 7500
rect 16163 7497 16175 7531
rect 16117 7491 16175 7497
rect 23474 7488 23480 7540
rect 23532 7488 23538 7540
rect 24670 7488 24676 7540
rect 24728 7488 24734 7540
rect 25774 7488 25780 7540
rect 25832 7528 25838 7540
rect 25869 7531 25927 7537
rect 25869 7528 25881 7531
rect 25832 7500 25881 7528
rect 25832 7488 25838 7500
rect 25869 7497 25881 7500
rect 25915 7497 25927 7531
rect 25869 7491 25927 7497
rect 26694 7488 26700 7540
rect 26752 7528 26758 7540
rect 26973 7531 27031 7537
rect 26973 7528 26985 7531
rect 26752 7500 26985 7528
rect 26752 7488 26758 7500
rect 26973 7497 26985 7500
rect 27019 7497 27031 7531
rect 26973 7491 27031 7497
rect 28166 7488 28172 7540
rect 28224 7488 28230 7540
rect 29546 7488 29552 7540
rect 29604 7488 29610 7540
rect 30466 7488 30472 7540
rect 30524 7488 30530 7540
rect 90542 7488 90548 7540
rect 90600 7488 90606 7540
rect 90726 7488 90732 7540
rect 90784 7488 90790 7540
rect 90910 7488 90916 7540
rect 90968 7488 90974 7540
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1489 7395 1547 7401
rect 1489 7392 1501 7395
rect 1360 7364 1501 7392
rect 1360 7352 1366 7364
rect 1489 7361 1501 7364
rect 1535 7392 1547 7395
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1535 7364 1961 7392
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 1857 7259 1915 7265
rect 1857 7256 1869 7259
rect 1719 7228 1869 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 1857 7225 1869 7228
rect 1903 7256 1915 7259
rect 28166 7256 28172 7268
rect 1903 7228 28172 7256
rect 1903 7225 1915 7228
rect 1857 7219 1915 7225
rect 28166 7216 28172 7228
rect 28224 7216 28230 7268
rect 1104 7098 108836 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 96374 7098
rect 96426 7046 96438 7098
rect 96490 7046 96502 7098
rect 96554 7046 96566 7098
rect 96618 7046 96630 7098
rect 96682 7046 105922 7098
rect 105974 7046 105986 7098
rect 106038 7046 106050 7098
rect 106102 7046 106114 7098
rect 106166 7046 106178 7098
rect 106230 7046 108836 7098
rect 1104 7024 108836 7046
rect 1104 6554 108836 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 66314 6554
rect 66366 6502 66378 6554
rect 66430 6502 66442 6554
rect 66494 6502 66506 6554
rect 66558 6502 66570 6554
rect 66622 6502 97034 6554
rect 97086 6502 97098 6554
rect 97150 6502 97162 6554
rect 97214 6502 97226 6554
rect 97278 6502 97290 6554
rect 97342 6502 108836 6554
rect 1104 6480 108836 6502
rect 1210 6264 1216 6316
rect 1268 6304 1274 6316
rect 1489 6307 1547 6313
rect 1489 6304 1501 6307
rect 1268 6276 1501 6304
rect 1268 6264 1274 6276
rect 1489 6273 1501 6276
rect 1535 6304 1547 6307
rect 1949 6307 2007 6313
rect 1949 6304 1961 6307
rect 1535 6276 1961 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 1949 6273 1961 6276
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 1673 6171 1731 6177
rect 1673 6137 1685 6171
rect 1719 6168 1731 6171
rect 1857 6171 1915 6177
rect 1857 6168 1869 6171
rect 1719 6140 1869 6168
rect 1719 6137 1731 6140
rect 1673 6131 1731 6137
rect 1857 6137 1869 6140
rect 1903 6168 1915 6171
rect 1903 6140 6914 6168
rect 1903 6137 1915 6140
rect 1857 6131 1915 6137
rect 6886 6100 6914 6140
rect 25866 6100 25872 6112
rect 6886 6072 25872 6100
rect 25866 6060 25872 6072
rect 25924 6060 25930 6112
rect 1104 6010 108836 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 96374 6010
rect 96426 5958 96438 6010
rect 96490 5958 96502 6010
rect 96554 5958 96566 6010
rect 96618 5958 96630 6010
rect 96682 5958 108836 6010
rect 1104 5936 108836 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1765 5899 1823 5905
rect 1765 5896 1777 5899
rect 1627 5868 1777 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 1765 5865 1777 5868
rect 1811 5896 1823 5899
rect 7466 5896 7472 5908
rect 1811 5868 7472 5896
rect 1811 5865 1823 5868
rect 1765 5859 1823 5865
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 1394 5652 1400 5704
rect 1452 5692 1458 5704
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1452 5664 1869 5692
rect 1452 5652 1458 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 1104 5466 108836 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 66314 5466
rect 66366 5414 66378 5466
rect 66430 5414 66442 5466
rect 66494 5414 66506 5466
rect 66558 5414 66570 5466
rect 66622 5414 97034 5466
rect 97086 5414 97098 5466
rect 97150 5414 97162 5466
rect 97214 5414 97226 5466
rect 97278 5414 97290 5466
rect 97342 5414 108836 5466
rect 1104 5392 108836 5414
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1489 5219 1547 5225
rect 1489 5216 1501 5219
rect 1360 5188 1501 5216
rect 1360 5176 1366 5188
rect 1489 5185 1501 5188
rect 1535 5216 1547 5219
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1535 5188 1961 5216
rect 1535 5185 1547 5188
rect 1489 5179 1547 5185
rect 1949 5185 1961 5188
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 1673 5083 1731 5089
rect 1673 5049 1685 5083
rect 1719 5080 1731 5083
rect 1857 5083 1915 5089
rect 1857 5080 1869 5083
rect 1719 5052 1869 5080
rect 1719 5049 1731 5052
rect 1673 5043 1731 5049
rect 1857 5049 1869 5052
rect 1903 5080 1915 5083
rect 1903 5052 6914 5080
rect 1903 5049 1915 5052
rect 1857 5043 1915 5049
rect 6886 5012 6914 5052
rect 23474 5012 23480 5024
rect 6886 4984 23480 5012
rect 23474 4972 23480 4984
rect 23532 4972 23538 5024
rect 1104 4922 108836 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 96374 4922
rect 96426 4870 96438 4922
rect 96490 4870 96502 4922
rect 96554 4870 96566 4922
rect 96618 4870 96630 4922
rect 96682 4870 108836 4922
rect 1104 4848 108836 4870
rect 1104 4378 108836 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 66314 4378
rect 66366 4326 66378 4378
rect 66430 4326 66442 4378
rect 66494 4326 66506 4378
rect 66558 4326 66570 4378
rect 66622 4326 97034 4378
rect 97086 4326 97098 4378
rect 97150 4326 97162 4378
rect 97214 4326 97226 4378
rect 97278 4326 97290 4378
rect 97342 4326 108836 4378
rect 1104 4304 108836 4326
rect 1104 3834 108836 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 96374 3834
rect 96426 3782 96438 3834
rect 96490 3782 96502 3834
rect 96554 3782 96566 3834
rect 96618 3782 96630 3834
rect 96682 3782 108836 3834
rect 1104 3760 108836 3782
rect 1104 3290 108836 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 66314 3290
rect 66366 3238 66378 3290
rect 66430 3238 66442 3290
rect 66494 3238 66506 3290
rect 66558 3238 66570 3290
rect 66622 3238 97034 3290
rect 97086 3238 97098 3290
rect 97150 3238 97162 3290
rect 97214 3238 97226 3290
rect 97278 3238 97290 3290
rect 97342 3238 108836 3290
rect 1104 3216 108836 3238
rect 1104 2746 108836 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 96374 2746
rect 96426 2694 96438 2746
rect 96490 2694 96502 2746
rect 96554 2694 96566 2746
rect 96618 2694 96630 2746
rect 96682 2694 108836 2746
rect 1104 2672 108836 2694
rect 31662 2592 31668 2644
rect 31720 2592 31726 2644
rect 32950 2592 32956 2644
rect 33008 2592 33014 2644
rect 34238 2592 34244 2644
rect 34296 2592 34302 2644
rect 35434 2592 35440 2644
rect 35492 2632 35498 2644
rect 35529 2635 35587 2641
rect 35529 2632 35541 2635
rect 35492 2604 35541 2632
rect 35492 2592 35498 2604
rect 35529 2601 35541 2604
rect 35575 2601 35587 2635
rect 35529 2595 35587 2601
rect 36354 2592 36360 2644
rect 36412 2592 36418 2644
rect 37458 2592 37464 2644
rect 37516 2592 37522 2644
rect 38746 2592 38752 2644
rect 38804 2592 38810 2644
rect 39942 2592 39948 2644
rect 40000 2632 40006 2644
rect 40037 2635 40095 2641
rect 40037 2632 40049 2635
rect 40000 2604 40049 2632
rect 40000 2592 40006 2604
rect 40037 2601 40049 2604
rect 40083 2601 40095 2635
rect 40037 2595 40095 2601
rect 41322 2592 41328 2644
rect 41380 2592 41386 2644
rect 42150 2592 42156 2644
rect 42208 2592 42214 2644
rect 43438 2592 43444 2644
rect 43496 2592 43502 2644
rect 31849 2431 31907 2437
rect 31849 2428 31861 2431
rect 31588 2400 31861 2428
rect 31588 2304 31616 2400
rect 31849 2397 31861 2400
rect 31895 2397 31907 2431
rect 33137 2431 33195 2437
rect 33137 2428 33149 2431
rect 31849 2391 31907 2397
rect 32876 2400 33149 2428
rect 32876 2304 32904 2400
rect 33137 2397 33149 2400
rect 33183 2397 33195 2431
rect 34425 2431 34483 2437
rect 34425 2428 34437 2431
rect 33137 2391 33195 2397
rect 34164 2400 34437 2428
rect 34164 2304 34192 2400
rect 34425 2397 34437 2400
rect 34471 2397 34483 2431
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 34425 2391 34483 2397
rect 35452 2400 35725 2428
rect 35452 2304 35480 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 35713 2391 35771 2397
rect 36096 2400 36185 2428
rect 36096 2304 36124 2400
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 37645 2431 37703 2437
rect 37645 2428 37657 2431
rect 36173 2391 36231 2397
rect 37384 2400 37657 2428
rect 37384 2304 37412 2400
rect 37645 2397 37657 2400
rect 37691 2397 37703 2431
rect 38933 2431 38991 2437
rect 38933 2428 38945 2431
rect 37645 2391 37703 2397
rect 38672 2400 38945 2428
rect 38672 2304 38700 2400
rect 38933 2397 38945 2400
rect 38979 2397 38991 2431
rect 40221 2431 40279 2437
rect 40221 2428 40233 2431
rect 38933 2391 38991 2397
rect 39960 2400 40233 2428
rect 39960 2304 39988 2400
rect 40221 2397 40233 2400
rect 40267 2397 40279 2431
rect 41509 2431 41567 2437
rect 41509 2428 41521 2431
rect 40221 2391 40279 2397
rect 41248 2400 41521 2428
rect 41248 2304 41276 2400
rect 41509 2397 41521 2400
rect 41555 2397 41567 2431
rect 41969 2431 42027 2437
rect 41969 2428 41981 2431
rect 41509 2391 41567 2397
rect 41892 2400 41981 2428
rect 41892 2304 41920 2400
rect 41969 2397 41981 2400
rect 42015 2397 42027 2431
rect 43257 2431 43315 2437
rect 43257 2428 43269 2431
rect 41969 2391 42027 2397
rect 43180 2400 43269 2428
rect 43180 2304 43208 2400
rect 43257 2397 43269 2400
rect 43303 2397 43315 2431
rect 43257 2391 43315 2397
rect 31570 2252 31576 2304
rect 31628 2252 31634 2304
rect 32858 2252 32864 2304
rect 32916 2252 32922 2304
rect 34146 2252 34152 2304
rect 34204 2252 34210 2304
rect 35434 2252 35440 2304
rect 35492 2252 35498 2304
rect 36078 2252 36084 2304
rect 36136 2252 36142 2304
rect 37366 2252 37372 2304
rect 37424 2252 37430 2304
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 39942 2252 39948 2304
rect 40000 2252 40006 2304
rect 41230 2252 41236 2304
rect 41288 2252 41294 2304
rect 41874 2252 41880 2304
rect 41932 2252 41938 2304
rect 43162 2252 43168 2304
rect 43220 2252 43226 2304
rect 1104 2202 108836 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 66314 2202
rect 66366 2150 66378 2202
rect 66430 2150 66442 2202
rect 66494 2150 66506 2202
rect 66558 2150 66570 2202
rect 66622 2150 97034 2202
rect 97086 2150 97098 2202
rect 97150 2150 97162 2202
rect 97214 2150 97226 2202
rect 97278 2150 97290 2202
rect 97342 2150 108836 2202
rect 1104 2128 108836 2150
<< via1 >>
rect 4214 147398 4266 147450
rect 4278 147398 4330 147450
rect 4342 147398 4394 147450
rect 4406 147398 4458 147450
rect 4470 147398 4522 147450
rect 34934 147398 34986 147450
rect 34998 147398 35050 147450
rect 35062 147398 35114 147450
rect 35126 147398 35178 147450
rect 35190 147398 35242 147450
rect 65654 147398 65706 147450
rect 65718 147398 65770 147450
rect 65782 147398 65834 147450
rect 65846 147398 65898 147450
rect 65910 147398 65962 147450
rect 96374 147398 96426 147450
rect 96438 147398 96490 147450
rect 96502 147398 96554 147450
rect 96566 147398 96618 147450
rect 96630 147398 96682 147450
rect 4874 146854 4926 146906
rect 4938 146854 4990 146906
rect 5002 146854 5054 146906
rect 5066 146854 5118 146906
rect 5130 146854 5182 146906
rect 35594 146854 35646 146906
rect 35658 146854 35710 146906
rect 35722 146854 35774 146906
rect 35786 146854 35838 146906
rect 35850 146854 35902 146906
rect 66314 146854 66366 146906
rect 66378 146854 66430 146906
rect 66442 146854 66494 146906
rect 66506 146854 66558 146906
rect 66570 146854 66622 146906
rect 97034 146854 97086 146906
rect 97098 146854 97150 146906
rect 97162 146854 97214 146906
rect 97226 146854 97278 146906
rect 97290 146854 97342 146906
rect 4214 146310 4266 146362
rect 4278 146310 4330 146362
rect 4342 146310 4394 146362
rect 4406 146310 4458 146362
rect 4470 146310 4522 146362
rect 34934 146310 34986 146362
rect 34998 146310 35050 146362
rect 35062 146310 35114 146362
rect 35126 146310 35178 146362
rect 35190 146310 35242 146362
rect 65654 146310 65706 146362
rect 65718 146310 65770 146362
rect 65782 146310 65834 146362
rect 65846 146310 65898 146362
rect 65910 146310 65962 146362
rect 96374 146310 96426 146362
rect 96438 146310 96490 146362
rect 96502 146310 96554 146362
rect 96566 146310 96618 146362
rect 96630 146310 96682 146362
rect 4874 145766 4926 145818
rect 4938 145766 4990 145818
rect 5002 145766 5054 145818
rect 5066 145766 5118 145818
rect 5130 145766 5182 145818
rect 35594 145766 35646 145818
rect 35658 145766 35710 145818
rect 35722 145766 35774 145818
rect 35786 145766 35838 145818
rect 35850 145766 35902 145818
rect 66314 145766 66366 145818
rect 66378 145766 66430 145818
rect 66442 145766 66494 145818
rect 66506 145766 66558 145818
rect 66570 145766 66622 145818
rect 97034 145766 97086 145818
rect 97098 145766 97150 145818
rect 97162 145766 97214 145818
rect 97226 145766 97278 145818
rect 97290 145766 97342 145818
rect 4214 145222 4266 145274
rect 4278 145222 4330 145274
rect 4342 145222 4394 145274
rect 4406 145222 4458 145274
rect 4470 145222 4522 145274
rect 34934 145222 34986 145274
rect 34998 145222 35050 145274
rect 35062 145222 35114 145274
rect 35126 145222 35178 145274
rect 35190 145222 35242 145274
rect 65654 145222 65706 145274
rect 65718 145222 65770 145274
rect 65782 145222 65834 145274
rect 65846 145222 65898 145274
rect 65910 145222 65962 145274
rect 96374 145222 96426 145274
rect 96438 145222 96490 145274
rect 96502 145222 96554 145274
rect 96566 145222 96618 145274
rect 96630 145222 96682 145274
rect 4874 144678 4926 144730
rect 4938 144678 4990 144730
rect 5002 144678 5054 144730
rect 5066 144678 5118 144730
rect 5130 144678 5182 144730
rect 35594 144678 35646 144730
rect 35658 144678 35710 144730
rect 35722 144678 35774 144730
rect 35786 144678 35838 144730
rect 35850 144678 35902 144730
rect 66314 144678 66366 144730
rect 66378 144678 66430 144730
rect 66442 144678 66494 144730
rect 66506 144678 66558 144730
rect 66570 144678 66622 144730
rect 97034 144678 97086 144730
rect 97098 144678 97150 144730
rect 97162 144678 97214 144730
rect 97226 144678 97278 144730
rect 97290 144678 97342 144730
rect 4214 144134 4266 144186
rect 4278 144134 4330 144186
rect 4342 144134 4394 144186
rect 4406 144134 4458 144186
rect 4470 144134 4522 144186
rect 34934 144134 34986 144186
rect 34998 144134 35050 144186
rect 35062 144134 35114 144186
rect 35126 144134 35178 144186
rect 35190 144134 35242 144186
rect 65654 144134 65706 144186
rect 65718 144134 65770 144186
rect 65782 144134 65834 144186
rect 65846 144134 65898 144186
rect 65910 144134 65962 144186
rect 96374 144134 96426 144186
rect 96438 144134 96490 144186
rect 96502 144134 96554 144186
rect 96566 144134 96618 144186
rect 96630 144134 96682 144186
rect 4874 143590 4926 143642
rect 4938 143590 4990 143642
rect 5002 143590 5054 143642
rect 5066 143590 5118 143642
rect 5130 143590 5182 143642
rect 35594 143590 35646 143642
rect 35658 143590 35710 143642
rect 35722 143590 35774 143642
rect 35786 143590 35838 143642
rect 35850 143590 35902 143642
rect 66314 143590 66366 143642
rect 66378 143590 66430 143642
rect 66442 143590 66494 143642
rect 66506 143590 66558 143642
rect 66570 143590 66622 143642
rect 97034 143590 97086 143642
rect 97098 143590 97150 143642
rect 97162 143590 97214 143642
rect 97226 143590 97278 143642
rect 97290 143590 97342 143642
rect 4214 143046 4266 143098
rect 4278 143046 4330 143098
rect 4342 143046 4394 143098
rect 4406 143046 4458 143098
rect 4470 143046 4522 143098
rect 34934 143046 34986 143098
rect 34998 143046 35050 143098
rect 35062 143046 35114 143098
rect 35126 143046 35178 143098
rect 35190 143046 35242 143098
rect 65654 143046 65706 143098
rect 65718 143046 65770 143098
rect 65782 143046 65834 143098
rect 65846 143046 65898 143098
rect 65910 143046 65962 143098
rect 96374 143046 96426 143098
rect 96438 143046 96490 143098
rect 96502 143046 96554 143098
rect 96566 143046 96618 143098
rect 96630 143046 96682 143098
rect 4874 142502 4926 142554
rect 4938 142502 4990 142554
rect 5002 142502 5054 142554
rect 5066 142502 5118 142554
rect 5130 142502 5182 142554
rect 35594 142502 35646 142554
rect 35658 142502 35710 142554
rect 35722 142502 35774 142554
rect 35786 142502 35838 142554
rect 35850 142502 35902 142554
rect 66314 142502 66366 142554
rect 66378 142502 66430 142554
rect 66442 142502 66494 142554
rect 66506 142502 66558 142554
rect 66570 142502 66622 142554
rect 97034 142502 97086 142554
rect 97098 142502 97150 142554
rect 97162 142502 97214 142554
rect 97226 142502 97278 142554
rect 97290 142502 97342 142554
rect 4214 141958 4266 142010
rect 4278 141958 4330 142010
rect 4342 141958 4394 142010
rect 4406 141958 4458 142010
rect 4470 141958 4522 142010
rect 34934 141958 34986 142010
rect 34998 141958 35050 142010
rect 35062 141958 35114 142010
rect 35126 141958 35178 142010
rect 35190 141958 35242 142010
rect 65654 141958 65706 142010
rect 65718 141958 65770 142010
rect 65782 141958 65834 142010
rect 65846 141958 65898 142010
rect 65910 141958 65962 142010
rect 96374 141958 96426 142010
rect 96438 141958 96490 142010
rect 96502 141958 96554 142010
rect 96566 141958 96618 142010
rect 96630 141958 96682 142010
rect 4874 141414 4926 141466
rect 4938 141414 4990 141466
rect 5002 141414 5054 141466
rect 5066 141414 5118 141466
rect 5130 141414 5182 141466
rect 35594 141414 35646 141466
rect 35658 141414 35710 141466
rect 35722 141414 35774 141466
rect 35786 141414 35838 141466
rect 35850 141414 35902 141466
rect 66314 141414 66366 141466
rect 66378 141414 66430 141466
rect 66442 141414 66494 141466
rect 66506 141414 66558 141466
rect 66570 141414 66622 141466
rect 97034 141414 97086 141466
rect 97098 141414 97150 141466
rect 97162 141414 97214 141466
rect 97226 141414 97278 141466
rect 97290 141414 97342 141466
rect 4214 140870 4266 140922
rect 4278 140870 4330 140922
rect 4342 140870 4394 140922
rect 4406 140870 4458 140922
rect 4470 140870 4522 140922
rect 34934 140870 34986 140922
rect 34998 140870 35050 140922
rect 35062 140870 35114 140922
rect 35126 140870 35178 140922
rect 35190 140870 35242 140922
rect 65654 140870 65706 140922
rect 65718 140870 65770 140922
rect 65782 140870 65834 140922
rect 65846 140870 65898 140922
rect 65910 140870 65962 140922
rect 96374 140870 96426 140922
rect 96438 140870 96490 140922
rect 96502 140870 96554 140922
rect 96566 140870 96618 140922
rect 96630 140870 96682 140922
rect 4874 140326 4926 140378
rect 4938 140326 4990 140378
rect 5002 140326 5054 140378
rect 5066 140326 5118 140378
rect 5130 140326 5182 140378
rect 35594 140326 35646 140378
rect 35658 140326 35710 140378
rect 35722 140326 35774 140378
rect 35786 140326 35838 140378
rect 35850 140326 35902 140378
rect 66314 140326 66366 140378
rect 66378 140326 66430 140378
rect 66442 140326 66494 140378
rect 66506 140326 66558 140378
rect 66570 140326 66622 140378
rect 97034 140326 97086 140378
rect 97098 140326 97150 140378
rect 97162 140326 97214 140378
rect 97226 140326 97278 140378
rect 97290 140326 97342 140378
rect 4214 139782 4266 139834
rect 4278 139782 4330 139834
rect 4342 139782 4394 139834
rect 4406 139782 4458 139834
rect 4470 139782 4522 139834
rect 34934 139782 34986 139834
rect 34998 139782 35050 139834
rect 35062 139782 35114 139834
rect 35126 139782 35178 139834
rect 35190 139782 35242 139834
rect 65654 139782 65706 139834
rect 65718 139782 65770 139834
rect 65782 139782 65834 139834
rect 65846 139782 65898 139834
rect 65910 139782 65962 139834
rect 96374 139782 96426 139834
rect 96438 139782 96490 139834
rect 96502 139782 96554 139834
rect 96566 139782 96618 139834
rect 96630 139782 96682 139834
rect 4874 139238 4926 139290
rect 4938 139238 4990 139290
rect 5002 139238 5054 139290
rect 5066 139238 5118 139290
rect 5130 139238 5182 139290
rect 35594 139238 35646 139290
rect 35658 139238 35710 139290
rect 35722 139238 35774 139290
rect 35786 139238 35838 139290
rect 35850 139238 35902 139290
rect 66314 139238 66366 139290
rect 66378 139238 66430 139290
rect 66442 139238 66494 139290
rect 66506 139238 66558 139290
rect 66570 139238 66622 139290
rect 97034 139238 97086 139290
rect 97098 139238 97150 139290
rect 97162 139238 97214 139290
rect 97226 139238 97278 139290
rect 97290 139238 97342 139290
rect 4214 138694 4266 138746
rect 4278 138694 4330 138746
rect 4342 138694 4394 138746
rect 4406 138694 4458 138746
rect 4470 138694 4522 138746
rect 34934 138694 34986 138746
rect 34998 138694 35050 138746
rect 35062 138694 35114 138746
rect 35126 138694 35178 138746
rect 35190 138694 35242 138746
rect 65654 138694 65706 138746
rect 65718 138694 65770 138746
rect 65782 138694 65834 138746
rect 65846 138694 65898 138746
rect 65910 138694 65962 138746
rect 96374 138694 96426 138746
rect 96438 138694 96490 138746
rect 96502 138694 96554 138746
rect 96566 138694 96618 138746
rect 96630 138694 96682 138746
rect 4874 138150 4926 138202
rect 4938 138150 4990 138202
rect 5002 138150 5054 138202
rect 5066 138150 5118 138202
rect 5130 138150 5182 138202
rect 35594 138150 35646 138202
rect 35658 138150 35710 138202
rect 35722 138150 35774 138202
rect 35786 138150 35838 138202
rect 35850 138150 35902 138202
rect 66314 138150 66366 138202
rect 66378 138150 66430 138202
rect 66442 138150 66494 138202
rect 66506 138150 66558 138202
rect 66570 138150 66622 138202
rect 97034 138150 97086 138202
rect 97098 138150 97150 138202
rect 97162 138150 97214 138202
rect 97226 138150 97278 138202
rect 97290 138150 97342 138202
rect 4214 137606 4266 137658
rect 4278 137606 4330 137658
rect 4342 137606 4394 137658
rect 4406 137606 4458 137658
rect 4470 137606 4522 137658
rect 34934 137606 34986 137658
rect 34998 137606 35050 137658
rect 35062 137606 35114 137658
rect 35126 137606 35178 137658
rect 35190 137606 35242 137658
rect 65654 137606 65706 137658
rect 65718 137606 65770 137658
rect 65782 137606 65834 137658
rect 65846 137606 65898 137658
rect 65910 137606 65962 137658
rect 96374 137606 96426 137658
rect 96438 137606 96490 137658
rect 96502 137606 96554 137658
rect 96566 137606 96618 137658
rect 96630 137606 96682 137658
rect 4874 137062 4926 137114
rect 4938 137062 4990 137114
rect 5002 137062 5054 137114
rect 5066 137062 5118 137114
rect 5130 137062 5182 137114
rect 35594 137062 35646 137114
rect 35658 137062 35710 137114
rect 35722 137062 35774 137114
rect 35786 137062 35838 137114
rect 35850 137062 35902 137114
rect 66314 137062 66366 137114
rect 66378 137062 66430 137114
rect 66442 137062 66494 137114
rect 66506 137062 66558 137114
rect 66570 137062 66622 137114
rect 97034 137062 97086 137114
rect 97098 137062 97150 137114
rect 97162 137062 97214 137114
rect 97226 137062 97278 137114
rect 97290 137062 97342 137114
rect 4214 136518 4266 136570
rect 4278 136518 4330 136570
rect 4342 136518 4394 136570
rect 4406 136518 4458 136570
rect 4470 136518 4522 136570
rect 34934 136518 34986 136570
rect 34998 136518 35050 136570
rect 35062 136518 35114 136570
rect 35126 136518 35178 136570
rect 35190 136518 35242 136570
rect 65654 136518 65706 136570
rect 65718 136518 65770 136570
rect 65782 136518 65834 136570
rect 65846 136518 65898 136570
rect 65910 136518 65962 136570
rect 96374 136518 96426 136570
rect 96438 136518 96490 136570
rect 96502 136518 96554 136570
rect 96566 136518 96618 136570
rect 96630 136518 96682 136570
rect 105922 136518 105974 136570
rect 105986 136518 106038 136570
rect 106050 136518 106102 136570
rect 106114 136518 106166 136570
rect 106178 136518 106230 136570
rect 9496 136076 9548 136128
rect 101956 136212 102008 136264
rect 38200 136187 38252 136196
rect 38200 136153 38209 136187
rect 38209 136153 38243 136187
rect 38243 136153 38252 136187
rect 38200 136144 38252 136153
rect 40684 136187 40736 136196
rect 40684 136153 40693 136187
rect 40693 136153 40727 136187
rect 40727 136153 40736 136187
rect 40684 136144 40736 136153
rect 42984 136187 43036 136196
rect 42984 136153 42993 136187
rect 42993 136153 43027 136187
rect 43027 136153 43036 136187
rect 42984 136144 43036 136153
rect 46020 136144 46072 136196
rect 48504 136144 48556 136196
rect 52368 136144 52420 136196
rect 55772 136187 55824 136196
rect 55772 136153 55781 136187
rect 55781 136153 55815 136187
rect 55815 136153 55824 136187
rect 55772 136144 55824 136153
rect 58164 136187 58216 136196
rect 58164 136153 58173 136187
rect 58173 136153 58207 136187
rect 58207 136153 58216 136187
rect 58164 136144 58216 136153
rect 60648 136187 60700 136196
rect 60648 136153 60657 136187
rect 60657 136153 60691 136187
rect 60691 136153 60700 136187
rect 60648 136144 60700 136153
rect 63132 136187 63184 136196
rect 63132 136153 63141 136187
rect 63141 136153 63175 136187
rect 63175 136153 63184 136187
rect 63132 136144 63184 136153
rect 64420 136144 64472 136196
rect 67548 136187 67600 136196
rect 67548 136153 67557 136187
rect 67557 136153 67591 136187
rect 67591 136153 67600 136187
rect 67548 136144 67600 136153
rect 69756 136187 69808 136196
rect 69756 136153 69765 136187
rect 69765 136153 69799 136187
rect 69799 136153 69808 136187
rect 69756 136144 69808 136153
rect 72148 136187 72200 136196
rect 72148 136153 72157 136187
rect 72157 136153 72191 136187
rect 72191 136153 72200 136187
rect 72148 136144 72200 136153
rect 74172 136187 74224 136196
rect 74172 136153 74181 136187
rect 74181 136153 74215 136187
rect 74215 136153 74224 136187
rect 74172 136144 74224 136153
rect 36084 136119 36136 136128
rect 36084 136085 36093 136119
rect 36093 136085 36127 136119
rect 36127 136085 36136 136119
rect 36084 136076 36136 136085
rect 38108 136119 38160 136128
rect 38108 136085 38117 136119
rect 38117 136085 38151 136119
rect 38151 136085 38160 136119
rect 38108 136076 38160 136085
rect 40592 136119 40644 136128
rect 40592 136085 40601 136119
rect 40601 136085 40635 136119
rect 40635 136085 40644 136119
rect 40592 136076 40644 136085
rect 42892 136119 42944 136128
rect 42892 136085 42901 136119
rect 42901 136085 42935 136119
rect 42935 136085 42944 136119
rect 42892 136076 42944 136085
rect 45192 136119 45244 136128
rect 45192 136085 45201 136119
rect 45201 136085 45235 136119
rect 45235 136085 45244 136119
rect 45192 136076 45244 136085
rect 56140 136119 56192 136128
rect 56140 136085 56149 136119
rect 56149 136085 56183 136119
rect 56183 136085 56192 136119
rect 56140 136076 56192 136085
rect 58532 136119 58584 136128
rect 58532 136085 58541 136119
rect 58541 136085 58575 136119
rect 58575 136085 58584 136119
rect 58532 136076 58584 136085
rect 61016 136119 61068 136128
rect 61016 136085 61025 136119
rect 61025 136085 61059 136119
rect 61059 136085 61068 136119
rect 61016 136076 61068 136085
rect 63500 136119 63552 136128
rect 63500 136085 63509 136119
rect 63509 136085 63543 136119
rect 63543 136085 63552 136119
rect 63500 136076 63552 136085
rect 65340 136119 65392 136128
rect 65340 136085 65349 136119
rect 65349 136085 65383 136119
rect 65383 136085 65392 136119
rect 65340 136076 65392 136085
rect 67916 136119 67968 136128
rect 67916 136085 67925 136119
rect 67925 136085 67959 136119
rect 67959 136085 67968 136119
rect 67916 136076 67968 136085
rect 70124 136119 70176 136128
rect 70124 136085 70133 136119
rect 70133 136085 70167 136119
rect 70167 136085 70176 136119
rect 70124 136076 70176 136085
rect 72516 136119 72568 136128
rect 72516 136085 72525 136119
rect 72525 136085 72559 136119
rect 72559 136085 72568 136119
rect 72516 136076 72568 136085
rect 77760 136076 77812 136128
rect 86132 136076 86184 136128
rect 87328 136119 87380 136128
rect 87328 136085 87337 136119
rect 87337 136085 87371 136119
rect 87371 136085 87380 136119
rect 87328 136076 87380 136085
rect 95976 136119 96028 136128
rect 95976 136085 95985 136119
rect 95985 136085 96019 136119
rect 96019 136085 96028 136119
rect 95976 136076 96028 136085
rect 4874 135974 4926 136026
rect 4938 135974 4990 136026
rect 5002 135974 5054 136026
rect 5066 135974 5118 136026
rect 5130 135974 5182 136026
rect 35594 135974 35646 136026
rect 35658 135974 35710 136026
rect 35722 135974 35774 136026
rect 35786 135974 35838 136026
rect 35850 135974 35902 136026
rect 66314 135974 66366 136026
rect 66378 135974 66430 136026
rect 66442 135974 66494 136026
rect 66506 135974 66558 136026
rect 66570 135974 66622 136026
rect 97034 135974 97086 136026
rect 97098 135974 97150 136026
rect 97162 135974 97214 136026
rect 97226 135974 97278 136026
rect 97290 135974 97342 136026
rect 106658 135974 106710 136026
rect 106722 135974 106774 136026
rect 106786 135974 106838 136026
rect 106850 135974 106902 136026
rect 106914 135974 106966 136026
rect 8116 135872 8168 135924
rect 45192 135872 45244 135924
rect 56140 135872 56192 135924
rect 102140 135872 102192 135924
rect 8208 135804 8260 135856
rect 42892 135804 42944 135856
rect 58532 135804 58584 135856
rect 103980 135804 104032 135856
rect 9588 135736 9640 135788
rect 40592 135736 40644 135788
rect 61016 135736 61068 135788
rect 102324 135736 102376 135788
rect 8024 135668 8076 135720
rect 38108 135668 38160 135720
rect 63500 135668 63552 135720
rect 102416 135668 102468 135720
rect 65340 135600 65392 135652
rect 103612 135600 103664 135652
rect 67916 135532 67968 135584
rect 103704 135532 103756 135584
rect 4214 135430 4266 135482
rect 4278 135430 4330 135482
rect 4342 135430 4394 135482
rect 4406 135430 4458 135482
rect 4470 135430 4522 135482
rect 70124 135464 70176 135516
rect 102508 135464 102560 135516
rect 72516 135396 72568 135448
rect 103888 135396 103940 135448
rect 105922 135430 105974 135482
rect 105986 135430 106038 135482
rect 106050 135430 106102 135482
rect 106114 135430 106166 135482
rect 106178 135430 106230 135482
rect 77760 135328 77812 135380
rect 103796 135328 103848 135380
rect 4874 134886 4926 134938
rect 4938 134886 4990 134938
rect 5002 134886 5054 134938
rect 5066 134886 5118 134938
rect 5130 134886 5182 134938
rect 106658 134886 106710 134938
rect 106722 134886 106774 134938
rect 106786 134886 106838 134938
rect 106850 134886 106902 134938
rect 106914 134886 106966 134938
rect 95976 134512 96028 134564
rect 103520 134512 103572 134564
rect 4214 134342 4266 134394
rect 4278 134342 4330 134394
rect 4342 134342 4394 134394
rect 4406 134342 4458 134394
rect 4470 134342 4522 134394
rect 105922 134342 105974 134394
rect 105986 134342 106038 134394
rect 106050 134342 106102 134394
rect 106114 134342 106166 134394
rect 106178 134342 106230 134394
rect 87328 133968 87380 134020
rect 102232 133968 102284 134020
rect 7932 133900 7984 133952
rect 36084 133900 36136 133952
rect 86132 133900 86184 133952
rect 102600 133900 102652 133952
rect 4874 133798 4926 133850
rect 4938 133798 4990 133850
rect 5002 133798 5054 133850
rect 5066 133798 5118 133850
rect 5130 133798 5182 133850
rect 106658 133798 106710 133850
rect 106722 133798 106774 133850
rect 106786 133798 106838 133850
rect 106850 133798 106902 133850
rect 106914 133798 106966 133850
rect 4214 133254 4266 133306
rect 4278 133254 4330 133306
rect 4342 133254 4394 133306
rect 4406 133254 4458 133306
rect 4470 133254 4522 133306
rect 105922 133254 105974 133306
rect 105986 133254 106038 133306
rect 106050 133254 106102 133306
rect 106114 133254 106166 133306
rect 106178 133254 106230 133306
rect 4874 132710 4926 132762
rect 4938 132710 4990 132762
rect 5002 132710 5054 132762
rect 5066 132710 5118 132762
rect 5130 132710 5182 132762
rect 106658 132710 106710 132762
rect 106722 132710 106774 132762
rect 106786 132710 106838 132762
rect 106850 132710 106902 132762
rect 106914 132710 106966 132762
rect 4214 132166 4266 132218
rect 4278 132166 4330 132218
rect 4342 132166 4394 132218
rect 4406 132166 4458 132218
rect 4470 132166 4522 132218
rect 105922 132166 105974 132218
rect 105986 132166 106038 132218
rect 106050 132166 106102 132218
rect 106114 132166 106166 132218
rect 106178 132166 106230 132218
rect 4874 131622 4926 131674
rect 4938 131622 4990 131674
rect 5002 131622 5054 131674
rect 5066 131622 5118 131674
rect 5130 131622 5182 131674
rect 106658 131622 106710 131674
rect 106722 131622 106774 131674
rect 106786 131622 106838 131674
rect 106850 131622 106902 131674
rect 106914 131622 106966 131674
rect 4214 131078 4266 131130
rect 4278 131078 4330 131130
rect 4342 131078 4394 131130
rect 4406 131078 4458 131130
rect 4470 131078 4522 131130
rect 105922 131078 105974 131130
rect 105986 131078 106038 131130
rect 106050 131078 106102 131130
rect 106114 131078 106166 131130
rect 106178 131078 106230 131130
rect 4874 130534 4926 130586
rect 4938 130534 4990 130586
rect 5002 130534 5054 130586
rect 5066 130534 5118 130586
rect 5130 130534 5182 130586
rect 106658 130534 106710 130586
rect 106722 130534 106774 130586
rect 106786 130534 106838 130586
rect 106850 130534 106902 130586
rect 106914 130534 106966 130586
rect 4214 129990 4266 130042
rect 4278 129990 4330 130042
rect 4342 129990 4394 130042
rect 4406 129990 4458 130042
rect 4470 129990 4522 130042
rect 105922 129990 105974 130042
rect 105986 129990 106038 130042
rect 106050 129990 106102 130042
rect 106114 129990 106166 130042
rect 106178 129990 106230 130042
rect 104348 129863 104400 129872
rect 104348 129829 104357 129863
rect 104357 129829 104391 129863
rect 104391 129829 104400 129863
rect 104348 129820 104400 129829
rect 4874 129446 4926 129498
rect 4938 129446 4990 129498
rect 5002 129446 5054 129498
rect 5066 129446 5118 129498
rect 5130 129446 5182 129498
rect 106658 129446 106710 129498
rect 106722 129446 106774 129498
rect 106786 129446 106838 129498
rect 106850 129446 106902 129498
rect 106914 129446 106966 129498
rect 4214 128902 4266 128954
rect 4278 128902 4330 128954
rect 4342 128902 4394 128954
rect 4406 128902 4458 128954
rect 4470 128902 4522 128954
rect 105922 128902 105974 128954
rect 105986 128902 106038 128954
rect 106050 128902 106102 128954
rect 106114 128902 106166 128954
rect 106178 128902 106230 128954
rect 4874 128358 4926 128410
rect 4938 128358 4990 128410
rect 5002 128358 5054 128410
rect 5066 128358 5118 128410
rect 5130 128358 5182 128410
rect 106658 128358 106710 128410
rect 106722 128358 106774 128410
rect 106786 128358 106838 128410
rect 106850 128358 106902 128410
rect 106914 128358 106966 128410
rect 4214 127814 4266 127866
rect 4278 127814 4330 127866
rect 4342 127814 4394 127866
rect 4406 127814 4458 127866
rect 4470 127814 4522 127866
rect 105922 127814 105974 127866
rect 105986 127814 106038 127866
rect 106050 127814 106102 127866
rect 106114 127814 106166 127866
rect 106178 127814 106230 127866
rect 4874 127270 4926 127322
rect 4938 127270 4990 127322
rect 5002 127270 5054 127322
rect 5066 127270 5118 127322
rect 5130 127270 5182 127322
rect 106658 127270 106710 127322
rect 106722 127270 106774 127322
rect 106786 127270 106838 127322
rect 106850 127270 106902 127322
rect 106914 127270 106966 127322
rect 4214 126726 4266 126778
rect 4278 126726 4330 126778
rect 4342 126726 4394 126778
rect 4406 126726 4458 126778
rect 4470 126726 4522 126778
rect 105922 126726 105974 126778
rect 105986 126726 106038 126778
rect 106050 126726 106102 126778
rect 106114 126726 106166 126778
rect 106178 126726 106230 126778
rect 4874 126182 4926 126234
rect 4938 126182 4990 126234
rect 5002 126182 5054 126234
rect 5066 126182 5118 126234
rect 5130 126182 5182 126234
rect 106658 126182 106710 126234
rect 106722 126182 106774 126234
rect 106786 126182 106838 126234
rect 106850 126182 106902 126234
rect 106914 126182 106966 126234
rect 4214 125638 4266 125690
rect 4278 125638 4330 125690
rect 4342 125638 4394 125690
rect 4406 125638 4458 125690
rect 4470 125638 4522 125690
rect 105922 125638 105974 125690
rect 105986 125638 106038 125690
rect 106050 125638 106102 125690
rect 106114 125638 106166 125690
rect 106178 125638 106230 125690
rect 4874 125094 4926 125146
rect 4938 125094 4990 125146
rect 5002 125094 5054 125146
rect 5066 125094 5118 125146
rect 5130 125094 5182 125146
rect 106658 125094 106710 125146
rect 106722 125094 106774 125146
rect 106786 125094 106838 125146
rect 106850 125094 106902 125146
rect 106914 125094 106966 125146
rect 4214 124550 4266 124602
rect 4278 124550 4330 124602
rect 4342 124550 4394 124602
rect 4406 124550 4458 124602
rect 4470 124550 4522 124602
rect 105922 124550 105974 124602
rect 105986 124550 106038 124602
rect 106050 124550 106102 124602
rect 106114 124550 106166 124602
rect 106178 124550 106230 124602
rect 4874 124006 4926 124058
rect 4938 124006 4990 124058
rect 5002 124006 5054 124058
rect 5066 124006 5118 124058
rect 5130 124006 5182 124058
rect 106658 124006 106710 124058
rect 106722 124006 106774 124058
rect 106786 124006 106838 124058
rect 106850 124006 106902 124058
rect 106914 124006 106966 124058
rect 4214 123462 4266 123514
rect 4278 123462 4330 123514
rect 4342 123462 4394 123514
rect 4406 123462 4458 123514
rect 4470 123462 4522 123514
rect 105922 123462 105974 123514
rect 105986 123462 106038 123514
rect 106050 123462 106102 123514
rect 106114 123462 106166 123514
rect 106178 123462 106230 123514
rect 4874 122918 4926 122970
rect 4938 122918 4990 122970
rect 5002 122918 5054 122970
rect 5066 122918 5118 122970
rect 5130 122918 5182 122970
rect 106658 122918 106710 122970
rect 106722 122918 106774 122970
rect 106786 122918 106838 122970
rect 106850 122918 106902 122970
rect 106914 122918 106966 122970
rect 4214 122374 4266 122426
rect 4278 122374 4330 122426
rect 4342 122374 4394 122426
rect 4406 122374 4458 122426
rect 4470 122374 4522 122426
rect 105922 122374 105974 122426
rect 105986 122374 106038 122426
rect 106050 122374 106102 122426
rect 106114 122374 106166 122426
rect 106178 122374 106230 122426
rect 4874 121830 4926 121882
rect 4938 121830 4990 121882
rect 5002 121830 5054 121882
rect 5066 121830 5118 121882
rect 5130 121830 5182 121882
rect 106658 121830 106710 121882
rect 106722 121830 106774 121882
rect 106786 121830 106838 121882
rect 106850 121830 106902 121882
rect 106914 121830 106966 121882
rect 4214 121286 4266 121338
rect 4278 121286 4330 121338
rect 4342 121286 4394 121338
rect 4406 121286 4458 121338
rect 4470 121286 4522 121338
rect 105922 121286 105974 121338
rect 105986 121286 106038 121338
rect 106050 121286 106102 121338
rect 106114 121286 106166 121338
rect 106178 121286 106230 121338
rect 4874 120742 4926 120794
rect 4938 120742 4990 120794
rect 5002 120742 5054 120794
rect 5066 120742 5118 120794
rect 5130 120742 5182 120794
rect 106658 120742 106710 120794
rect 106722 120742 106774 120794
rect 106786 120742 106838 120794
rect 106850 120742 106902 120794
rect 106914 120742 106966 120794
rect 4214 120198 4266 120250
rect 4278 120198 4330 120250
rect 4342 120198 4394 120250
rect 4406 120198 4458 120250
rect 4470 120198 4522 120250
rect 105922 120198 105974 120250
rect 105986 120198 106038 120250
rect 106050 120198 106102 120250
rect 106114 120198 106166 120250
rect 106178 120198 106230 120250
rect 4874 119654 4926 119706
rect 4938 119654 4990 119706
rect 5002 119654 5054 119706
rect 5066 119654 5118 119706
rect 5130 119654 5182 119706
rect 106658 119654 106710 119706
rect 106722 119654 106774 119706
rect 106786 119654 106838 119706
rect 106850 119654 106902 119706
rect 106914 119654 106966 119706
rect 4214 119110 4266 119162
rect 4278 119110 4330 119162
rect 4342 119110 4394 119162
rect 4406 119110 4458 119162
rect 4470 119110 4522 119162
rect 105922 119110 105974 119162
rect 105986 119110 106038 119162
rect 106050 119110 106102 119162
rect 106114 119110 106166 119162
rect 106178 119110 106230 119162
rect 4874 118566 4926 118618
rect 4938 118566 4990 118618
rect 5002 118566 5054 118618
rect 5066 118566 5118 118618
rect 5130 118566 5182 118618
rect 106658 118566 106710 118618
rect 106722 118566 106774 118618
rect 106786 118566 106838 118618
rect 106850 118566 106902 118618
rect 106914 118566 106966 118618
rect 4214 118022 4266 118074
rect 4278 118022 4330 118074
rect 4342 118022 4394 118074
rect 4406 118022 4458 118074
rect 4470 118022 4522 118074
rect 105922 118022 105974 118074
rect 105986 118022 106038 118074
rect 106050 118022 106102 118074
rect 106114 118022 106166 118074
rect 106178 118022 106230 118074
rect 4874 117478 4926 117530
rect 4938 117478 4990 117530
rect 5002 117478 5054 117530
rect 5066 117478 5118 117530
rect 5130 117478 5182 117530
rect 106658 117478 106710 117530
rect 106722 117478 106774 117530
rect 106786 117478 106838 117530
rect 106850 117478 106902 117530
rect 106914 117478 106966 117530
rect 4214 116934 4266 116986
rect 4278 116934 4330 116986
rect 4342 116934 4394 116986
rect 4406 116934 4458 116986
rect 4470 116934 4522 116986
rect 105922 116934 105974 116986
rect 105986 116934 106038 116986
rect 106050 116934 106102 116986
rect 106114 116934 106166 116986
rect 106178 116934 106230 116986
rect 4874 116390 4926 116442
rect 4938 116390 4990 116442
rect 5002 116390 5054 116442
rect 5066 116390 5118 116442
rect 5130 116390 5182 116442
rect 106658 116390 106710 116442
rect 106722 116390 106774 116442
rect 106786 116390 106838 116442
rect 106850 116390 106902 116442
rect 106914 116390 106966 116442
rect 4214 115846 4266 115898
rect 4278 115846 4330 115898
rect 4342 115846 4394 115898
rect 4406 115846 4458 115898
rect 4470 115846 4522 115898
rect 105922 115846 105974 115898
rect 105986 115846 106038 115898
rect 106050 115846 106102 115898
rect 106114 115846 106166 115898
rect 106178 115846 106230 115898
rect 4874 115302 4926 115354
rect 4938 115302 4990 115354
rect 5002 115302 5054 115354
rect 5066 115302 5118 115354
rect 5130 115302 5182 115354
rect 106658 115302 106710 115354
rect 106722 115302 106774 115354
rect 106786 115302 106838 115354
rect 106850 115302 106902 115354
rect 106914 115302 106966 115354
rect 4214 114758 4266 114810
rect 4278 114758 4330 114810
rect 4342 114758 4394 114810
rect 4406 114758 4458 114810
rect 4470 114758 4522 114810
rect 105922 114758 105974 114810
rect 105986 114758 106038 114810
rect 106050 114758 106102 114810
rect 106114 114758 106166 114810
rect 106178 114758 106230 114810
rect 4874 114214 4926 114266
rect 4938 114214 4990 114266
rect 5002 114214 5054 114266
rect 5066 114214 5118 114266
rect 5130 114214 5182 114266
rect 106658 114214 106710 114266
rect 106722 114214 106774 114266
rect 106786 114214 106838 114266
rect 106850 114214 106902 114266
rect 106914 114214 106966 114266
rect 4214 113670 4266 113722
rect 4278 113670 4330 113722
rect 4342 113670 4394 113722
rect 4406 113670 4458 113722
rect 4470 113670 4522 113722
rect 105922 113670 105974 113722
rect 105986 113670 106038 113722
rect 106050 113670 106102 113722
rect 106114 113670 106166 113722
rect 106178 113670 106230 113722
rect 4874 113126 4926 113178
rect 4938 113126 4990 113178
rect 5002 113126 5054 113178
rect 5066 113126 5118 113178
rect 5130 113126 5182 113178
rect 106658 113126 106710 113178
rect 106722 113126 106774 113178
rect 106786 113126 106838 113178
rect 106850 113126 106902 113178
rect 106914 113126 106966 113178
rect 4214 112582 4266 112634
rect 4278 112582 4330 112634
rect 4342 112582 4394 112634
rect 4406 112582 4458 112634
rect 4470 112582 4522 112634
rect 105922 112582 105974 112634
rect 105986 112582 106038 112634
rect 106050 112582 106102 112634
rect 106114 112582 106166 112634
rect 106178 112582 106230 112634
rect 4874 112038 4926 112090
rect 4938 112038 4990 112090
rect 5002 112038 5054 112090
rect 5066 112038 5118 112090
rect 5130 112038 5182 112090
rect 106658 112038 106710 112090
rect 106722 112038 106774 112090
rect 106786 112038 106838 112090
rect 106850 112038 106902 112090
rect 106914 112038 106966 112090
rect 4214 111494 4266 111546
rect 4278 111494 4330 111546
rect 4342 111494 4394 111546
rect 4406 111494 4458 111546
rect 4470 111494 4522 111546
rect 105922 111494 105974 111546
rect 105986 111494 106038 111546
rect 106050 111494 106102 111546
rect 106114 111494 106166 111546
rect 106178 111494 106230 111546
rect 8392 111324 8444 111376
rect 1308 111188 1360 111240
rect 4874 110950 4926 111002
rect 4938 110950 4990 111002
rect 5002 110950 5054 111002
rect 5066 110950 5118 111002
rect 5130 110950 5182 111002
rect 106658 110950 106710 111002
rect 106722 110950 106774 111002
rect 106786 110950 106838 111002
rect 106850 110950 106902 111002
rect 106914 110950 106966 111002
rect 4214 110406 4266 110458
rect 4278 110406 4330 110458
rect 4342 110406 4394 110458
rect 4406 110406 4458 110458
rect 4470 110406 4522 110458
rect 105922 110406 105974 110458
rect 105986 110406 106038 110458
rect 106050 110406 106102 110458
rect 106114 110406 106166 110458
rect 106178 110406 106230 110458
rect 4874 109862 4926 109914
rect 4938 109862 4990 109914
rect 5002 109862 5054 109914
rect 5066 109862 5118 109914
rect 5130 109862 5182 109914
rect 106658 109862 106710 109914
rect 106722 109862 106774 109914
rect 106786 109862 106838 109914
rect 106850 109862 106902 109914
rect 106914 109862 106966 109914
rect 1308 109624 1360 109676
rect 8392 109488 8444 109540
rect 4214 109318 4266 109370
rect 4278 109318 4330 109370
rect 4342 109318 4394 109370
rect 4406 109318 4458 109370
rect 4470 109318 4522 109370
rect 105922 109318 105974 109370
rect 105986 109318 106038 109370
rect 106050 109318 106102 109370
rect 106114 109318 106166 109370
rect 106178 109318 106230 109370
rect 4874 108774 4926 108826
rect 4938 108774 4990 108826
rect 5002 108774 5054 108826
rect 5066 108774 5118 108826
rect 5130 108774 5182 108826
rect 106658 108774 106710 108826
rect 106722 108774 106774 108826
rect 106786 108774 106838 108826
rect 106850 108774 106902 108826
rect 106914 108774 106966 108826
rect 1308 108536 1360 108588
rect 8392 108400 8444 108452
rect 4214 108230 4266 108282
rect 4278 108230 4330 108282
rect 4342 108230 4394 108282
rect 4406 108230 4458 108282
rect 4470 108230 4522 108282
rect 105922 108230 105974 108282
rect 105986 108230 106038 108282
rect 106050 108230 106102 108282
rect 106114 108230 106166 108282
rect 106178 108230 106230 108282
rect 4874 107686 4926 107738
rect 4938 107686 4990 107738
rect 5002 107686 5054 107738
rect 5066 107686 5118 107738
rect 5130 107686 5182 107738
rect 106658 107686 106710 107738
rect 106722 107686 106774 107738
rect 106786 107686 106838 107738
rect 106850 107686 106902 107738
rect 106914 107686 106966 107738
rect 4214 107142 4266 107194
rect 4278 107142 4330 107194
rect 4342 107142 4394 107194
rect 4406 107142 4458 107194
rect 4470 107142 4522 107194
rect 105922 107142 105974 107194
rect 105986 107142 106038 107194
rect 106050 107142 106102 107194
rect 106114 107142 106166 107194
rect 106178 107142 106230 107194
rect 8392 106972 8444 107024
rect 1216 106836 1268 106888
rect 4874 106598 4926 106650
rect 4938 106598 4990 106650
rect 5002 106598 5054 106650
rect 5066 106598 5118 106650
rect 5130 106598 5182 106650
rect 106658 106598 106710 106650
rect 106722 106598 106774 106650
rect 106786 106598 106838 106650
rect 106850 106598 106902 106650
rect 106914 106598 106966 106650
rect 4214 106054 4266 106106
rect 4278 106054 4330 106106
rect 4342 106054 4394 106106
rect 4406 106054 4458 106106
rect 4470 106054 4522 106106
rect 105922 106054 105974 106106
rect 105986 106054 106038 106106
rect 106050 106054 106102 106106
rect 106114 106054 106166 106106
rect 106178 106054 106230 106106
rect 8392 105884 8444 105936
rect 1308 105748 1360 105800
rect 4874 105510 4926 105562
rect 4938 105510 4990 105562
rect 5002 105510 5054 105562
rect 5066 105510 5118 105562
rect 5130 105510 5182 105562
rect 106658 105510 106710 105562
rect 106722 105510 106774 105562
rect 106786 105510 106838 105562
rect 106850 105510 106902 105562
rect 106914 105510 106966 105562
rect 4214 104966 4266 105018
rect 4278 104966 4330 105018
rect 4342 104966 4394 105018
rect 4406 104966 4458 105018
rect 4470 104966 4522 105018
rect 105922 104966 105974 105018
rect 105986 104966 106038 105018
rect 106050 104966 106102 105018
rect 106114 104966 106166 105018
rect 106178 104966 106230 105018
rect 4874 104422 4926 104474
rect 4938 104422 4990 104474
rect 5002 104422 5054 104474
rect 5066 104422 5118 104474
rect 5130 104422 5182 104474
rect 106658 104422 106710 104474
rect 106722 104422 106774 104474
rect 106786 104422 106838 104474
rect 106850 104422 106902 104474
rect 106914 104422 106966 104474
rect 1308 104184 1360 104236
rect 8392 104048 8444 104100
rect 4214 103878 4266 103930
rect 4278 103878 4330 103930
rect 4342 103878 4394 103930
rect 4406 103878 4458 103930
rect 4470 103878 4522 103930
rect 105922 103878 105974 103930
rect 105986 103878 106038 103930
rect 106050 103878 106102 103930
rect 106114 103878 106166 103930
rect 106178 103878 106230 103930
rect 4874 103334 4926 103386
rect 4938 103334 4990 103386
rect 5002 103334 5054 103386
rect 5066 103334 5118 103386
rect 5130 103334 5182 103386
rect 106658 103334 106710 103386
rect 106722 103334 106774 103386
rect 106786 103334 106838 103386
rect 106850 103334 106902 103386
rect 106914 103334 106966 103386
rect 4214 102790 4266 102842
rect 4278 102790 4330 102842
rect 4342 102790 4394 102842
rect 4406 102790 4458 102842
rect 4470 102790 4522 102842
rect 105922 102790 105974 102842
rect 105986 102790 106038 102842
rect 106050 102790 106102 102842
rect 106114 102790 106166 102842
rect 106178 102790 106230 102842
rect 4874 102246 4926 102298
rect 4938 102246 4990 102298
rect 5002 102246 5054 102298
rect 5066 102246 5118 102298
rect 5130 102246 5182 102298
rect 106658 102246 106710 102298
rect 106722 102246 106774 102298
rect 106786 102246 106838 102298
rect 106850 102246 106902 102298
rect 106914 102246 106966 102298
rect 4214 101702 4266 101754
rect 4278 101702 4330 101754
rect 4342 101702 4394 101754
rect 4406 101702 4458 101754
rect 4470 101702 4522 101754
rect 105922 101702 105974 101754
rect 105986 101702 106038 101754
rect 106050 101702 106102 101754
rect 106114 101702 106166 101754
rect 106178 101702 106230 101754
rect 4874 101158 4926 101210
rect 4938 101158 4990 101210
rect 5002 101158 5054 101210
rect 5066 101158 5118 101210
rect 5130 101158 5182 101210
rect 106658 101158 106710 101210
rect 106722 101158 106774 101210
rect 106786 101158 106838 101210
rect 106850 101158 106902 101210
rect 106914 101158 106966 101210
rect 4214 100614 4266 100666
rect 4278 100614 4330 100666
rect 4342 100614 4394 100666
rect 4406 100614 4458 100666
rect 4470 100614 4522 100666
rect 105922 100614 105974 100666
rect 105986 100614 106038 100666
rect 106050 100614 106102 100666
rect 106114 100614 106166 100666
rect 106178 100614 106230 100666
rect 4874 100070 4926 100122
rect 4938 100070 4990 100122
rect 5002 100070 5054 100122
rect 5066 100070 5118 100122
rect 5130 100070 5182 100122
rect 106658 100070 106710 100122
rect 106722 100070 106774 100122
rect 106786 100070 106838 100122
rect 106850 100070 106902 100122
rect 106914 100070 106966 100122
rect 4214 99526 4266 99578
rect 4278 99526 4330 99578
rect 4342 99526 4394 99578
rect 4406 99526 4458 99578
rect 4470 99526 4522 99578
rect 105922 99526 105974 99578
rect 105986 99526 106038 99578
rect 106050 99526 106102 99578
rect 106114 99526 106166 99578
rect 106178 99526 106230 99578
rect 4874 98982 4926 99034
rect 4938 98982 4990 99034
rect 5002 98982 5054 99034
rect 5066 98982 5118 99034
rect 5130 98982 5182 99034
rect 106658 98982 106710 99034
rect 106722 98982 106774 99034
rect 106786 98982 106838 99034
rect 106850 98982 106902 99034
rect 106914 98982 106966 99034
rect 4214 98438 4266 98490
rect 4278 98438 4330 98490
rect 4342 98438 4394 98490
rect 4406 98438 4458 98490
rect 4470 98438 4522 98490
rect 105922 98438 105974 98490
rect 105986 98438 106038 98490
rect 106050 98438 106102 98490
rect 106114 98438 106166 98490
rect 106178 98438 106230 98490
rect 4874 97894 4926 97946
rect 4938 97894 4990 97946
rect 5002 97894 5054 97946
rect 5066 97894 5118 97946
rect 5130 97894 5182 97946
rect 106658 97894 106710 97946
rect 106722 97894 106774 97946
rect 106786 97894 106838 97946
rect 106850 97894 106902 97946
rect 106914 97894 106966 97946
rect 4214 97350 4266 97402
rect 4278 97350 4330 97402
rect 4342 97350 4394 97402
rect 4406 97350 4458 97402
rect 4470 97350 4522 97402
rect 105922 97350 105974 97402
rect 105986 97350 106038 97402
rect 106050 97350 106102 97402
rect 106114 97350 106166 97402
rect 106178 97350 106230 97402
rect 4874 96806 4926 96858
rect 4938 96806 4990 96858
rect 5002 96806 5054 96858
rect 5066 96806 5118 96858
rect 5130 96806 5182 96858
rect 106658 96806 106710 96858
rect 106722 96806 106774 96858
rect 106786 96806 106838 96858
rect 106850 96806 106902 96858
rect 106914 96806 106966 96858
rect 4214 96262 4266 96314
rect 4278 96262 4330 96314
rect 4342 96262 4394 96314
rect 4406 96262 4458 96314
rect 4470 96262 4522 96314
rect 105922 96262 105974 96314
rect 105986 96262 106038 96314
rect 106050 96262 106102 96314
rect 106114 96262 106166 96314
rect 106178 96262 106230 96314
rect 4874 95718 4926 95770
rect 4938 95718 4990 95770
rect 5002 95718 5054 95770
rect 5066 95718 5118 95770
rect 5130 95718 5182 95770
rect 106658 95718 106710 95770
rect 106722 95718 106774 95770
rect 106786 95718 106838 95770
rect 106850 95718 106902 95770
rect 106914 95718 106966 95770
rect 102692 95276 102744 95328
rect 4214 95174 4266 95226
rect 4278 95174 4330 95226
rect 4342 95174 4394 95226
rect 4406 95174 4458 95226
rect 4470 95174 4522 95226
rect 105922 95174 105974 95226
rect 105986 95174 106038 95226
rect 106050 95174 106102 95226
rect 106114 95174 106166 95226
rect 106178 95174 106230 95226
rect 4874 94630 4926 94682
rect 4938 94630 4990 94682
rect 5002 94630 5054 94682
rect 5066 94630 5118 94682
rect 5130 94630 5182 94682
rect 106658 94630 106710 94682
rect 106722 94630 106774 94682
rect 106786 94630 106838 94682
rect 106850 94630 106902 94682
rect 106914 94630 106966 94682
rect 4214 94086 4266 94138
rect 4278 94086 4330 94138
rect 4342 94086 4394 94138
rect 4406 94086 4458 94138
rect 4470 94086 4522 94138
rect 105922 94086 105974 94138
rect 105986 94086 106038 94138
rect 106050 94086 106102 94138
rect 106114 94086 106166 94138
rect 106178 94086 106230 94138
rect 103060 93848 103112 93900
rect 4874 93542 4926 93594
rect 4938 93542 4990 93594
rect 5002 93542 5054 93594
rect 5066 93542 5118 93594
rect 5130 93542 5182 93594
rect 106658 93542 106710 93594
rect 106722 93542 106774 93594
rect 106786 93542 106838 93594
rect 106850 93542 106902 93594
rect 106914 93542 106966 93594
rect 4214 92998 4266 93050
rect 4278 92998 4330 93050
rect 4342 92998 4394 93050
rect 4406 92998 4458 93050
rect 4470 92998 4522 93050
rect 105922 92998 105974 93050
rect 105986 92998 106038 93050
rect 106050 92998 106102 93050
rect 106114 92998 106166 93050
rect 106178 92998 106230 93050
rect 102968 92556 103020 92608
rect 4874 92454 4926 92506
rect 4938 92454 4990 92506
rect 5002 92454 5054 92506
rect 5066 92454 5118 92506
rect 5130 92454 5182 92506
rect 106658 92454 106710 92506
rect 106722 92454 106774 92506
rect 106786 92454 106838 92506
rect 106850 92454 106902 92506
rect 106914 92454 106966 92506
rect 4214 91910 4266 91962
rect 4278 91910 4330 91962
rect 4342 91910 4394 91962
rect 4406 91910 4458 91962
rect 4470 91910 4522 91962
rect 105922 91910 105974 91962
rect 105986 91910 106038 91962
rect 106050 91910 106102 91962
rect 106114 91910 106166 91962
rect 106178 91910 106230 91962
rect 4874 91366 4926 91418
rect 4938 91366 4990 91418
rect 5002 91366 5054 91418
rect 5066 91366 5118 91418
rect 5130 91366 5182 91418
rect 106658 91366 106710 91418
rect 106722 91366 106774 91418
rect 106786 91366 106838 91418
rect 106850 91366 106902 91418
rect 106914 91366 106966 91418
rect 104348 91171 104400 91180
rect 104348 91137 104357 91171
rect 104357 91137 104391 91171
rect 104391 91137 104400 91171
rect 104348 91128 104400 91137
rect 103520 90924 103572 90976
rect 104164 90924 104216 90976
rect 4214 90822 4266 90874
rect 4278 90822 4330 90874
rect 4342 90822 4394 90874
rect 4406 90822 4458 90874
rect 4470 90822 4522 90874
rect 105922 90822 105974 90874
rect 105986 90822 106038 90874
rect 106050 90822 106102 90874
rect 106114 90822 106166 90874
rect 106178 90822 106230 90874
rect 104348 90423 104400 90432
rect 104348 90389 104357 90423
rect 104357 90389 104391 90423
rect 104391 90389 104400 90423
rect 104348 90380 104400 90389
rect 4874 90278 4926 90330
rect 4938 90278 4990 90330
rect 5002 90278 5054 90330
rect 5066 90278 5118 90330
rect 5130 90278 5182 90330
rect 106658 90278 106710 90330
rect 106722 90278 106774 90330
rect 106786 90278 106838 90330
rect 106850 90278 106902 90330
rect 106914 90278 106966 90330
rect 4214 89734 4266 89786
rect 4278 89734 4330 89786
rect 4342 89734 4394 89786
rect 4406 89734 4458 89786
rect 4470 89734 4522 89786
rect 105922 89734 105974 89786
rect 105986 89734 106038 89786
rect 106050 89734 106102 89786
rect 106114 89734 106166 89786
rect 106178 89734 106230 89786
rect 4874 89190 4926 89242
rect 4938 89190 4990 89242
rect 5002 89190 5054 89242
rect 5066 89190 5118 89242
rect 5130 89190 5182 89242
rect 106658 89190 106710 89242
rect 106722 89190 106774 89242
rect 106786 89190 106838 89242
rect 106850 89190 106902 89242
rect 106914 89190 106966 89242
rect 1308 88952 1360 89004
rect 7564 88816 7616 88868
rect 4214 88646 4266 88698
rect 4278 88646 4330 88698
rect 4342 88646 4394 88698
rect 4406 88646 4458 88698
rect 4470 88646 4522 88698
rect 105922 88646 105974 88698
rect 105986 88646 106038 88698
rect 106050 88646 106102 88698
rect 106114 88646 106166 88698
rect 106178 88646 106230 88698
rect 4874 88102 4926 88154
rect 4938 88102 4990 88154
rect 5002 88102 5054 88154
rect 5066 88102 5118 88154
rect 5130 88102 5182 88154
rect 106658 88102 106710 88154
rect 106722 88102 106774 88154
rect 106786 88102 106838 88154
rect 106850 88102 106902 88154
rect 106914 88102 106966 88154
rect 1216 87864 1268 87916
rect 8944 87728 8996 87780
rect 4214 87558 4266 87610
rect 4278 87558 4330 87610
rect 4342 87558 4394 87610
rect 4406 87558 4458 87610
rect 4470 87558 4522 87610
rect 105922 87558 105974 87610
rect 105986 87558 106038 87610
rect 106050 87558 106102 87610
rect 106114 87558 106166 87610
rect 106178 87558 106230 87610
rect 1216 87184 1268 87236
rect 1860 87159 1912 87168
rect 1860 87125 1869 87159
rect 1869 87125 1903 87159
rect 1903 87125 1912 87159
rect 1860 87116 1912 87125
rect 4874 87014 4926 87066
rect 4938 87014 4990 87066
rect 5002 87014 5054 87066
rect 5066 87014 5118 87066
rect 5130 87014 5182 87066
rect 106658 87014 106710 87066
rect 106722 87014 106774 87066
rect 106786 87014 106838 87066
rect 106850 87014 106902 87066
rect 106914 87014 106966 87066
rect 1308 86776 1360 86828
rect 8668 86640 8720 86692
rect 4214 86470 4266 86522
rect 4278 86470 4330 86522
rect 4342 86470 4394 86522
rect 4406 86470 4458 86522
rect 4470 86470 4522 86522
rect 105922 86470 105974 86522
rect 105986 86470 106038 86522
rect 106050 86470 106102 86522
rect 106114 86470 106166 86522
rect 106178 86470 106230 86522
rect 1308 86164 1360 86216
rect 1860 86096 1912 86148
rect 8576 86096 8628 86148
rect 6000 86028 6052 86080
rect 4874 85926 4926 85978
rect 4938 85926 4990 85978
rect 5002 85926 5054 85978
rect 5066 85926 5118 85978
rect 5130 85926 5182 85978
rect 106658 85926 106710 85978
rect 106722 85926 106774 85978
rect 106786 85926 106838 85978
rect 106850 85926 106902 85978
rect 106914 85926 106966 85978
rect 4214 85382 4266 85434
rect 4278 85382 4330 85434
rect 4342 85382 4394 85434
rect 4406 85382 4458 85434
rect 4470 85382 4522 85434
rect 105922 85382 105974 85434
rect 105986 85382 106038 85434
rect 106050 85382 106102 85434
rect 106114 85382 106166 85434
rect 106178 85382 106230 85434
rect 1216 85008 1268 85060
rect 1768 84983 1820 84992
rect 1768 84949 1777 84983
rect 1777 84949 1811 84983
rect 1811 84949 1820 84983
rect 1768 84940 1820 84949
rect 4874 84838 4926 84890
rect 4938 84838 4990 84890
rect 5002 84838 5054 84890
rect 5066 84838 5118 84890
rect 5130 84838 5182 84890
rect 106658 84838 106710 84890
rect 106722 84838 106774 84890
rect 106786 84838 106838 84890
rect 106850 84838 106902 84890
rect 106914 84838 106966 84890
rect 1308 84600 1360 84652
rect 1860 84464 1912 84516
rect 4214 84294 4266 84346
rect 4278 84294 4330 84346
rect 4342 84294 4394 84346
rect 4406 84294 4458 84346
rect 4470 84294 4522 84346
rect 105922 84294 105974 84346
rect 105986 84294 106038 84346
rect 106050 84294 106102 84346
rect 106114 84294 106166 84346
rect 106178 84294 106230 84346
rect 1952 84124 2004 84176
rect 9404 84124 9456 84176
rect 1308 83920 1360 83972
rect 8484 83920 8536 83972
rect 4874 83750 4926 83802
rect 4938 83750 4990 83802
rect 5002 83750 5054 83802
rect 5066 83750 5118 83802
rect 5130 83750 5182 83802
rect 106658 83750 106710 83802
rect 106722 83750 106774 83802
rect 106786 83750 106838 83802
rect 106850 83750 106902 83802
rect 106914 83750 106966 83802
rect 1308 83512 1360 83564
rect 2504 83308 2556 83360
rect 4214 83206 4266 83258
rect 4278 83206 4330 83258
rect 4342 83206 4394 83258
rect 4406 83206 4458 83258
rect 4470 83206 4522 83258
rect 105922 83206 105974 83258
rect 105986 83206 106038 83258
rect 106050 83206 106102 83258
rect 106114 83206 106166 83258
rect 106178 83206 106230 83258
rect 1860 82764 1912 82816
rect 9220 82764 9272 82816
rect 4874 82662 4926 82714
rect 4938 82662 4990 82714
rect 5002 82662 5054 82714
rect 5066 82662 5118 82714
rect 5130 82662 5182 82714
rect 106658 82662 106710 82714
rect 106722 82662 106774 82714
rect 106786 82662 106838 82714
rect 106850 82662 106902 82714
rect 106914 82662 106966 82714
rect 1216 82424 1268 82476
rect 2412 82220 2464 82272
rect 4214 82118 4266 82170
rect 4278 82118 4330 82170
rect 4342 82118 4394 82170
rect 4406 82118 4458 82170
rect 4470 82118 4522 82170
rect 105922 82118 105974 82170
rect 105986 82118 106038 82170
rect 106050 82118 106102 82170
rect 106114 82118 106166 82170
rect 106178 82118 106230 82170
rect 1216 81744 1268 81796
rect 1860 81719 1912 81728
rect 1860 81685 1869 81719
rect 1869 81685 1903 81719
rect 1903 81685 1912 81719
rect 1860 81676 1912 81685
rect 4874 81574 4926 81626
rect 4938 81574 4990 81626
rect 5002 81574 5054 81626
rect 5066 81574 5118 81626
rect 5130 81574 5182 81626
rect 106658 81574 106710 81626
rect 106722 81574 106774 81626
rect 106786 81574 106838 81626
rect 106850 81574 106902 81626
rect 106914 81574 106966 81626
rect 1308 81336 1360 81388
rect 1860 81200 1912 81252
rect 9772 81200 9824 81252
rect 5632 81132 5684 81184
rect 4214 81030 4266 81082
rect 4278 81030 4330 81082
rect 4342 81030 4394 81082
rect 4406 81030 4458 81082
rect 4470 81030 4522 81082
rect 105922 81030 105974 81082
rect 105986 81030 106038 81082
rect 106050 81030 106102 81082
rect 106114 81030 106166 81082
rect 106178 81030 106230 81082
rect 2412 80792 2464 80844
rect 9864 80792 9916 80844
rect 1308 80724 1360 80776
rect 2504 80656 2556 80708
rect 9956 80656 10008 80708
rect 5540 80588 5592 80640
rect 4874 80486 4926 80538
rect 4938 80486 4990 80538
rect 5002 80486 5054 80538
rect 5066 80486 5118 80538
rect 5130 80486 5182 80538
rect 106658 80486 106710 80538
rect 106722 80486 106774 80538
rect 106786 80486 106838 80538
rect 106850 80486 106902 80538
rect 106914 80486 106966 80538
rect 1308 80316 1360 80368
rect 4214 79942 4266 79994
rect 4278 79942 4330 79994
rect 4342 79942 4394 79994
rect 4406 79942 4458 79994
rect 4470 79942 4522 79994
rect 9956 79976 10008 80028
rect 40960 79976 41012 80028
rect 9864 79908 9916 79960
rect 39764 79908 39816 79960
rect 105922 79942 105974 79994
rect 105986 79942 106038 79994
rect 106050 79942 106102 79994
rect 106114 79942 106166 79994
rect 106178 79942 106230 79994
rect 9772 79840 9824 79892
rect 38660 79840 38712 79892
rect 8944 79772 8996 79824
rect 36268 79772 36320 79824
rect 8576 79704 8628 79756
rect 34704 79704 34756 79756
rect 9220 79636 9272 79688
rect 32312 79636 32364 79688
rect 1216 79568 1268 79620
rect 37004 79500 37056 79552
rect 4874 79398 4926 79450
rect 4938 79398 4990 79450
rect 5002 79398 5054 79450
rect 5066 79398 5118 79450
rect 5130 79398 5182 79450
rect 106658 79398 106710 79450
rect 106722 79398 106774 79450
rect 106786 79398 106838 79450
rect 106850 79398 106902 79450
rect 106914 79398 106966 79450
rect 61108 79296 61160 79348
rect 101956 79296 102008 79348
rect 1308 79160 1360 79212
rect 42156 78956 42208 79008
rect 88892 78956 88944 79008
rect 108488 78999 108540 79008
rect 108488 78965 108497 78999
rect 108497 78965 108531 78999
rect 108531 78965 108540 78999
rect 108488 78956 108540 78965
rect 4214 78854 4266 78906
rect 4278 78854 4330 78906
rect 4342 78854 4394 78906
rect 4406 78854 4458 78906
rect 4470 78854 4522 78906
rect 105922 78854 105974 78906
rect 105986 78854 106038 78906
rect 106050 78854 106102 78906
rect 106114 78854 106166 78906
rect 106178 78854 106230 78906
rect 96528 78548 96580 78600
rect 102140 78548 102192 78600
rect 1308 78480 1360 78532
rect 79232 78480 79284 78532
rect 91652 78480 91704 78532
rect 29552 78412 29604 78464
rect 76656 78412 76708 78464
rect 89812 78412 89864 78464
rect 108120 78455 108172 78464
rect 108120 78421 108129 78455
rect 108129 78421 108163 78455
rect 108163 78421 108172 78455
rect 108120 78412 108172 78421
rect 108488 78455 108540 78464
rect 108488 78421 108497 78455
rect 108497 78421 108531 78455
rect 108531 78421 108540 78455
rect 108488 78412 108540 78421
rect 4874 78310 4926 78362
rect 4938 78310 4990 78362
rect 5002 78310 5054 78362
rect 5066 78310 5118 78362
rect 5130 78310 5182 78362
rect 71964 78344 72016 78396
rect 85672 78344 85724 78396
rect 22744 78276 22796 78328
rect 22100 78208 22152 78260
rect 2320 78140 2372 78192
rect 1308 78072 1360 78124
rect 25044 78072 25096 78124
rect 73528 78276 73580 78328
rect 80060 78276 80112 78328
rect 106658 78310 106710 78362
rect 106722 78310 106774 78362
rect 106786 78310 106838 78362
rect 106850 78310 106902 78362
rect 106914 78310 106966 78362
rect 26056 78208 26108 78260
rect 30288 78208 30340 78260
rect 69756 78208 69808 78260
rect 102416 78208 102468 78260
rect 34796 78140 34848 78192
rect 63960 78140 64012 78192
rect 81348 78140 81400 78192
rect 20812 78004 20864 78056
rect 27252 78004 27304 78056
rect 21272 77936 21324 77988
rect 30564 77936 30616 77988
rect 31484 78072 31536 78124
rect 33968 78072 34020 78124
rect 63592 78072 63644 78124
rect 71136 78072 71188 78124
rect 74448 78072 74500 78124
rect 88984 78072 89036 78124
rect 30748 78004 30800 78056
rect 39856 78004 39908 78056
rect 58624 78004 58676 78056
rect 43260 77936 43312 77988
rect 43812 77936 43864 77988
rect 53564 77936 53616 77988
rect 62488 77936 62540 77988
rect 31484 77868 31536 77920
rect 31668 77868 31720 77920
rect 36084 77868 36136 77920
rect 56140 77868 56192 77920
rect 64144 77868 64196 77920
rect 69112 78004 69164 78056
rect 85948 78004 86000 78056
rect 87328 78004 87380 78056
rect 102600 78072 102652 78124
rect 93124 78004 93176 78056
rect 107660 78004 107712 78056
rect 66076 77936 66128 77988
rect 73436 77936 73488 77988
rect 80888 77936 80940 77988
rect 94228 77936 94280 77988
rect 67640 77868 67692 77920
rect 70400 77868 70452 77920
rect 87052 77868 87104 77920
rect 90732 77868 90784 77920
rect 99656 77868 99708 77920
rect 105820 77868 105872 77920
rect 108488 77911 108540 77920
rect 108488 77877 108497 77911
rect 108497 77877 108531 77911
rect 108531 77877 108540 77911
rect 108488 77868 108540 77877
rect 4214 77766 4266 77818
rect 4278 77766 4330 77818
rect 4342 77766 4394 77818
rect 4406 77766 4458 77818
rect 4470 77766 4522 77818
rect 34934 77766 34986 77818
rect 34998 77766 35050 77818
rect 35062 77766 35114 77818
rect 35126 77766 35178 77818
rect 35190 77766 35242 77818
rect 65654 77766 65706 77818
rect 65718 77766 65770 77818
rect 65782 77766 65834 77818
rect 65846 77766 65898 77818
rect 65910 77766 65962 77818
rect 96374 77766 96426 77818
rect 96438 77766 96490 77818
rect 96502 77766 96554 77818
rect 96566 77766 96618 77818
rect 96630 77766 96682 77818
rect 105922 77766 105974 77818
rect 105986 77766 106038 77818
rect 106050 77766 106102 77818
rect 106114 77766 106166 77818
rect 106178 77766 106230 77818
rect 17868 77596 17920 77648
rect 21548 77571 21600 77580
rect 6828 77324 6880 77376
rect 16028 77324 16080 77376
rect 21548 77537 21557 77571
rect 21557 77537 21591 77571
rect 21591 77537 21600 77571
rect 21548 77528 21600 77537
rect 22744 77571 22796 77580
rect 22744 77537 22753 77571
rect 22753 77537 22787 77571
rect 22787 77537 22796 77571
rect 22744 77528 22796 77537
rect 27528 77664 27580 77716
rect 27620 77707 27672 77716
rect 27620 77673 27629 77707
rect 27629 77673 27663 77707
rect 27663 77673 27672 77707
rect 27620 77664 27672 77673
rect 28172 77707 28224 77716
rect 28172 77673 28181 77707
rect 28181 77673 28215 77707
rect 28215 77673 28224 77707
rect 28172 77664 28224 77673
rect 29552 77707 29604 77716
rect 29552 77673 29561 77707
rect 29561 77673 29595 77707
rect 29595 77673 29604 77707
rect 29552 77664 29604 77673
rect 30472 77707 30524 77716
rect 30472 77673 30481 77707
rect 30481 77673 30515 77707
rect 30515 77673 30524 77707
rect 30472 77664 30524 77673
rect 30564 77664 30616 77716
rect 31668 77707 31720 77716
rect 31668 77673 31677 77707
rect 31677 77673 31711 77707
rect 31711 77673 31720 77707
rect 31668 77664 31720 77673
rect 32312 77664 32364 77716
rect 32956 77664 33008 77716
rect 33968 77707 34020 77716
rect 33968 77673 33977 77707
rect 33977 77673 34011 77707
rect 34011 77673 34020 77707
rect 33968 77664 34020 77673
rect 34704 77707 34756 77716
rect 34704 77673 34713 77707
rect 34713 77673 34747 77707
rect 34747 77673 34756 77707
rect 34704 77664 34756 77673
rect 34796 77664 34848 77716
rect 35256 77664 35308 77716
rect 40684 77664 40736 77716
rect 24676 77639 24728 77648
rect 24676 77605 24685 77639
rect 24685 77605 24719 77639
rect 24719 77605 24728 77639
rect 24676 77596 24728 77605
rect 24768 77596 24820 77648
rect 25044 77639 25096 77648
rect 25044 77605 25053 77639
rect 25053 77605 25087 77639
rect 25087 77605 25096 77639
rect 25044 77596 25096 77605
rect 26792 77596 26844 77648
rect 20812 77392 20864 77444
rect 21272 77435 21324 77444
rect 21272 77401 21281 77435
rect 21281 77401 21315 77435
rect 21315 77401 21324 77435
rect 21272 77392 21324 77401
rect 21364 77324 21416 77376
rect 26792 77503 26844 77512
rect 26792 77469 26801 77503
rect 26801 77469 26835 77503
rect 26835 77469 26844 77503
rect 31208 77571 31260 77580
rect 31208 77537 31217 77571
rect 31217 77537 31251 77571
rect 31251 77537 31260 77571
rect 31208 77528 31260 77537
rect 32956 77528 33008 77580
rect 38660 77639 38712 77648
rect 38660 77605 38669 77639
rect 38669 77605 38703 77639
rect 38703 77605 38712 77639
rect 38660 77596 38712 77605
rect 39764 77596 39816 77648
rect 39856 77639 39908 77648
rect 39856 77605 39865 77639
rect 39865 77605 39899 77639
rect 39899 77605 39908 77639
rect 39856 77596 39908 77605
rect 40868 77639 40920 77648
rect 40868 77605 40877 77639
rect 40877 77605 40911 77639
rect 40911 77605 40920 77639
rect 40868 77596 40920 77605
rect 40960 77596 41012 77648
rect 42156 77639 42208 77648
rect 42156 77605 42165 77639
rect 42165 77605 42199 77639
rect 42199 77605 42208 77639
rect 42156 77596 42208 77605
rect 62488 77639 62540 77648
rect 62488 77605 62497 77639
rect 62497 77605 62531 77639
rect 62531 77605 62540 77639
rect 62488 77596 62540 77605
rect 43812 77571 43864 77580
rect 43812 77537 43821 77571
rect 43821 77537 43855 77571
rect 43855 77537 43864 77571
rect 43812 77528 43864 77537
rect 63960 77639 64012 77648
rect 63960 77605 63969 77639
rect 63969 77605 64003 77639
rect 64003 77605 64012 77639
rect 63960 77596 64012 77605
rect 64972 77596 65024 77648
rect 64052 77571 64104 77580
rect 64052 77537 64061 77571
rect 64061 77537 64095 77571
rect 64095 77537 64104 77571
rect 64052 77528 64104 77537
rect 64144 77528 64196 77580
rect 67640 77639 67692 77648
rect 67640 77605 67649 77639
rect 67649 77605 67683 77639
rect 67683 77605 67692 77639
rect 67640 77596 67692 77605
rect 26792 77460 26844 77469
rect 35256 77503 35308 77512
rect 35256 77469 35265 77503
rect 35265 77469 35299 77503
rect 35299 77469 35308 77503
rect 35256 77460 35308 77469
rect 35348 77503 35400 77512
rect 35348 77469 35357 77503
rect 35357 77469 35391 77503
rect 35391 77469 35400 77503
rect 35348 77460 35400 77469
rect 36268 77460 36320 77512
rect 37004 77503 37056 77512
rect 37004 77469 37013 77503
rect 37013 77469 37047 77503
rect 37047 77469 37056 77503
rect 37004 77460 37056 77469
rect 40040 77460 40092 77512
rect 26056 77392 26108 77444
rect 39948 77392 40000 77444
rect 46112 77460 46164 77512
rect 61108 77503 61160 77512
rect 61108 77469 61117 77503
rect 61117 77469 61151 77503
rect 61151 77469 61160 77503
rect 61108 77460 61160 77469
rect 63316 77503 63368 77512
rect 63316 77469 63325 77503
rect 63325 77469 63359 77503
rect 63359 77469 63368 77503
rect 63316 77460 63368 77469
rect 48596 77392 48648 77444
rect 51080 77392 51132 77444
rect 62488 77392 62540 77444
rect 31576 77324 31628 77376
rect 32680 77367 32732 77376
rect 32680 77333 32689 77367
rect 32689 77333 32723 77367
rect 32723 77333 32732 77367
rect 32680 77324 32732 77333
rect 35992 77324 36044 77376
rect 37280 77367 37332 77376
rect 37280 77333 37289 77367
rect 37289 77333 37323 77367
rect 37323 77333 37332 77367
rect 37280 77324 37332 77333
rect 37740 77367 37792 77376
rect 37740 77333 37749 77367
rect 37749 77333 37783 77367
rect 37783 77333 37792 77367
rect 37740 77324 37792 77333
rect 40132 77324 40184 77376
rect 42432 77367 42484 77376
rect 42432 77333 42441 77367
rect 42441 77333 42475 77367
rect 42475 77333 42484 77367
rect 42432 77324 42484 77333
rect 42892 77367 42944 77376
rect 42892 77333 42901 77367
rect 42901 77333 42935 77367
rect 42935 77333 42944 77367
rect 42892 77324 42944 77333
rect 64052 77324 64104 77376
rect 64972 77324 65024 77376
rect 68284 77571 68336 77580
rect 68284 77537 68293 77571
rect 68293 77537 68327 77571
rect 68327 77537 68336 77571
rect 68284 77528 68336 77537
rect 68468 77571 68520 77580
rect 68468 77537 68477 77571
rect 68477 77537 68511 77571
rect 68511 77537 68520 77571
rect 68468 77528 68520 77537
rect 65892 77503 65944 77512
rect 65892 77469 65901 77503
rect 65901 77469 65935 77503
rect 65935 77469 65944 77503
rect 65892 77460 65944 77469
rect 67364 77460 67416 77512
rect 69112 77639 69164 77648
rect 69112 77605 69121 77639
rect 69121 77605 69155 77639
rect 69155 77605 69164 77639
rect 69112 77596 69164 77605
rect 69204 77528 69256 77580
rect 70400 77707 70452 77716
rect 70400 77673 70409 77707
rect 70409 77673 70443 77707
rect 70443 77673 70452 77707
rect 70400 77664 70452 77673
rect 70952 77707 71004 77716
rect 70952 77673 70961 77707
rect 70961 77673 70995 77707
rect 70995 77673 71004 77707
rect 70952 77664 71004 77673
rect 71044 77664 71096 77716
rect 69756 77571 69808 77580
rect 69756 77537 69765 77571
rect 69765 77537 69799 77571
rect 69799 77537 69808 77571
rect 69756 77528 69808 77537
rect 71136 77639 71188 77648
rect 71136 77605 71145 77639
rect 71145 77605 71179 77639
rect 71179 77605 71188 77639
rect 71136 77596 71188 77605
rect 71964 77707 72016 77716
rect 71964 77673 71973 77707
rect 71973 77673 72007 77707
rect 72007 77673 72016 77707
rect 71964 77664 72016 77673
rect 74448 77707 74500 77716
rect 74448 77673 74457 77707
rect 74457 77673 74491 77707
rect 74491 77673 74500 77707
rect 74448 77664 74500 77673
rect 76656 77707 76708 77716
rect 76656 77673 76665 77707
rect 76665 77673 76699 77707
rect 76699 77673 76708 77707
rect 76656 77664 76708 77673
rect 78772 77664 78824 77716
rect 79232 77707 79284 77716
rect 79232 77673 79241 77707
rect 79241 77673 79275 77707
rect 79275 77673 79284 77707
rect 79232 77664 79284 77673
rect 80060 77707 80112 77716
rect 80060 77673 80069 77707
rect 80069 77673 80103 77707
rect 80103 77673 80112 77707
rect 80060 77664 80112 77673
rect 73804 77571 73856 77580
rect 73804 77537 73813 77571
rect 73813 77537 73847 77571
rect 73847 77537 73856 77571
rect 73804 77528 73856 77537
rect 73988 77571 74040 77580
rect 73988 77537 73997 77571
rect 73997 77537 74031 77571
rect 74031 77537 74040 77571
rect 73988 77528 74040 77537
rect 74632 77503 74684 77512
rect 74632 77469 74641 77503
rect 74641 77469 74675 77503
rect 74675 77469 74684 77503
rect 74632 77460 74684 77469
rect 71320 77392 71372 77444
rect 68284 77324 68336 77376
rect 69204 77324 69256 77376
rect 69756 77324 69808 77376
rect 69848 77367 69900 77376
rect 69848 77333 69857 77367
rect 69857 77333 69891 77367
rect 69891 77333 69900 77367
rect 69848 77324 69900 77333
rect 71136 77324 71188 77376
rect 73436 77392 73488 77444
rect 71688 77324 71740 77376
rect 73804 77324 73856 77376
rect 76196 77571 76248 77580
rect 76196 77537 76205 77571
rect 76205 77537 76239 77571
rect 76239 77537 76248 77571
rect 76196 77528 76248 77537
rect 78772 77571 78824 77580
rect 78772 77537 78781 77571
rect 78781 77537 78815 77571
rect 78815 77537 78824 77571
rect 78772 77528 78824 77537
rect 80888 77639 80940 77648
rect 80888 77605 80897 77639
rect 80897 77605 80931 77639
rect 80931 77605 80940 77639
rect 80888 77596 80940 77605
rect 103796 77664 103848 77716
rect 86592 77596 86644 77648
rect 87328 77639 87380 77648
rect 87328 77605 87337 77639
rect 87337 77605 87371 77639
rect 87371 77605 87380 77639
rect 87328 77596 87380 77605
rect 90732 77639 90784 77648
rect 90732 77605 90741 77639
rect 90741 77605 90775 77639
rect 90775 77605 90784 77639
rect 90732 77596 90784 77605
rect 93124 77639 93176 77648
rect 93124 77605 93133 77639
rect 93133 77605 93167 77639
rect 93167 77605 93176 77639
rect 93124 77596 93176 77605
rect 86500 77571 86552 77580
rect 86500 77537 86509 77571
rect 86509 77537 86543 77571
rect 86543 77537 86552 77571
rect 86500 77528 86552 77537
rect 89076 77528 89128 77580
rect 80060 77460 80112 77512
rect 81532 77392 81584 77444
rect 83096 77435 83148 77444
rect 83096 77401 83105 77435
rect 83105 77401 83139 77435
rect 83139 77401 83148 77435
rect 83096 77392 83148 77401
rect 83832 77503 83884 77512
rect 83832 77469 83841 77503
rect 83841 77469 83875 77503
rect 83875 77469 83884 77503
rect 83832 77460 83884 77469
rect 84292 77392 84344 77444
rect 86408 77460 86460 77512
rect 86868 77460 86920 77512
rect 75644 77324 75696 77376
rect 76196 77324 76248 77376
rect 76288 77367 76340 77376
rect 76288 77333 76297 77367
rect 76297 77333 76331 77367
rect 76331 77333 76340 77367
rect 76288 77324 76340 77333
rect 83648 77367 83700 77376
rect 83648 77333 83657 77367
rect 83657 77333 83691 77367
rect 83691 77333 83700 77367
rect 83648 77324 83700 77333
rect 84016 77367 84068 77376
rect 84016 77333 84025 77367
rect 84025 77333 84059 77367
rect 84059 77333 84068 77367
rect 84016 77324 84068 77333
rect 86500 77324 86552 77376
rect 87236 77392 87288 77444
rect 88984 77392 89036 77444
rect 89720 77392 89772 77444
rect 89444 77324 89496 77376
rect 91652 77435 91704 77444
rect 91652 77401 91661 77435
rect 91661 77401 91695 77435
rect 91695 77401 91704 77435
rect 91652 77392 91704 77401
rect 92664 77392 92716 77444
rect 92020 77324 92072 77376
rect 94228 77435 94280 77444
rect 94228 77401 94237 77435
rect 94237 77401 94271 77435
rect 94271 77401 94280 77435
rect 94228 77392 94280 77401
rect 95240 77392 95292 77444
rect 99656 77528 99708 77580
rect 108120 77528 108172 77580
rect 106280 77392 106332 77444
rect 104164 77324 104216 77376
rect 4874 77222 4926 77274
rect 4938 77222 4990 77274
rect 5002 77222 5054 77274
rect 5066 77222 5118 77274
rect 5130 77222 5182 77274
rect 35594 77222 35646 77274
rect 35658 77222 35710 77274
rect 35722 77222 35774 77274
rect 35786 77222 35838 77274
rect 35850 77222 35902 77274
rect 66314 77222 66366 77274
rect 66378 77222 66430 77274
rect 66442 77222 66494 77274
rect 66506 77222 66558 77274
rect 66570 77222 66622 77274
rect 97034 77222 97086 77274
rect 97098 77222 97150 77274
rect 97162 77222 97214 77274
rect 97226 77222 97278 77274
rect 97290 77222 97342 77274
rect 106658 77222 106710 77274
rect 106722 77222 106774 77274
rect 106786 77222 106838 77274
rect 106850 77222 106902 77274
rect 106914 77222 106966 77274
rect 1768 77120 1820 77172
rect 23480 77120 23532 77172
rect 27252 77120 27304 77172
rect 68560 77120 68612 77172
rect 76288 77120 76340 77172
rect 81532 77163 81584 77172
rect 81532 77129 81541 77163
rect 81541 77129 81575 77163
rect 81575 77129 81584 77163
rect 81532 77120 81584 77129
rect 83096 77120 83148 77172
rect 24768 77052 24820 77104
rect 27436 77052 27488 77104
rect 27528 77052 27580 77104
rect 69204 77095 69256 77104
rect 69204 77061 69213 77095
rect 69213 77061 69247 77095
rect 69247 77061 69256 77095
rect 69204 77052 69256 77061
rect 75644 77095 75696 77104
rect 75644 77061 75653 77095
rect 75653 77061 75687 77095
rect 75687 77061 75696 77095
rect 75644 77052 75696 77061
rect 1216 76984 1268 77036
rect 26792 76984 26844 77036
rect 24308 76959 24360 76968
rect 24308 76925 24317 76959
rect 24317 76925 24351 76959
rect 24351 76925 24360 76959
rect 24308 76916 24360 76925
rect 24584 76959 24636 76968
rect 24584 76925 24593 76959
rect 24593 76925 24627 76959
rect 24627 76925 24636 76959
rect 24584 76916 24636 76925
rect 30472 76916 30524 76968
rect 22008 76848 22060 76900
rect 22100 76780 22152 76832
rect 22836 76823 22888 76832
rect 22836 76789 22845 76823
rect 22845 76789 22879 76823
rect 22879 76789 22888 76823
rect 22836 76780 22888 76789
rect 26792 76823 26844 76832
rect 26792 76789 26801 76823
rect 26801 76789 26835 76823
rect 26835 76789 26844 76823
rect 26792 76780 26844 76789
rect 30564 76823 30616 76832
rect 30564 76789 30573 76823
rect 30573 76789 30607 76823
rect 30607 76789 30616 76823
rect 30564 76780 30616 76789
rect 61108 76780 61160 76832
rect 69848 76848 69900 76900
rect 83832 76984 83884 77036
rect 83924 76916 83976 76968
rect 88432 77120 88484 77172
rect 88892 77163 88944 77172
rect 88892 77129 88901 77163
rect 88901 77129 88935 77163
rect 88935 77129 88944 77163
rect 88892 77120 88944 77129
rect 92020 77163 92072 77172
rect 92020 77129 92029 77163
rect 92029 77129 92063 77163
rect 92063 77129 92072 77163
rect 92020 77120 92072 77129
rect 85764 77052 85816 77104
rect 88524 77052 88576 77104
rect 95240 77052 95292 77104
rect 85580 76984 85632 77036
rect 86408 76984 86460 77036
rect 86500 76984 86552 77036
rect 86868 77027 86920 77036
rect 86868 76993 86877 77027
rect 86877 76993 86911 77027
rect 86911 76993 86920 77027
rect 86868 76984 86920 76993
rect 88984 76984 89036 77036
rect 89444 77027 89496 77036
rect 89444 76993 89453 77027
rect 89453 76993 89487 77027
rect 89487 76993 89496 77027
rect 89444 76984 89496 76993
rect 91468 76984 91520 77036
rect 106280 76984 106332 77036
rect 85672 76916 85724 76968
rect 89812 76916 89864 76968
rect 82820 76780 82872 76832
rect 84016 76780 84068 76832
rect 86776 76848 86828 76900
rect 105820 76848 105872 76900
rect 108488 76891 108540 76900
rect 108488 76857 108497 76891
rect 108497 76857 108531 76891
rect 108531 76857 108540 76891
rect 108488 76848 108540 76857
rect 85580 76780 85632 76832
rect 86132 76823 86184 76832
rect 86132 76789 86141 76823
rect 86141 76789 86175 76823
rect 86175 76789 86184 76823
rect 86132 76780 86184 76789
rect 86592 76780 86644 76832
rect 87236 76780 87288 76832
rect 89904 76780 89956 76832
rect 91468 76823 91520 76832
rect 91468 76789 91477 76823
rect 91477 76789 91511 76823
rect 91511 76789 91520 76823
rect 91468 76780 91520 76789
rect 4214 76678 4266 76730
rect 4278 76678 4330 76730
rect 4342 76678 4394 76730
rect 4406 76678 4458 76730
rect 4470 76678 4522 76730
rect 34934 76678 34986 76730
rect 34998 76678 35050 76730
rect 35062 76678 35114 76730
rect 35126 76678 35178 76730
rect 35190 76678 35242 76730
rect 65654 76678 65706 76730
rect 65718 76678 65770 76730
rect 65782 76678 65834 76730
rect 65846 76678 65898 76730
rect 65910 76678 65962 76730
rect 96374 76678 96426 76730
rect 96438 76678 96490 76730
rect 96502 76678 96554 76730
rect 96566 76678 96618 76730
rect 96630 76678 96682 76730
rect 21548 76619 21600 76628
rect 21548 76585 21557 76619
rect 21557 76585 21591 76619
rect 21591 76585 21600 76619
rect 21548 76576 21600 76585
rect 23480 76619 23532 76628
rect 23480 76585 23489 76619
rect 23489 76585 23523 76619
rect 23523 76585 23532 76619
rect 23480 76576 23532 76585
rect 24584 76576 24636 76628
rect 26792 76576 26844 76628
rect 27436 76576 27488 76628
rect 84292 76576 84344 76628
rect 85764 76619 85816 76628
rect 85764 76585 85773 76619
rect 85773 76585 85807 76619
rect 85807 76585 85816 76619
rect 85764 76576 85816 76585
rect 85948 76619 86000 76628
rect 85948 76585 85957 76619
rect 85957 76585 85991 76619
rect 85991 76585 86000 76619
rect 85948 76576 86000 76585
rect 86132 76576 86184 76628
rect 23020 76508 23072 76560
rect 24768 76508 24820 76560
rect 32680 76440 32732 76492
rect 83648 76440 83700 76492
rect 86868 76440 86920 76492
rect 88524 76619 88576 76628
rect 88524 76585 88533 76619
rect 88533 76585 88567 76619
rect 88567 76585 88576 76619
rect 88524 76576 88576 76585
rect 88984 76619 89036 76628
rect 88984 76585 88993 76619
rect 88993 76585 89027 76619
rect 89027 76585 89036 76619
rect 88984 76576 89036 76585
rect 92664 76576 92716 76628
rect 89720 76508 89772 76560
rect 102232 76440 102284 76492
rect 17868 76372 17920 76424
rect 30564 76372 30616 76424
rect 30288 76304 30340 76356
rect 848 76236 900 76288
rect 82820 76372 82872 76424
rect 73988 76236 74040 76288
rect 83280 76347 83332 76356
rect 83280 76313 83289 76347
rect 83289 76313 83323 76347
rect 83323 76313 83332 76347
rect 83280 76304 83332 76313
rect 85580 76236 85632 76288
rect 86408 76304 86460 76356
rect 86960 76304 87012 76356
rect 87144 76236 87196 76288
rect 88432 76415 88484 76424
rect 88432 76381 88441 76415
rect 88441 76381 88475 76415
rect 88475 76381 88484 76415
rect 88432 76372 88484 76381
rect 89168 76372 89220 76424
rect 89720 76415 89772 76424
rect 89720 76381 89729 76415
rect 89729 76381 89763 76415
rect 89763 76381 89772 76415
rect 89720 76372 89772 76381
rect 107660 76372 107712 76424
rect 108120 76304 108172 76356
rect 89168 76279 89220 76288
rect 89168 76245 89177 76279
rect 89177 76245 89211 76279
rect 89211 76245 89220 76279
rect 89168 76236 89220 76245
rect 89720 76236 89772 76288
rect 91468 76236 91520 76288
rect 108488 76279 108540 76288
rect 108488 76245 108497 76279
rect 108497 76245 108531 76279
rect 108531 76245 108540 76279
rect 108488 76236 108540 76245
rect 4874 76134 4926 76186
rect 4938 76134 4990 76186
rect 5002 76134 5054 76186
rect 5066 76134 5118 76186
rect 5130 76134 5182 76186
rect 35594 76134 35646 76186
rect 35658 76134 35710 76186
rect 35722 76134 35774 76186
rect 35786 76134 35838 76186
rect 35850 76134 35902 76186
rect 66314 76134 66366 76186
rect 66378 76134 66430 76186
rect 66442 76134 66494 76186
rect 66506 76134 66558 76186
rect 66570 76134 66622 76186
rect 97034 76134 97086 76186
rect 97098 76134 97150 76186
rect 97162 76134 97214 76186
rect 97226 76134 97278 76186
rect 97290 76134 97342 76186
rect 2320 76032 2372 76084
rect 82820 76032 82872 76084
rect 83924 76075 83976 76084
rect 24308 75964 24360 76016
rect 37280 75964 37332 76016
rect 81348 75964 81400 76016
rect 83280 75964 83332 76016
rect 83924 76041 83933 76075
rect 83933 76041 83967 76075
rect 83967 76041 83976 76075
rect 83924 76032 83976 76041
rect 84292 76032 84344 76084
rect 86684 76032 86736 76084
rect 86776 76032 86828 76084
rect 87236 75964 87288 76016
rect 87420 75964 87472 76016
rect 84292 75939 84344 75948
rect 84292 75905 84301 75939
rect 84301 75905 84335 75939
rect 84335 75905 84344 75939
rect 84292 75896 84344 75905
rect 89904 75896 89956 75948
rect 108120 76075 108172 76084
rect 108120 76041 108129 76075
rect 108129 76041 108163 76075
rect 108163 76041 108172 76075
rect 108120 76032 108172 76041
rect 108488 76075 108540 76084
rect 108488 76041 108497 76075
rect 108497 76041 108531 76075
rect 108531 76041 108540 76075
rect 108488 76032 108540 76041
rect 90732 75896 90784 75948
rect 71780 75828 71832 75880
rect 86684 75871 86736 75880
rect 86684 75837 86693 75871
rect 86693 75837 86727 75871
rect 86727 75837 86736 75871
rect 86684 75828 86736 75837
rect 87052 75828 87104 75880
rect 88708 75828 88760 75880
rect 89076 75828 89128 75880
rect 86592 75760 86644 75812
rect 1400 75735 1452 75744
rect 1400 75701 1409 75735
rect 1409 75701 1443 75735
rect 1443 75701 1452 75735
rect 1400 75692 1452 75701
rect 86316 75735 86368 75744
rect 86316 75701 86325 75735
rect 86325 75701 86359 75735
rect 86359 75701 86368 75735
rect 86316 75692 86368 75701
rect 90180 75692 90232 75744
rect 90456 75692 90508 75744
rect 102692 75760 102744 75812
rect 108120 75692 108172 75744
rect 4214 75590 4266 75642
rect 4278 75590 4330 75642
rect 4342 75590 4394 75642
rect 4406 75590 4458 75642
rect 4470 75590 4522 75642
rect 34934 75590 34986 75642
rect 34998 75590 35050 75642
rect 35062 75590 35114 75642
rect 35126 75590 35178 75642
rect 35190 75590 35242 75642
rect 65654 75590 65706 75642
rect 65718 75590 65770 75642
rect 65782 75590 65834 75642
rect 65846 75590 65898 75642
rect 65910 75590 65962 75642
rect 96374 75590 96426 75642
rect 96438 75590 96490 75642
rect 96502 75590 96554 75642
rect 96566 75590 96618 75642
rect 96630 75590 96682 75642
rect 86684 75488 86736 75540
rect 88708 75488 88760 75540
rect 89904 75488 89956 75540
rect 90364 75488 90416 75540
rect 87420 75420 87472 75472
rect 848 75148 900 75200
rect 67364 75216 67416 75268
rect 86960 75352 87012 75404
rect 82176 75327 82228 75336
rect 82176 75293 82185 75327
rect 82185 75293 82219 75327
rect 82219 75293 82228 75327
rect 82176 75284 82228 75293
rect 86592 75327 86644 75336
rect 86592 75293 86601 75327
rect 86601 75293 86635 75327
rect 86635 75293 86644 75327
rect 86592 75284 86644 75293
rect 90456 75284 90508 75336
rect 22008 75148 22060 75200
rect 82084 75191 82136 75200
rect 82084 75157 82093 75191
rect 82093 75157 82127 75191
rect 82127 75157 82136 75191
rect 82084 75148 82136 75157
rect 87144 75216 87196 75268
rect 90824 75259 90876 75268
rect 90824 75225 90833 75259
rect 90833 75225 90867 75259
rect 90867 75225 90876 75259
rect 90824 75216 90876 75225
rect 84384 75191 84436 75200
rect 84384 75157 84393 75191
rect 84393 75157 84427 75191
rect 84427 75157 84436 75191
rect 84384 75148 84436 75157
rect 87052 75148 87104 75200
rect 90456 75191 90508 75200
rect 90456 75157 90465 75191
rect 90465 75157 90499 75191
rect 90499 75157 90508 75191
rect 90456 75148 90508 75157
rect 90732 75148 90784 75200
rect 108488 75191 108540 75200
rect 108488 75157 108497 75191
rect 108497 75157 108531 75191
rect 108531 75157 108540 75191
rect 108488 75148 108540 75157
rect 4874 75046 4926 75098
rect 4938 75046 4990 75098
rect 5002 75046 5054 75098
rect 5066 75046 5118 75098
rect 5130 75046 5182 75098
rect 35594 75046 35646 75098
rect 35658 75046 35710 75098
rect 35722 75046 35774 75098
rect 35786 75046 35838 75098
rect 35850 75046 35902 75098
rect 66314 75046 66366 75098
rect 66378 75046 66430 75098
rect 66442 75046 66494 75098
rect 66506 75046 66558 75098
rect 66570 75046 66622 75098
rect 97034 75046 97086 75098
rect 97098 75046 97150 75098
rect 97162 75046 97214 75098
rect 97226 75046 97278 75098
rect 97290 75046 97342 75098
rect 82176 74944 82228 74996
rect 82820 74944 82872 74996
rect 84384 74944 84436 74996
rect 102140 74944 102192 74996
rect 4214 74502 4266 74554
rect 4278 74502 4330 74554
rect 4342 74502 4394 74554
rect 4406 74502 4458 74554
rect 4470 74502 4522 74554
rect 34934 74502 34986 74554
rect 34998 74502 35050 74554
rect 35062 74502 35114 74554
rect 35126 74502 35178 74554
rect 35190 74502 35242 74554
rect 65654 74502 65706 74554
rect 65718 74502 65770 74554
rect 65782 74502 65834 74554
rect 65846 74502 65898 74554
rect 65910 74502 65962 74554
rect 96374 74502 96426 74554
rect 96438 74502 96490 74554
rect 96502 74502 96554 74554
rect 96566 74502 96618 74554
rect 96630 74502 96682 74554
rect 848 74332 900 74384
rect 22836 74196 22888 74248
rect 85580 74196 85632 74248
rect 108488 74103 108540 74112
rect 108488 74069 108497 74103
rect 108497 74069 108531 74103
rect 108531 74069 108540 74103
rect 108488 74060 108540 74069
rect 4874 73958 4926 74010
rect 4938 73958 4990 74010
rect 5002 73958 5054 74010
rect 5066 73958 5118 74010
rect 5130 73958 5182 74010
rect 35594 73958 35646 74010
rect 35658 73958 35710 74010
rect 35722 73958 35774 74010
rect 35786 73958 35838 74010
rect 35850 73958 35902 74010
rect 66314 73958 66366 74010
rect 66378 73958 66430 74010
rect 66442 73958 66494 74010
rect 66506 73958 66558 74010
rect 66570 73958 66622 74010
rect 97034 73958 97086 74010
rect 97098 73958 97150 74010
rect 97162 73958 97214 74010
rect 97226 73958 97278 74010
rect 97290 73958 97342 74010
rect 21364 73720 21416 73772
rect 848 73584 900 73636
rect 102140 73516 102192 73568
rect 108488 73559 108540 73568
rect 108488 73525 108497 73559
rect 108497 73525 108531 73559
rect 108531 73525 108540 73559
rect 108488 73516 108540 73525
rect 4214 73414 4266 73466
rect 4278 73414 4330 73466
rect 4342 73414 4394 73466
rect 4406 73414 4458 73466
rect 4470 73414 4522 73466
rect 34934 73414 34986 73466
rect 34998 73414 35050 73466
rect 35062 73414 35114 73466
rect 35126 73414 35178 73466
rect 35190 73414 35242 73466
rect 65654 73414 65706 73466
rect 65718 73414 65770 73466
rect 65782 73414 65834 73466
rect 65846 73414 65898 73466
rect 65910 73414 65962 73466
rect 96374 73414 96426 73466
rect 96438 73414 96490 73466
rect 96502 73414 96554 73466
rect 96566 73414 96618 73466
rect 96630 73414 96682 73466
rect 1768 73355 1820 73364
rect 1768 73321 1777 73355
rect 1777 73321 1811 73355
rect 1811 73321 1820 73355
rect 1768 73312 1820 73321
rect 108120 73355 108172 73364
rect 108120 73321 108129 73355
rect 108129 73321 108163 73355
rect 108163 73321 108172 73355
rect 108120 73312 108172 73321
rect 88984 73244 89036 73296
rect 90272 73244 90324 73296
rect 90640 73244 90692 73296
rect 1768 73108 1820 73160
rect 90180 73108 90232 73160
rect 90456 73108 90508 73160
rect 90640 73108 90692 73160
rect 108120 73108 108172 73160
rect 848 72972 900 73024
rect 108488 73015 108540 73024
rect 108488 72981 108497 73015
rect 108497 72981 108531 73015
rect 108531 72981 108540 73015
rect 108488 72972 108540 72981
rect 4874 72870 4926 72922
rect 4938 72870 4990 72922
rect 5002 72870 5054 72922
rect 5066 72870 5118 72922
rect 5130 72870 5182 72922
rect 35594 72870 35646 72922
rect 35658 72870 35710 72922
rect 35722 72870 35774 72922
rect 35786 72870 35838 72922
rect 35850 72870 35902 72922
rect 66314 72870 66366 72922
rect 66378 72870 66430 72922
rect 66442 72870 66494 72922
rect 66506 72870 66558 72922
rect 66570 72870 66622 72922
rect 97034 72870 97086 72922
rect 97098 72870 97150 72922
rect 97162 72870 97214 72922
rect 97226 72870 97278 72922
rect 97290 72870 97342 72922
rect 1124 72632 1176 72684
rect 7288 72632 7340 72684
rect 26792 72700 26844 72752
rect 44180 72675 44232 72684
rect 44180 72641 44189 72675
rect 44189 72641 44223 72675
rect 44223 72641 44232 72675
rect 74080 72700 74132 72752
rect 77208 72700 77260 72752
rect 44180 72632 44232 72641
rect 28172 72428 28224 72480
rect 75092 72564 75144 72616
rect 57796 72496 57848 72548
rect 82084 72564 82136 72616
rect 95148 72428 95200 72480
rect 104348 72428 104400 72480
rect 4214 72326 4266 72378
rect 4278 72326 4330 72378
rect 4342 72326 4394 72378
rect 4406 72326 4458 72378
rect 4470 72326 4522 72378
rect 34934 72326 34986 72378
rect 34998 72326 35050 72378
rect 35062 72326 35114 72378
rect 35126 72326 35178 72378
rect 35190 72326 35242 72378
rect 65654 72326 65706 72378
rect 65718 72326 65770 72378
rect 65782 72326 65834 72378
rect 65846 72326 65898 72378
rect 65910 72326 65962 72378
rect 96374 72326 96426 72378
rect 96438 72326 96490 72378
rect 96502 72326 96554 72378
rect 96566 72326 96618 72378
rect 96630 72326 96682 72378
rect 44180 72224 44232 72276
rect 74080 72224 74132 72276
rect 73988 72020 74040 72072
rect 74356 72020 74408 72072
rect 9588 71952 9640 72004
rect 57796 71995 57848 72004
rect 57796 71961 57805 71995
rect 57805 71961 57839 71995
rect 57839 71961 57848 71995
rect 57796 71952 57848 71961
rect 74356 71927 74408 71936
rect 74356 71893 74365 71927
rect 74365 71893 74399 71927
rect 74399 71893 74408 71927
rect 74356 71884 74408 71893
rect 94320 72224 94372 72276
rect 95148 72224 95200 72276
rect 90824 72020 90876 72072
rect 90364 71952 90416 72004
rect 92388 71952 92440 72004
rect 102876 71952 102928 72004
rect 87696 71884 87748 71936
rect 91836 71927 91888 71936
rect 91836 71893 91845 71927
rect 91845 71893 91879 71927
rect 91879 71893 91888 71927
rect 91836 71884 91888 71893
rect 92112 71927 92164 71936
rect 92112 71893 92121 71927
rect 92121 71893 92155 71927
rect 92155 71893 92164 71927
rect 92112 71884 92164 71893
rect 4874 71782 4926 71834
rect 4938 71782 4990 71834
rect 5002 71782 5054 71834
rect 5066 71782 5118 71834
rect 5130 71782 5182 71834
rect 35594 71782 35646 71834
rect 35658 71782 35710 71834
rect 35722 71782 35774 71834
rect 35786 71782 35838 71834
rect 35850 71782 35902 71834
rect 66314 71782 66366 71834
rect 66378 71782 66430 71834
rect 66442 71782 66494 71834
rect 66506 71782 66558 71834
rect 66570 71782 66622 71834
rect 97034 71782 97086 71834
rect 97098 71782 97150 71834
rect 97162 71782 97214 71834
rect 97226 71782 97278 71834
rect 97290 71782 97342 71834
rect 90732 71723 90784 71732
rect 90732 71689 90741 71723
rect 90741 71689 90775 71723
rect 90775 71689 90784 71723
rect 90732 71680 90784 71689
rect 91100 71544 91152 71596
rect 91836 71587 91888 71596
rect 91836 71553 91845 71587
rect 91845 71553 91879 71587
rect 91879 71553 91888 71587
rect 91836 71544 91888 71553
rect 102232 71340 102284 71392
rect 4214 71238 4266 71290
rect 4278 71238 4330 71290
rect 4342 71238 4394 71290
rect 4406 71238 4458 71290
rect 4470 71238 4522 71290
rect 34934 71238 34986 71290
rect 34998 71238 35050 71290
rect 35062 71238 35114 71290
rect 35126 71238 35178 71290
rect 35190 71238 35242 71290
rect 65654 71238 65706 71290
rect 65718 71238 65770 71290
rect 65782 71238 65834 71290
rect 65846 71238 65898 71290
rect 65910 71238 65962 71290
rect 96374 71238 96426 71290
rect 96438 71238 96490 71290
rect 96502 71238 96554 71290
rect 96566 71238 96618 71290
rect 96630 71238 96682 71290
rect 91100 71136 91152 71188
rect 74632 71000 74684 71052
rect 78036 71000 78088 71052
rect 88708 71043 88760 71052
rect 88708 71009 88717 71043
rect 88717 71009 88751 71043
rect 88751 71009 88760 71043
rect 88708 71000 88760 71009
rect 75092 70932 75144 70984
rect 87144 70932 87196 70984
rect 87880 70975 87932 70984
rect 87880 70941 87889 70975
rect 87889 70941 87923 70975
rect 87923 70941 87932 70975
rect 87880 70932 87932 70941
rect 88984 70907 89036 70916
rect 88984 70873 88993 70907
rect 88993 70873 89027 70907
rect 89027 70873 89036 70907
rect 88984 70864 89036 70873
rect 4874 70694 4926 70746
rect 4938 70694 4990 70746
rect 5002 70694 5054 70746
rect 5066 70694 5118 70746
rect 5130 70694 5182 70746
rect 35594 70694 35646 70746
rect 35658 70694 35710 70746
rect 35722 70694 35774 70746
rect 35786 70694 35838 70746
rect 35850 70694 35902 70746
rect 66314 70694 66366 70746
rect 66378 70694 66430 70746
rect 66442 70694 66494 70746
rect 66506 70694 66558 70746
rect 66570 70694 66622 70746
rect 97034 70694 97086 70746
rect 97098 70694 97150 70746
rect 97162 70694 97214 70746
rect 97226 70694 97278 70746
rect 97290 70694 97342 70746
rect 78036 70635 78088 70644
rect 78036 70601 78045 70635
rect 78045 70601 78079 70635
rect 78079 70601 78088 70635
rect 78036 70592 78088 70601
rect 77208 70388 77260 70440
rect 85672 70388 85724 70440
rect 4214 70150 4266 70202
rect 4278 70150 4330 70202
rect 4342 70150 4394 70202
rect 4406 70150 4458 70202
rect 4470 70150 4522 70202
rect 34934 70150 34986 70202
rect 34998 70150 35050 70202
rect 35062 70150 35114 70202
rect 35126 70150 35178 70202
rect 35190 70150 35242 70202
rect 65654 70150 65706 70202
rect 65718 70150 65770 70202
rect 65782 70150 65834 70202
rect 65846 70150 65898 70202
rect 65910 70150 65962 70202
rect 96374 70150 96426 70202
rect 96438 70150 96490 70202
rect 96502 70150 96554 70202
rect 96566 70150 96618 70202
rect 96630 70150 96682 70202
rect 4874 69606 4926 69658
rect 4938 69606 4990 69658
rect 5002 69606 5054 69658
rect 5066 69606 5118 69658
rect 5130 69606 5182 69658
rect 35594 69606 35646 69658
rect 35658 69606 35710 69658
rect 35722 69606 35774 69658
rect 35786 69606 35838 69658
rect 35850 69606 35902 69658
rect 66314 69606 66366 69658
rect 66378 69606 66430 69658
rect 66442 69606 66494 69658
rect 66506 69606 66558 69658
rect 66570 69606 66622 69658
rect 97034 69606 97086 69658
rect 97098 69606 97150 69658
rect 97162 69606 97214 69658
rect 97226 69606 97278 69658
rect 97290 69606 97342 69658
rect 88984 69164 89036 69216
rect 89168 69164 89220 69216
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 34934 69062 34986 69114
rect 34998 69062 35050 69114
rect 35062 69062 35114 69114
rect 35126 69062 35178 69114
rect 35190 69062 35242 69114
rect 65654 69062 65706 69114
rect 65718 69062 65770 69114
rect 65782 69062 65834 69114
rect 65846 69062 65898 69114
rect 65910 69062 65962 69114
rect 96374 69062 96426 69114
rect 96438 69062 96490 69114
rect 96502 69062 96554 69114
rect 96566 69062 96618 69114
rect 96630 69062 96682 69114
rect 88984 68892 89036 68944
rect 89812 68892 89864 68944
rect 74356 68688 74408 68740
rect 88984 68799 89036 68808
rect 88984 68765 88993 68799
rect 88993 68765 89027 68799
rect 89027 68765 89036 68799
rect 88984 68756 89036 68765
rect 87880 68688 87932 68740
rect 88248 68688 88300 68740
rect 89812 68799 89864 68808
rect 89812 68765 89821 68799
rect 89821 68765 89855 68799
rect 89855 68765 89864 68799
rect 89812 68756 89864 68765
rect 90640 68756 90692 68808
rect 92388 68799 92440 68808
rect 92388 68765 92397 68799
rect 92397 68765 92431 68799
rect 92431 68765 92440 68799
rect 92388 68756 92440 68765
rect 91100 68620 91152 68672
rect 107936 68620 107988 68672
rect 4874 68518 4926 68570
rect 4938 68518 4990 68570
rect 5002 68518 5054 68570
rect 5066 68518 5118 68570
rect 5130 68518 5182 68570
rect 35594 68518 35646 68570
rect 35658 68518 35710 68570
rect 35722 68518 35774 68570
rect 35786 68518 35838 68570
rect 35850 68518 35902 68570
rect 66314 68518 66366 68570
rect 66378 68518 66430 68570
rect 66442 68518 66494 68570
rect 66506 68518 66558 68570
rect 66570 68518 66622 68570
rect 97034 68518 97086 68570
rect 97098 68518 97150 68570
rect 97162 68518 97214 68570
rect 97226 68518 97278 68570
rect 97290 68518 97342 68570
rect 85488 68280 85540 68332
rect 88248 68280 88300 68332
rect 86960 68076 87012 68128
rect 90732 68076 90784 68128
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 34934 67974 34986 68026
rect 34998 67974 35050 68026
rect 35062 67974 35114 68026
rect 35126 67974 35178 68026
rect 35190 67974 35242 68026
rect 65654 67974 65706 68026
rect 65718 67974 65770 68026
rect 65782 67974 65834 68026
rect 65846 67974 65898 68026
rect 65910 67974 65962 68026
rect 96374 67974 96426 68026
rect 96438 67974 96490 68026
rect 96502 67974 96554 68026
rect 96566 67974 96618 68026
rect 96630 67974 96682 68026
rect 90548 67915 90600 67924
rect 90548 67881 90557 67915
rect 90557 67881 90591 67915
rect 90591 67881 90600 67915
rect 90548 67872 90600 67881
rect 107936 67915 107988 67924
rect 107936 67881 107945 67915
rect 107945 67881 107979 67915
rect 107979 67881 107988 67915
rect 107936 67872 107988 67881
rect 101956 67804 102008 67856
rect 84384 67668 84436 67720
rect 85488 67668 85540 67720
rect 88432 67668 88484 67720
rect 87052 67600 87104 67652
rect 89352 67600 89404 67652
rect 89812 67668 89864 67720
rect 90548 67668 90600 67720
rect 91560 67736 91612 67788
rect 92112 67736 92164 67788
rect 91100 67711 91152 67720
rect 91100 67677 91109 67711
rect 91109 67677 91143 67711
rect 91143 67677 91152 67711
rect 91100 67668 91152 67677
rect 92388 67711 92440 67720
rect 92388 67677 92397 67711
rect 92397 67677 92431 67711
rect 92431 67677 92440 67711
rect 92388 67668 92440 67677
rect 108488 67711 108540 67720
rect 108488 67677 108497 67711
rect 108497 67677 108531 67711
rect 108531 67677 108540 67711
rect 108488 67668 108540 67677
rect 102968 67600 103020 67652
rect 89996 67532 90048 67584
rect 91100 67532 91152 67584
rect 4874 67430 4926 67482
rect 4938 67430 4990 67482
rect 5002 67430 5054 67482
rect 5066 67430 5118 67482
rect 5130 67430 5182 67482
rect 35594 67430 35646 67482
rect 35658 67430 35710 67482
rect 35722 67430 35774 67482
rect 35786 67430 35838 67482
rect 35850 67430 35902 67482
rect 66314 67430 66366 67482
rect 66378 67430 66430 67482
rect 66442 67430 66494 67482
rect 66506 67430 66558 67482
rect 66570 67430 66622 67482
rect 97034 67430 97086 67482
rect 97098 67430 97150 67482
rect 97162 67430 97214 67482
rect 97226 67430 97278 67482
rect 97290 67430 97342 67482
rect 88708 67328 88760 67380
rect 89720 67328 89772 67380
rect 90180 67328 90232 67380
rect 84384 67235 84436 67244
rect 84384 67201 84393 67235
rect 84393 67201 84427 67235
rect 84427 67201 84436 67235
rect 84384 67192 84436 67201
rect 87052 67192 87104 67244
rect 89168 67260 89220 67312
rect 91100 67328 91152 67380
rect 92388 67328 92440 67380
rect 88708 67192 88760 67244
rect 89352 67235 89404 67244
rect 89352 67201 89361 67235
rect 89361 67201 89395 67235
rect 89395 67201 89404 67235
rect 89352 67192 89404 67201
rect 89536 67192 89588 67244
rect 90732 67260 90784 67312
rect 89260 67124 89312 67176
rect 89904 67056 89956 67108
rect 84384 66988 84436 67040
rect 85580 66988 85632 67040
rect 88432 66988 88484 67040
rect 88892 66988 88944 67040
rect 89812 67031 89864 67040
rect 89812 66997 89821 67031
rect 89821 66997 89855 67031
rect 89855 66997 89864 67031
rect 89812 66988 89864 66997
rect 90272 67124 90324 67176
rect 91560 67124 91612 67176
rect 95884 66988 95936 67040
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 96374 66886 96426 66938
rect 96438 66886 96490 66938
rect 96502 66886 96554 66938
rect 96566 66886 96618 66938
rect 96630 66886 96682 66938
rect 82084 66784 82136 66836
rect 89260 66784 89312 66836
rect 89352 66716 89404 66768
rect 88156 66648 88208 66700
rect 89168 66691 89220 66700
rect 89168 66657 89177 66691
rect 89177 66657 89211 66691
rect 89211 66657 89220 66691
rect 89168 66648 89220 66657
rect 89260 66580 89312 66632
rect 89904 66648 89956 66700
rect 90640 66716 90692 66768
rect 89996 66580 90048 66632
rect 90272 66623 90324 66632
rect 90272 66589 90281 66623
rect 90281 66589 90315 66623
rect 90315 66589 90324 66623
rect 90272 66580 90324 66589
rect 84292 66555 84344 66564
rect 84292 66521 84301 66555
rect 84301 66521 84335 66555
rect 84335 66521 84344 66555
rect 84292 66512 84344 66521
rect 84384 66512 84436 66564
rect 86960 66512 87012 66564
rect 88892 66555 88944 66564
rect 88892 66521 88901 66555
rect 88901 66521 88935 66555
rect 88935 66521 88944 66555
rect 88892 66512 88944 66521
rect 88984 66512 89036 66564
rect 89352 66555 89404 66564
rect 89352 66521 89361 66555
rect 89361 66521 89395 66555
rect 89395 66521 89404 66555
rect 89352 66512 89404 66521
rect 90640 66580 90692 66632
rect 91284 66580 91336 66632
rect 91376 66580 91428 66632
rect 102324 66580 102376 66632
rect 88708 66444 88760 66496
rect 89720 66444 89772 66496
rect 90548 66555 90600 66564
rect 90548 66521 90557 66555
rect 90557 66521 90591 66555
rect 90591 66521 90600 66555
rect 90548 66512 90600 66521
rect 89996 66444 90048 66496
rect 90456 66444 90508 66496
rect 91928 66487 91980 66496
rect 91928 66453 91937 66487
rect 91937 66453 91971 66487
rect 91971 66453 91980 66487
rect 91928 66444 91980 66453
rect 4874 66342 4926 66394
rect 4938 66342 4990 66394
rect 5002 66342 5054 66394
rect 5066 66342 5118 66394
rect 5130 66342 5182 66394
rect 35594 66342 35646 66394
rect 35658 66342 35710 66394
rect 35722 66342 35774 66394
rect 35786 66342 35838 66394
rect 35850 66342 35902 66394
rect 66314 66342 66366 66394
rect 66378 66342 66430 66394
rect 66442 66342 66494 66394
rect 66506 66342 66558 66394
rect 66570 66342 66622 66394
rect 97034 66342 97086 66394
rect 97098 66342 97150 66394
rect 97162 66342 97214 66394
rect 97226 66342 97278 66394
rect 97290 66342 97342 66394
rect 106658 66342 106710 66394
rect 106722 66342 106774 66394
rect 106786 66342 106838 66394
rect 106850 66342 106902 66394
rect 106914 66342 106966 66394
rect 84292 66240 84344 66292
rect 88432 66283 88484 66292
rect 88432 66249 88441 66283
rect 88441 66249 88475 66283
rect 88475 66249 88484 66283
rect 88432 66240 88484 66249
rect 89444 66240 89496 66292
rect 89720 66240 89772 66292
rect 89904 66240 89956 66292
rect 89996 66240 90048 66292
rect 90732 66240 90784 66292
rect 91008 66283 91060 66292
rect 91008 66249 91017 66283
rect 91017 66249 91051 66283
rect 91051 66249 91060 66283
rect 91008 66240 91060 66249
rect 36084 66215 36136 66224
rect 36084 66181 36093 66215
rect 36093 66181 36127 66215
rect 36127 66181 36136 66215
rect 36084 66172 36136 66181
rect 37924 66172 37976 66224
rect 38476 66172 38528 66224
rect 41144 66215 41196 66224
rect 41144 66181 41153 66215
rect 41153 66181 41187 66215
rect 41187 66181 41196 66215
rect 41144 66172 41196 66181
rect 43628 66215 43680 66224
rect 43628 66181 43637 66215
rect 43637 66181 43671 66215
rect 43671 66181 43680 66215
rect 43628 66172 43680 66181
rect 46112 66215 46164 66224
rect 46112 66181 46121 66215
rect 46121 66181 46155 66215
rect 46155 66181 46164 66215
rect 46112 66172 46164 66181
rect 48596 66215 48648 66224
rect 48596 66181 48605 66215
rect 48605 66181 48639 66215
rect 48639 66181 48648 66215
rect 48596 66172 48648 66181
rect 51080 66215 51132 66224
rect 51080 66181 51089 66215
rect 51089 66181 51123 66215
rect 51123 66181 51132 66215
rect 51080 66172 51132 66181
rect 53564 66215 53616 66224
rect 53564 66181 53573 66215
rect 53573 66181 53607 66215
rect 53607 66181 53616 66215
rect 53564 66172 53616 66181
rect 56140 66215 56192 66224
rect 56140 66181 56149 66215
rect 56149 66181 56183 66215
rect 56183 66181 56192 66215
rect 56140 66172 56192 66181
rect 58624 66215 58676 66224
rect 58624 66181 58633 66215
rect 58633 66181 58667 66215
rect 58667 66181 58676 66215
rect 58624 66172 58676 66181
rect 61108 66215 61160 66224
rect 61108 66181 61117 66215
rect 61117 66181 61151 66215
rect 61151 66181 61160 66215
rect 61108 66172 61160 66181
rect 63592 66215 63644 66224
rect 63592 66181 63601 66215
rect 63601 66181 63635 66215
rect 63635 66181 63644 66215
rect 63592 66172 63644 66181
rect 66076 66215 66128 66224
rect 66076 66181 66085 66215
rect 66085 66181 66119 66215
rect 66119 66181 66128 66215
rect 66076 66172 66128 66181
rect 68560 66215 68612 66224
rect 68560 66181 68569 66215
rect 68569 66181 68603 66215
rect 68603 66181 68612 66215
rect 68560 66172 68612 66181
rect 71044 66215 71096 66224
rect 71044 66181 71053 66215
rect 71053 66181 71087 66215
rect 71087 66181 71096 66215
rect 71044 66172 71096 66181
rect 73528 66215 73580 66224
rect 73528 66181 73537 66215
rect 73537 66181 73571 66215
rect 73571 66181 73580 66215
rect 73528 66172 73580 66181
rect 85580 66172 85632 66224
rect 87604 66172 87656 66224
rect 85672 66147 85724 66156
rect 85672 66113 85681 66147
rect 85681 66113 85715 66147
rect 85715 66113 85724 66147
rect 85672 66104 85724 66113
rect 88156 66104 88208 66156
rect 87604 66036 87656 66088
rect 88064 66036 88116 66088
rect 88984 66079 89036 66088
rect 88984 66045 88993 66079
rect 88993 66045 89027 66079
rect 89027 66045 89036 66079
rect 88984 66036 89036 66045
rect 90456 66172 90508 66224
rect 90916 66172 90968 66224
rect 89444 66079 89496 66088
rect 86224 65943 86276 65952
rect 86224 65909 86233 65943
rect 86233 65909 86267 65943
rect 86267 65909 86276 65943
rect 86224 65900 86276 65909
rect 87880 65900 87932 65952
rect 89444 66045 89453 66079
rect 89453 66045 89487 66079
rect 89487 66045 89496 66079
rect 89444 66036 89496 66045
rect 90364 66147 90416 66156
rect 90364 66113 90373 66147
rect 90373 66113 90407 66147
rect 90407 66113 90416 66147
rect 90364 66104 90416 66113
rect 91376 66240 91428 66292
rect 91928 66240 91980 66292
rect 102140 66240 102192 66292
rect 91560 66215 91612 66224
rect 91560 66181 91587 66215
rect 91587 66181 91612 66215
rect 91560 66172 91612 66181
rect 91192 66147 91244 66156
rect 91192 66113 91201 66147
rect 91201 66113 91235 66147
rect 91235 66113 91244 66147
rect 91192 66104 91244 66113
rect 89260 65968 89312 66020
rect 89352 65968 89404 66020
rect 90640 66036 90692 66088
rect 90732 66036 90784 66088
rect 94320 66215 94372 66224
rect 94320 66181 94329 66215
rect 94329 66181 94363 66215
rect 94363 66181 94372 66215
rect 94320 66172 94372 66181
rect 91928 66147 91980 66156
rect 91928 66113 91937 66147
rect 91937 66113 91971 66147
rect 91971 66113 91980 66147
rect 91928 66104 91980 66113
rect 90640 65900 90692 65952
rect 91284 65900 91336 65952
rect 91560 65943 91612 65952
rect 91560 65909 91569 65943
rect 91569 65909 91603 65943
rect 91603 65909 91612 65943
rect 91560 65900 91612 65909
rect 92296 65943 92348 65952
rect 92296 65909 92305 65943
rect 92305 65909 92339 65943
rect 92339 65909 92348 65943
rect 92296 65900 92348 65909
rect 95884 65943 95936 65952
rect 95884 65909 95893 65943
rect 95893 65909 95927 65943
rect 95927 65909 95936 65943
rect 95884 65900 95936 65909
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 96374 65798 96426 65850
rect 96438 65798 96490 65850
rect 96502 65798 96554 65850
rect 96566 65798 96618 65850
rect 96630 65798 96682 65850
rect 105922 65798 105974 65850
rect 105986 65798 106038 65850
rect 106050 65798 106102 65850
rect 106114 65798 106166 65850
rect 106178 65798 106230 65850
rect 86224 65696 86276 65748
rect 90364 65696 90416 65748
rect 90548 65696 90600 65748
rect 91560 65696 91612 65748
rect 88432 65628 88484 65680
rect 91192 65628 91244 65680
rect 92296 65628 92348 65680
rect 103520 65628 103572 65680
rect 89812 65492 89864 65544
rect 103612 65492 103664 65544
rect 4874 65254 4926 65306
rect 4938 65254 4990 65306
rect 5002 65254 5054 65306
rect 5066 65254 5118 65306
rect 5130 65254 5182 65306
rect 106658 65254 106710 65306
rect 106722 65254 106774 65306
rect 106786 65254 106838 65306
rect 106850 65254 106902 65306
rect 106914 65254 106966 65306
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 105922 64710 105974 64762
rect 105986 64710 106038 64762
rect 106050 64710 106102 64762
rect 106114 64710 106166 64762
rect 106178 64710 106230 64762
rect 4874 64166 4926 64218
rect 4938 64166 4990 64218
rect 5002 64166 5054 64218
rect 5066 64166 5118 64218
rect 5130 64166 5182 64218
rect 106658 64166 106710 64218
rect 106722 64166 106774 64218
rect 106786 64166 106838 64218
rect 106850 64166 106902 64218
rect 106914 64166 106966 64218
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 105922 63622 105974 63674
rect 105986 63622 106038 63674
rect 106050 63622 106102 63674
rect 106114 63622 106166 63674
rect 106178 63622 106230 63674
rect 4874 63078 4926 63130
rect 4938 63078 4990 63130
rect 5002 63078 5054 63130
rect 5066 63078 5118 63130
rect 5130 63078 5182 63130
rect 106658 63078 106710 63130
rect 106722 63078 106774 63130
rect 106786 63078 106838 63130
rect 106850 63078 106902 63130
rect 106914 63078 106966 63130
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 105922 62534 105974 62586
rect 105986 62534 106038 62586
rect 106050 62534 106102 62586
rect 106114 62534 106166 62586
rect 106178 62534 106230 62586
rect 4874 61990 4926 62042
rect 4938 61990 4990 62042
rect 5002 61990 5054 62042
rect 5066 61990 5118 62042
rect 5130 61990 5182 62042
rect 106658 61990 106710 62042
rect 106722 61990 106774 62042
rect 106786 61990 106838 62042
rect 106850 61990 106902 62042
rect 106914 61990 106966 62042
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 105922 61446 105974 61498
rect 105986 61446 106038 61498
rect 106050 61446 106102 61498
rect 106114 61446 106166 61498
rect 106178 61446 106230 61498
rect 4874 60902 4926 60954
rect 4938 60902 4990 60954
rect 5002 60902 5054 60954
rect 5066 60902 5118 60954
rect 5130 60902 5182 60954
rect 106658 60902 106710 60954
rect 106722 60902 106774 60954
rect 106786 60902 106838 60954
rect 106850 60902 106902 60954
rect 106914 60902 106966 60954
rect 7288 60707 7340 60716
rect 7288 60673 7297 60707
rect 7297 60673 7331 60707
rect 7331 60673 7340 60707
rect 7288 60664 7340 60673
rect 6828 60596 6880 60648
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 105922 60358 105974 60410
rect 105986 60358 106038 60410
rect 106050 60358 106102 60410
rect 106114 60358 106166 60410
rect 106178 60358 106230 60410
rect 6828 60256 6880 60308
rect 7288 60052 7340 60104
rect 104348 60095 104400 60104
rect 104348 60061 104357 60095
rect 104357 60061 104391 60095
rect 104391 60061 104400 60095
rect 104348 60052 104400 60061
rect 4874 59814 4926 59866
rect 4938 59814 4990 59866
rect 5002 59814 5054 59866
rect 5066 59814 5118 59866
rect 5130 59814 5182 59866
rect 106658 59814 106710 59866
rect 106722 59814 106774 59866
rect 106786 59814 106838 59866
rect 106850 59814 106902 59866
rect 106914 59814 106966 59866
rect 6828 59712 6880 59764
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 105922 59270 105974 59322
rect 105986 59270 106038 59322
rect 106050 59270 106102 59322
rect 106114 59270 106166 59322
rect 106178 59270 106230 59322
rect 4874 58726 4926 58778
rect 4938 58726 4990 58778
rect 5002 58726 5054 58778
rect 5066 58726 5118 58778
rect 5130 58726 5182 58778
rect 106658 58726 106710 58778
rect 106722 58726 106774 58778
rect 106786 58726 106838 58778
rect 106850 58726 106902 58778
rect 106914 58726 106966 58778
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 105922 58182 105974 58234
rect 105986 58182 106038 58234
rect 106050 58182 106102 58234
rect 106114 58182 106166 58234
rect 106178 58182 106230 58234
rect 4874 57638 4926 57690
rect 4938 57638 4990 57690
rect 5002 57638 5054 57690
rect 5066 57638 5118 57690
rect 5130 57638 5182 57690
rect 106658 57638 106710 57690
rect 106722 57638 106774 57690
rect 106786 57638 106838 57690
rect 106850 57638 106902 57690
rect 106914 57638 106966 57690
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 105922 57094 105974 57146
rect 105986 57094 106038 57146
rect 106050 57094 106102 57146
rect 106114 57094 106166 57146
rect 106178 57094 106230 57146
rect 4874 56550 4926 56602
rect 4938 56550 4990 56602
rect 5002 56550 5054 56602
rect 5066 56550 5118 56602
rect 5130 56550 5182 56602
rect 106658 56550 106710 56602
rect 106722 56550 106774 56602
rect 106786 56550 106838 56602
rect 106850 56550 106902 56602
rect 106914 56550 106966 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 105922 56006 105974 56058
rect 105986 56006 106038 56058
rect 106050 56006 106102 56058
rect 106114 56006 106166 56058
rect 106178 56006 106230 56058
rect 4874 55462 4926 55514
rect 4938 55462 4990 55514
rect 5002 55462 5054 55514
rect 5066 55462 5118 55514
rect 5130 55462 5182 55514
rect 106658 55462 106710 55514
rect 106722 55462 106774 55514
rect 106786 55462 106838 55514
rect 106850 55462 106902 55514
rect 106914 55462 106966 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 105922 54918 105974 54970
rect 105986 54918 106038 54970
rect 106050 54918 106102 54970
rect 106114 54918 106166 54970
rect 106178 54918 106230 54970
rect 4874 54374 4926 54426
rect 4938 54374 4990 54426
rect 5002 54374 5054 54426
rect 5066 54374 5118 54426
rect 5130 54374 5182 54426
rect 106658 54374 106710 54426
rect 106722 54374 106774 54426
rect 106786 54374 106838 54426
rect 106850 54374 106902 54426
rect 106914 54374 106966 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 105922 53830 105974 53882
rect 105986 53830 106038 53882
rect 106050 53830 106102 53882
rect 106114 53830 106166 53882
rect 106178 53830 106230 53882
rect 4874 53286 4926 53338
rect 4938 53286 4990 53338
rect 5002 53286 5054 53338
rect 5066 53286 5118 53338
rect 5130 53286 5182 53338
rect 106658 53286 106710 53338
rect 106722 53286 106774 53338
rect 106786 53286 106838 53338
rect 106850 53286 106902 53338
rect 106914 53286 106966 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 105922 52742 105974 52794
rect 105986 52742 106038 52794
rect 106050 52742 106102 52794
rect 106114 52742 106166 52794
rect 106178 52742 106230 52794
rect 4874 52198 4926 52250
rect 4938 52198 4990 52250
rect 5002 52198 5054 52250
rect 5066 52198 5118 52250
rect 5130 52198 5182 52250
rect 106658 52198 106710 52250
rect 106722 52198 106774 52250
rect 106786 52198 106838 52250
rect 106850 52198 106902 52250
rect 106914 52198 106966 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 105922 51654 105974 51706
rect 105986 51654 106038 51706
rect 106050 51654 106102 51706
rect 106114 51654 106166 51706
rect 106178 51654 106230 51706
rect 4874 51110 4926 51162
rect 4938 51110 4990 51162
rect 5002 51110 5054 51162
rect 5066 51110 5118 51162
rect 5130 51110 5182 51162
rect 106658 51110 106710 51162
rect 106722 51110 106774 51162
rect 106786 51110 106838 51162
rect 106850 51110 106902 51162
rect 106914 51110 106966 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 105922 50566 105974 50618
rect 105986 50566 106038 50618
rect 106050 50566 106102 50618
rect 106114 50566 106166 50618
rect 106178 50566 106230 50618
rect 4874 50022 4926 50074
rect 4938 50022 4990 50074
rect 5002 50022 5054 50074
rect 5066 50022 5118 50074
rect 5130 50022 5182 50074
rect 106658 50022 106710 50074
rect 106722 50022 106774 50074
rect 106786 50022 106838 50074
rect 106850 50022 106902 50074
rect 106914 50022 106966 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 105922 49478 105974 49530
rect 105986 49478 106038 49530
rect 106050 49478 106102 49530
rect 106114 49478 106166 49530
rect 106178 49478 106230 49530
rect 4874 48934 4926 48986
rect 4938 48934 4990 48986
rect 5002 48934 5054 48986
rect 5066 48934 5118 48986
rect 5130 48934 5182 48986
rect 106658 48934 106710 48986
rect 106722 48934 106774 48986
rect 106786 48934 106838 48986
rect 106850 48934 106902 48986
rect 106914 48934 106966 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 105922 48390 105974 48442
rect 105986 48390 106038 48442
rect 106050 48390 106102 48442
rect 106114 48390 106166 48442
rect 106178 48390 106230 48442
rect 4874 47846 4926 47898
rect 4938 47846 4990 47898
rect 5002 47846 5054 47898
rect 5066 47846 5118 47898
rect 5130 47846 5182 47898
rect 106658 47846 106710 47898
rect 106722 47846 106774 47898
rect 106786 47846 106838 47898
rect 106850 47846 106902 47898
rect 106914 47846 106966 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 105922 47302 105974 47354
rect 105986 47302 106038 47354
rect 106050 47302 106102 47354
rect 106114 47302 106166 47354
rect 106178 47302 106230 47354
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 106658 46758 106710 46810
rect 106722 46758 106774 46810
rect 106786 46758 106838 46810
rect 106850 46758 106902 46810
rect 106914 46758 106966 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 105922 46214 105974 46266
rect 105986 46214 106038 46266
rect 106050 46214 106102 46266
rect 106114 46214 106166 46266
rect 106178 46214 106230 46266
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 106658 45670 106710 45722
rect 106722 45670 106774 45722
rect 106786 45670 106838 45722
rect 106850 45670 106902 45722
rect 106914 45670 106966 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 105922 45126 105974 45178
rect 105986 45126 106038 45178
rect 106050 45126 106102 45178
rect 106114 45126 106166 45178
rect 106178 45126 106230 45178
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 106658 44582 106710 44634
rect 106722 44582 106774 44634
rect 106786 44582 106838 44634
rect 106850 44582 106902 44634
rect 106914 44582 106966 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 105922 44038 105974 44090
rect 105986 44038 106038 44090
rect 106050 44038 106102 44090
rect 106114 44038 106166 44090
rect 106178 44038 106230 44090
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 106658 43494 106710 43546
rect 106722 43494 106774 43546
rect 106786 43494 106838 43546
rect 106850 43494 106902 43546
rect 106914 43494 106966 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 105922 42950 105974 43002
rect 105986 42950 106038 43002
rect 106050 42950 106102 43002
rect 106114 42950 106166 43002
rect 106178 42950 106230 43002
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 106658 42406 106710 42458
rect 106722 42406 106774 42458
rect 106786 42406 106838 42458
rect 106850 42406 106902 42458
rect 106914 42406 106966 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 105922 41862 105974 41914
rect 105986 41862 106038 41914
rect 106050 41862 106102 41914
rect 106114 41862 106166 41914
rect 106178 41862 106230 41914
rect 7564 41463 7616 41472
rect 7564 41429 7573 41463
rect 7573 41429 7607 41463
rect 7607 41429 7616 41463
rect 7564 41420 7616 41429
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 106658 41318 106710 41370
rect 106722 41318 106774 41370
rect 106786 41318 106838 41370
rect 106850 41318 106902 41370
rect 106914 41318 106966 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 105922 40774 105974 40826
rect 105986 40774 106038 40826
rect 106050 40774 106102 40826
rect 106114 40774 106166 40826
rect 106178 40774 106230 40826
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 106658 40230 106710 40282
rect 106722 40230 106774 40282
rect 106786 40230 106838 40282
rect 106850 40230 106902 40282
rect 106914 40230 106966 40282
rect 3424 39992 3476 40044
rect 7564 39992 7616 40044
rect 7288 39788 7340 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 105922 39686 105974 39738
rect 105986 39686 106038 39738
rect 106050 39686 106102 39738
rect 106114 39686 106166 39738
rect 106178 39686 106230 39738
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 106658 39142 106710 39194
rect 106722 39142 106774 39194
rect 106786 39142 106838 39194
rect 106850 39142 106902 39194
rect 106914 39142 106966 39194
rect 7564 38743 7616 38752
rect 7564 38709 7573 38743
rect 7573 38709 7607 38743
rect 7607 38709 7616 38743
rect 7564 38700 7616 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 105922 38598 105974 38650
rect 105986 38598 106038 38650
rect 106050 38598 106102 38650
rect 106114 38598 106166 38650
rect 106178 38598 106230 38650
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 106658 38054 106710 38106
rect 106722 38054 106774 38106
rect 106786 38054 106838 38106
rect 106850 38054 106902 38106
rect 106914 38054 106966 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 105922 37510 105974 37562
rect 105986 37510 106038 37562
rect 106050 37510 106102 37562
rect 106114 37510 106166 37562
rect 106178 37510 106230 37562
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 106658 36966 106710 37018
rect 106722 36966 106774 37018
rect 106786 36966 106838 37018
rect 106850 36966 106902 37018
rect 106914 36966 106966 37018
rect 7564 36635 7616 36644
rect 7564 36601 7573 36635
rect 7573 36601 7607 36635
rect 7607 36601 7616 36635
rect 7564 36592 7616 36601
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 105922 36422 105974 36474
rect 105986 36422 106038 36474
rect 106050 36422 106102 36474
rect 106114 36422 106166 36474
rect 106178 36422 106230 36474
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 106658 35878 106710 35930
rect 106722 35878 106774 35930
rect 106786 35878 106838 35930
rect 106850 35878 106902 35930
rect 106914 35878 106966 35930
rect 7472 35479 7524 35488
rect 7472 35445 7481 35479
rect 7481 35445 7515 35479
rect 7515 35445 7524 35479
rect 7472 35436 7524 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 105922 35334 105974 35386
rect 105986 35334 106038 35386
rect 106050 35334 106102 35386
rect 106114 35334 106166 35386
rect 106178 35334 106230 35386
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 106658 34790 106710 34842
rect 106722 34790 106774 34842
rect 106786 34790 106838 34842
rect 106850 34790 106902 34842
rect 106914 34790 106966 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 105922 34246 105974 34298
rect 105986 34246 106038 34298
rect 106050 34246 106102 34298
rect 106114 34246 106166 34298
rect 106178 34246 106230 34298
rect 7564 33915 7616 33924
rect 7564 33881 7573 33915
rect 7573 33881 7607 33915
rect 7607 33881 7616 33915
rect 7564 33872 7616 33881
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 106658 33702 106710 33754
rect 106722 33702 106774 33754
rect 106786 33702 106838 33754
rect 106850 33702 106902 33754
rect 106914 33702 106966 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 105922 33158 105974 33210
rect 105986 33158 106038 33210
rect 106050 33158 106102 33210
rect 106114 33158 106166 33210
rect 106178 33158 106230 33210
rect 1768 33056 1820 33108
rect 7564 33056 7616 33108
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 106658 32614 106710 32666
rect 106722 32614 106774 32666
rect 106786 32614 106838 32666
rect 106850 32614 106902 32666
rect 106914 32614 106966 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 105922 32070 105974 32122
rect 105986 32070 106038 32122
rect 106050 32070 106102 32122
rect 106114 32070 106166 32122
rect 106178 32070 106230 32122
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 106658 31526 106710 31578
rect 106722 31526 106774 31578
rect 106786 31526 106838 31578
rect 106850 31526 106902 31578
rect 106914 31526 106966 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 105922 30982 105974 31034
rect 105986 30982 106038 31034
rect 106050 30982 106102 31034
rect 106114 30982 106166 31034
rect 106178 30982 106230 31034
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 106658 30438 106710 30490
rect 106722 30438 106774 30490
rect 106786 30438 106838 30490
rect 106850 30438 106902 30490
rect 106914 30438 106966 30490
rect 1584 30268 1636 30320
rect 7472 30268 7524 30320
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 105922 29894 105974 29946
rect 105986 29894 106038 29946
rect 106050 29894 106102 29946
rect 106114 29894 106166 29946
rect 106178 29894 106230 29946
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 106658 29350 106710 29402
rect 106722 29350 106774 29402
rect 106786 29350 106838 29402
rect 106850 29350 106902 29402
rect 106914 29350 106966 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 105922 28806 105974 28858
rect 105986 28806 106038 28858
rect 106050 28806 106102 28858
rect 106114 28806 106166 28858
rect 106178 28806 106230 28858
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 106658 28262 106710 28314
rect 106722 28262 106774 28314
rect 106786 28262 106838 28314
rect 106850 28262 106902 28314
rect 106914 28262 106966 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 105922 27718 105974 27770
rect 105986 27718 106038 27770
rect 106050 27718 106102 27770
rect 106114 27718 106166 27770
rect 106178 27718 106230 27770
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 106658 27174 106710 27226
rect 106722 27174 106774 27226
rect 106786 27174 106838 27226
rect 106850 27174 106902 27226
rect 106914 27174 106966 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 105922 26630 105974 26682
rect 105986 26630 106038 26682
rect 106050 26630 106102 26682
rect 106114 26630 106166 26682
rect 106178 26630 106230 26682
rect 1676 26256 1728 26308
rect 7380 26256 7432 26308
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 106658 26086 106710 26138
rect 106722 26086 106774 26138
rect 106786 26086 106838 26138
rect 106850 26086 106902 26138
rect 106914 26086 106966 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 105922 25542 105974 25594
rect 105986 25542 106038 25594
rect 106050 25542 106102 25594
rect 106114 25542 106166 25594
rect 106178 25542 106230 25594
rect 102600 25100 102652 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 106658 24998 106710 25050
rect 106722 24998 106774 25050
rect 106786 24998 106838 25050
rect 106850 24998 106902 25050
rect 106914 24998 106966 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 105922 24454 105974 24506
rect 105986 24454 106038 24506
rect 106050 24454 106102 24506
rect 106114 24454 106166 24506
rect 106178 24454 106230 24506
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 106658 23910 106710 23962
rect 106722 23910 106774 23962
rect 106786 23910 106838 23962
rect 106850 23910 106902 23962
rect 106914 23910 106966 23962
rect 101956 23808 102008 23860
rect 1860 23604 1912 23656
rect 7564 23604 7616 23656
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 105922 23366 105974 23418
rect 105986 23366 106038 23418
rect 106050 23366 106102 23418
rect 106114 23366 106166 23418
rect 106178 23366 106230 23418
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 106658 22822 106710 22874
rect 106722 22822 106774 22874
rect 106786 22822 106838 22874
rect 106850 22822 106902 22874
rect 106914 22822 106966 22874
rect 102324 22720 102376 22772
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 105922 22278 105974 22330
rect 105986 22278 106038 22330
rect 106050 22278 106102 22330
rect 106114 22278 106166 22330
rect 106178 22278 106230 22330
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 106658 21734 106710 21786
rect 106722 21734 106774 21786
rect 106786 21734 106838 21786
rect 106850 21734 106902 21786
rect 106914 21734 106966 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 105922 21190 105974 21242
rect 105986 21190 106038 21242
rect 106050 21190 106102 21242
rect 106114 21190 106166 21242
rect 106178 21190 106230 21242
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 106658 20646 106710 20698
rect 106722 20646 106774 20698
rect 106786 20646 106838 20698
rect 106850 20646 106902 20698
rect 106914 20646 106966 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 105922 20102 105974 20154
rect 105986 20102 106038 20154
rect 106050 20102 106102 20154
rect 106114 20102 106166 20154
rect 106178 20102 106230 20154
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 106658 19558 106710 19610
rect 106722 19558 106774 19610
rect 106786 19558 106838 19610
rect 106850 19558 106902 19610
rect 106914 19558 106966 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 105922 19014 105974 19066
rect 105986 19014 106038 19066
rect 106050 19014 106102 19066
rect 106114 19014 106166 19066
rect 106178 19014 106230 19066
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 106658 18470 106710 18522
rect 106722 18470 106774 18522
rect 106786 18470 106838 18522
rect 106850 18470 106902 18522
rect 106914 18470 106966 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 105922 17926 105974 17978
rect 105986 17926 106038 17978
rect 106050 17926 106102 17978
rect 106114 17926 106166 17978
rect 106178 17926 106230 17978
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 106658 17382 106710 17434
rect 106722 17382 106774 17434
rect 106786 17382 106838 17434
rect 106850 17382 106902 17434
rect 106914 17382 106966 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 105922 16838 105974 16890
rect 105986 16838 106038 16890
rect 106050 16838 106102 16890
rect 106114 16838 106166 16890
rect 106178 16838 106230 16890
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 106658 16294 106710 16346
rect 106722 16294 106774 16346
rect 106786 16294 106838 16346
rect 106850 16294 106902 16346
rect 106914 16294 106966 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 105922 15750 105974 15802
rect 105986 15750 106038 15802
rect 106050 15750 106102 15802
rect 106114 15750 106166 15802
rect 106178 15750 106230 15802
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 106658 15206 106710 15258
rect 106722 15206 106774 15258
rect 106786 15206 106838 15258
rect 106850 15206 106902 15258
rect 106914 15206 106966 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 105922 14662 105974 14714
rect 105986 14662 106038 14714
rect 106050 14662 106102 14714
rect 106114 14662 106166 14714
rect 106178 14662 106230 14714
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 106658 14118 106710 14170
rect 106722 14118 106774 14170
rect 106786 14118 106838 14170
rect 106850 14118 106902 14170
rect 106914 14118 106966 14170
rect 3424 14016 3476 14068
rect 1492 13923 1544 13932
rect 1492 13889 1501 13923
rect 1501 13889 1535 13923
rect 1535 13889 1544 13923
rect 1492 13880 1544 13889
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 105922 13574 105974 13626
rect 105986 13574 106038 13626
rect 106050 13574 106102 13626
rect 106114 13574 106166 13626
rect 106178 13574 106230 13626
rect 1860 13515 1912 13524
rect 1860 13481 1869 13515
rect 1869 13481 1903 13515
rect 1903 13481 1912 13515
rect 1860 13472 1912 13481
rect 1308 13200 1360 13252
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 106658 13030 106710 13082
rect 106722 13030 106774 13082
rect 106786 13030 106838 13082
rect 106850 13030 106902 13082
rect 106914 13030 106966 13082
rect 1676 12903 1728 12912
rect 1676 12869 1685 12903
rect 1685 12869 1719 12903
rect 1719 12869 1728 12903
rect 1676 12860 1728 12869
rect 1492 12835 1544 12844
rect 1492 12801 1501 12835
rect 1501 12801 1535 12835
rect 1535 12801 1544 12835
rect 1492 12792 1544 12801
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 105922 12486 105974 12538
rect 105986 12486 106038 12538
rect 106050 12486 106102 12538
rect 106114 12486 106166 12538
rect 106178 12486 106230 12538
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 106658 11942 106710 11994
rect 106722 11942 106774 11994
rect 106786 11942 106838 11994
rect 106850 11942 106902 11994
rect 106914 11942 106966 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 1216 11704 1268 11756
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 105922 11398 105974 11450
rect 105986 11398 106038 11450
rect 106050 11398 106102 11450
rect 106114 11398 106166 11450
rect 106178 11398 106230 11450
rect 7288 11296 7340 11348
rect 1492 11067 1544 11076
rect 1492 11033 1501 11067
rect 1501 11033 1535 11067
rect 1535 11033 1544 11067
rect 1492 11024 1544 11033
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 106658 10854 106710 10906
rect 106722 10854 106774 10906
rect 106786 10854 106838 10906
rect 106850 10854 106902 10906
rect 106914 10854 106966 10906
rect 1768 10795 1820 10804
rect 1768 10761 1777 10795
rect 1777 10761 1811 10795
rect 1811 10761 1820 10795
rect 1768 10752 1820 10761
rect 1308 10616 1360 10668
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 105922 10310 105974 10362
rect 105986 10310 106038 10362
rect 106050 10310 106102 10362
rect 106114 10310 106166 10362
rect 106178 10310 106230 10362
rect 1492 9979 1544 9988
rect 1492 9945 1501 9979
rect 1501 9945 1535 9979
rect 1535 9945 1544 9979
rect 1492 9936 1544 9945
rect 29552 9868 29604 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 106658 9766 106710 9818
rect 106722 9766 106774 9818
rect 106786 9766 106838 9818
rect 106850 9766 106902 9818
rect 106914 9766 106966 9818
rect 9588 9596 9640 9648
rect 16120 9596 16172 9648
rect 90548 9596 90600 9648
rect 103612 9596 103664 9648
rect 6920 9528 6972 9580
rect 16028 9528 16080 9580
rect 90916 9528 90968 9580
rect 103520 9528 103572 9580
rect 90732 9460 90784 9512
rect 102140 9460 102192 9512
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 105922 9222 105974 9274
rect 105986 9222 106038 9274
rect 106050 9222 106102 9274
rect 106114 9222 106166 9274
rect 106178 9222 106230 9274
rect 1308 8848 1360 8900
rect 26700 8780 26752 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 106658 8678 106710 8730
rect 106722 8678 106774 8730
rect 106786 8678 106838 8730
rect 106850 8678 106902 8730
rect 106914 8678 106966 8730
rect 2044 8372 2096 8424
rect 24676 8304 24728 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 105922 8134 105974 8186
rect 105986 8134 106038 8186
rect 106050 8134 106102 8186
rect 106114 8134 106166 8186
rect 106178 8134 106230 8186
rect 1952 8075 2004 8084
rect 1952 8041 1961 8075
rect 1961 8041 1995 8075
rect 1995 8041 2004 8075
rect 1952 8032 2004 8041
rect 1308 7760 1360 7812
rect 30472 7692 30524 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 66314 7590 66366 7642
rect 66378 7590 66430 7642
rect 66442 7590 66494 7642
rect 66506 7590 66558 7642
rect 66570 7590 66622 7642
rect 97034 7590 97086 7642
rect 97098 7590 97150 7642
rect 97162 7590 97214 7642
rect 97226 7590 97278 7642
rect 97290 7590 97342 7642
rect 106658 7590 106710 7642
rect 106722 7590 106774 7642
rect 106786 7590 106838 7642
rect 106850 7590 106902 7642
rect 106914 7590 106966 7642
rect 16028 7488 16080 7540
rect 23480 7531 23532 7540
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 24676 7531 24728 7540
rect 24676 7497 24685 7531
rect 24685 7497 24719 7531
rect 24719 7497 24728 7531
rect 24676 7488 24728 7497
rect 25780 7488 25832 7540
rect 26700 7488 26752 7540
rect 28172 7531 28224 7540
rect 28172 7497 28181 7531
rect 28181 7497 28215 7531
rect 28215 7497 28224 7531
rect 28172 7488 28224 7497
rect 29552 7531 29604 7540
rect 29552 7497 29561 7531
rect 29561 7497 29595 7531
rect 29595 7497 29604 7531
rect 29552 7488 29604 7497
rect 30472 7531 30524 7540
rect 30472 7497 30481 7531
rect 30481 7497 30515 7531
rect 30515 7497 30524 7531
rect 30472 7488 30524 7497
rect 90548 7531 90600 7540
rect 90548 7497 90557 7531
rect 90557 7497 90591 7531
rect 90591 7497 90600 7531
rect 90548 7488 90600 7497
rect 90732 7531 90784 7540
rect 90732 7497 90741 7531
rect 90741 7497 90775 7531
rect 90775 7497 90784 7531
rect 90732 7488 90784 7497
rect 90916 7531 90968 7540
rect 90916 7497 90925 7531
rect 90925 7497 90959 7531
rect 90959 7497 90968 7531
rect 90916 7488 90968 7497
rect 1308 7352 1360 7404
rect 28172 7216 28224 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 96374 7046 96426 7098
rect 96438 7046 96490 7098
rect 96502 7046 96554 7098
rect 96566 7046 96618 7098
rect 96630 7046 96682 7098
rect 105922 7046 105974 7098
rect 105986 7046 106038 7098
rect 106050 7046 106102 7098
rect 106114 7046 106166 7098
rect 106178 7046 106230 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 66314 6502 66366 6554
rect 66378 6502 66430 6554
rect 66442 6502 66494 6554
rect 66506 6502 66558 6554
rect 66570 6502 66622 6554
rect 97034 6502 97086 6554
rect 97098 6502 97150 6554
rect 97162 6502 97214 6554
rect 97226 6502 97278 6554
rect 97290 6502 97342 6554
rect 1216 6264 1268 6316
rect 25872 6060 25924 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 96374 5958 96426 6010
rect 96438 5958 96490 6010
rect 96502 5958 96554 6010
rect 96566 5958 96618 6010
rect 96630 5958 96682 6010
rect 7472 5856 7524 5908
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 66314 5414 66366 5466
rect 66378 5414 66430 5466
rect 66442 5414 66494 5466
rect 66506 5414 66558 5466
rect 66570 5414 66622 5466
rect 97034 5414 97086 5466
rect 97098 5414 97150 5466
rect 97162 5414 97214 5466
rect 97226 5414 97278 5466
rect 97290 5414 97342 5466
rect 1308 5176 1360 5228
rect 23480 4972 23532 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 96374 4870 96426 4922
rect 96438 4870 96490 4922
rect 96502 4870 96554 4922
rect 96566 4870 96618 4922
rect 96630 4870 96682 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 66314 4326 66366 4378
rect 66378 4326 66430 4378
rect 66442 4326 66494 4378
rect 66506 4326 66558 4378
rect 66570 4326 66622 4378
rect 97034 4326 97086 4378
rect 97098 4326 97150 4378
rect 97162 4326 97214 4378
rect 97226 4326 97278 4378
rect 97290 4326 97342 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 96374 3782 96426 3834
rect 96438 3782 96490 3834
rect 96502 3782 96554 3834
rect 96566 3782 96618 3834
rect 96630 3782 96682 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 66314 3238 66366 3290
rect 66378 3238 66430 3290
rect 66442 3238 66494 3290
rect 66506 3238 66558 3290
rect 66570 3238 66622 3290
rect 97034 3238 97086 3290
rect 97098 3238 97150 3290
rect 97162 3238 97214 3290
rect 97226 3238 97278 3290
rect 97290 3238 97342 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 96374 2694 96426 2746
rect 96438 2694 96490 2746
rect 96502 2694 96554 2746
rect 96566 2694 96618 2746
rect 96630 2694 96682 2746
rect 31668 2635 31720 2644
rect 31668 2601 31677 2635
rect 31677 2601 31711 2635
rect 31711 2601 31720 2635
rect 31668 2592 31720 2601
rect 32956 2635 33008 2644
rect 32956 2601 32965 2635
rect 32965 2601 32999 2635
rect 32999 2601 33008 2635
rect 32956 2592 33008 2601
rect 34244 2635 34296 2644
rect 34244 2601 34253 2635
rect 34253 2601 34287 2635
rect 34287 2601 34296 2635
rect 34244 2592 34296 2601
rect 35440 2592 35492 2644
rect 36360 2635 36412 2644
rect 36360 2601 36369 2635
rect 36369 2601 36403 2635
rect 36403 2601 36412 2635
rect 36360 2592 36412 2601
rect 37464 2635 37516 2644
rect 37464 2601 37473 2635
rect 37473 2601 37507 2635
rect 37507 2601 37516 2635
rect 37464 2592 37516 2601
rect 38752 2635 38804 2644
rect 38752 2601 38761 2635
rect 38761 2601 38795 2635
rect 38795 2601 38804 2635
rect 38752 2592 38804 2601
rect 39948 2592 40000 2644
rect 41328 2635 41380 2644
rect 41328 2601 41337 2635
rect 41337 2601 41371 2635
rect 41371 2601 41380 2635
rect 41328 2592 41380 2601
rect 42156 2635 42208 2644
rect 42156 2601 42165 2635
rect 42165 2601 42199 2635
rect 42199 2601 42208 2635
rect 42156 2592 42208 2601
rect 43444 2635 43496 2644
rect 43444 2601 43453 2635
rect 43453 2601 43487 2635
rect 43487 2601 43496 2635
rect 43444 2592 43496 2601
rect 31576 2295 31628 2304
rect 31576 2261 31585 2295
rect 31585 2261 31619 2295
rect 31619 2261 31628 2295
rect 31576 2252 31628 2261
rect 32864 2295 32916 2304
rect 32864 2261 32873 2295
rect 32873 2261 32907 2295
rect 32907 2261 32916 2295
rect 32864 2252 32916 2261
rect 34152 2295 34204 2304
rect 34152 2261 34161 2295
rect 34161 2261 34195 2295
rect 34195 2261 34204 2295
rect 34152 2252 34204 2261
rect 35440 2295 35492 2304
rect 35440 2261 35449 2295
rect 35449 2261 35483 2295
rect 35483 2261 35492 2295
rect 35440 2252 35492 2261
rect 36084 2295 36136 2304
rect 36084 2261 36093 2295
rect 36093 2261 36127 2295
rect 36127 2261 36136 2295
rect 36084 2252 36136 2261
rect 37372 2295 37424 2304
rect 37372 2261 37381 2295
rect 37381 2261 37415 2295
rect 37415 2261 37424 2295
rect 37372 2252 37424 2261
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 39948 2295 40000 2304
rect 39948 2261 39957 2295
rect 39957 2261 39991 2295
rect 39991 2261 40000 2295
rect 39948 2252 40000 2261
rect 41236 2295 41288 2304
rect 41236 2261 41245 2295
rect 41245 2261 41279 2295
rect 41279 2261 41288 2295
rect 41236 2252 41288 2261
rect 41880 2295 41932 2304
rect 41880 2261 41889 2295
rect 41889 2261 41923 2295
rect 41923 2261 41932 2295
rect 41880 2252 41932 2261
rect 43168 2295 43220 2304
rect 43168 2261 43177 2295
rect 43177 2261 43211 2295
rect 43211 2261 43220 2295
rect 43168 2252 43220 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 66314 2150 66366 2202
rect 66378 2150 66430 2202
rect 66442 2150 66494 2202
rect 66506 2150 66558 2202
rect 66570 2150 66622 2202
rect 97034 2150 97086 2202
rect 97098 2150 97150 2202
rect 97162 2150 97214 2202
rect 97226 2150 97278 2202
rect 97290 2150 97342 2202
<< metal2 >>
rect 4214 147452 4522 147461
rect 4214 147450 4220 147452
rect 4276 147450 4300 147452
rect 4356 147450 4380 147452
rect 4436 147450 4460 147452
rect 4516 147450 4522 147452
rect 4276 147398 4278 147450
rect 4458 147398 4460 147450
rect 4214 147396 4220 147398
rect 4276 147396 4300 147398
rect 4356 147396 4380 147398
rect 4436 147396 4460 147398
rect 4516 147396 4522 147398
rect 4214 147387 4522 147396
rect 34934 147452 35242 147461
rect 34934 147450 34940 147452
rect 34996 147450 35020 147452
rect 35076 147450 35100 147452
rect 35156 147450 35180 147452
rect 35236 147450 35242 147452
rect 34996 147398 34998 147450
rect 35178 147398 35180 147450
rect 34934 147396 34940 147398
rect 34996 147396 35020 147398
rect 35076 147396 35100 147398
rect 35156 147396 35180 147398
rect 35236 147396 35242 147398
rect 34934 147387 35242 147396
rect 65654 147452 65962 147461
rect 65654 147450 65660 147452
rect 65716 147450 65740 147452
rect 65796 147450 65820 147452
rect 65876 147450 65900 147452
rect 65956 147450 65962 147452
rect 65716 147398 65718 147450
rect 65898 147398 65900 147450
rect 65654 147396 65660 147398
rect 65716 147396 65740 147398
rect 65796 147396 65820 147398
rect 65876 147396 65900 147398
rect 65956 147396 65962 147398
rect 65654 147387 65962 147396
rect 96374 147452 96682 147461
rect 96374 147450 96380 147452
rect 96436 147450 96460 147452
rect 96516 147450 96540 147452
rect 96596 147450 96620 147452
rect 96676 147450 96682 147452
rect 96436 147398 96438 147450
rect 96618 147398 96620 147450
rect 96374 147396 96380 147398
rect 96436 147396 96460 147398
rect 96516 147396 96540 147398
rect 96596 147396 96620 147398
rect 96676 147396 96682 147398
rect 96374 147387 96682 147396
rect 4874 146908 5182 146917
rect 4874 146906 4880 146908
rect 4936 146906 4960 146908
rect 5016 146906 5040 146908
rect 5096 146906 5120 146908
rect 5176 146906 5182 146908
rect 4936 146854 4938 146906
rect 5118 146854 5120 146906
rect 4874 146852 4880 146854
rect 4936 146852 4960 146854
rect 5016 146852 5040 146854
rect 5096 146852 5120 146854
rect 5176 146852 5182 146854
rect 4874 146843 5182 146852
rect 35594 146908 35902 146917
rect 35594 146906 35600 146908
rect 35656 146906 35680 146908
rect 35736 146906 35760 146908
rect 35816 146906 35840 146908
rect 35896 146906 35902 146908
rect 35656 146854 35658 146906
rect 35838 146854 35840 146906
rect 35594 146852 35600 146854
rect 35656 146852 35680 146854
rect 35736 146852 35760 146854
rect 35816 146852 35840 146854
rect 35896 146852 35902 146854
rect 35594 146843 35902 146852
rect 66314 146908 66622 146917
rect 66314 146906 66320 146908
rect 66376 146906 66400 146908
rect 66456 146906 66480 146908
rect 66536 146906 66560 146908
rect 66616 146906 66622 146908
rect 66376 146854 66378 146906
rect 66558 146854 66560 146906
rect 66314 146852 66320 146854
rect 66376 146852 66400 146854
rect 66456 146852 66480 146854
rect 66536 146852 66560 146854
rect 66616 146852 66622 146854
rect 66314 146843 66622 146852
rect 97034 146908 97342 146917
rect 97034 146906 97040 146908
rect 97096 146906 97120 146908
rect 97176 146906 97200 146908
rect 97256 146906 97280 146908
rect 97336 146906 97342 146908
rect 97096 146854 97098 146906
rect 97278 146854 97280 146906
rect 97034 146852 97040 146854
rect 97096 146852 97120 146854
rect 97176 146852 97200 146854
rect 97256 146852 97280 146854
rect 97336 146852 97342 146854
rect 97034 146843 97342 146852
rect 4214 146364 4522 146373
rect 4214 146362 4220 146364
rect 4276 146362 4300 146364
rect 4356 146362 4380 146364
rect 4436 146362 4460 146364
rect 4516 146362 4522 146364
rect 4276 146310 4278 146362
rect 4458 146310 4460 146362
rect 4214 146308 4220 146310
rect 4276 146308 4300 146310
rect 4356 146308 4380 146310
rect 4436 146308 4460 146310
rect 4516 146308 4522 146310
rect 4214 146299 4522 146308
rect 34934 146364 35242 146373
rect 34934 146362 34940 146364
rect 34996 146362 35020 146364
rect 35076 146362 35100 146364
rect 35156 146362 35180 146364
rect 35236 146362 35242 146364
rect 34996 146310 34998 146362
rect 35178 146310 35180 146362
rect 34934 146308 34940 146310
rect 34996 146308 35020 146310
rect 35076 146308 35100 146310
rect 35156 146308 35180 146310
rect 35236 146308 35242 146310
rect 34934 146299 35242 146308
rect 65654 146364 65962 146373
rect 65654 146362 65660 146364
rect 65716 146362 65740 146364
rect 65796 146362 65820 146364
rect 65876 146362 65900 146364
rect 65956 146362 65962 146364
rect 65716 146310 65718 146362
rect 65898 146310 65900 146362
rect 65654 146308 65660 146310
rect 65716 146308 65740 146310
rect 65796 146308 65820 146310
rect 65876 146308 65900 146310
rect 65956 146308 65962 146310
rect 65654 146299 65962 146308
rect 96374 146364 96682 146373
rect 96374 146362 96380 146364
rect 96436 146362 96460 146364
rect 96516 146362 96540 146364
rect 96596 146362 96620 146364
rect 96676 146362 96682 146364
rect 96436 146310 96438 146362
rect 96618 146310 96620 146362
rect 96374 146308 96380 146310
rect 96436 146308 96460 146310
rect 96516 146308 96540 146310
rect 96596 146308 96620 146310
rect 96676 146308 96682 146310
rect 96374 146299 96682 146308
rect 4874 145820 5182 145829
rect 4874 145818 4880 145820
rect 4936 145818 4960 145820
rect 5016 145818 5040 145820
rect 5096 145818 5120 145820
rect 5176 145818 5182 145820
rect 4936 145766 4938 145818
rect 5118 145766 5120 145818
rect 4874 145764 4880 145766
rect 4936 145764 4960 145766
rect 5016 145764 5040 145766
rect 5096 145764 5120 145766
rect 5176 145764 5182 145766
rect 4874 145755 5182 145764
rect 35594 145820 35902 145829
rect 35594 145818 35600 145820
rect 35656 145818 35680 145820
rect 35736 145818 35760 145820
rect 35816 145818 35840 145820
rect 35896 145818 35902 145820
rect 35656 145766 35658 145818
rect 35838 145766 35840 145818
rect 35594 145764 35600 145766
rect 35656 145764 35680 145766
rect 35736 145764 35760 145766
rect 35816 145764 35840 145766
rect 35896 145764 35902 145766
rect 35594 145755 35902 145764
rect 66314 145820 66622 145829
rect 66314 145818 66320 145820
rect 66376 145818 66400 145820
rect 66456 145818 66480 145820
rect 66536 145818 66560 145820
rect 66616 145818 66622 145820
rect 66376 145766 66378 145818
rect 66558 145766 66560 145818
rect 66314 145764 66320 145766
rect 66376 145764 66400 145766
rect 66456 145764 66480 145766
rect 66536 145764 66560 145766
rect 66616 145764 66622 145766
rect 66314 145755 66622 145764
rect 97034 145820 97342 145829
rect 97034 145818 97040 145820
rect 97096 145818 97120 145820
rect 97176 145818 97200 145820
rect 97256 145818 97280 145820
rect 97336 145818 97342 145820
rect 97096 145766 97098 145818
rect 97278 145766 97280 145818
rect 97034 145764 97040 145766
rect 97096 145764 97120 145766
rect 97176 145764 97200 145766
rect 97256 145764 97280 145766
rect 97336 145764 97342 145766
rect 97034 145755 97342 145764
rect 4214 145276 4522 145285
rect 4214 145274 4220 145276
rect 4276 145274 4300 145276
rect 4356 145274 4380 145276
rect 4436 145274 4460 145276
rect 4516 145274 4522 145276
rect 4276 145222 4278 145274
rect 4458 145222 4460 145274
rect 4214 145220 4220 145222
rect 4276 145220 4300 145222
rect 4356 145220 4380 145222
rect 4436 145220 4460 145222
rect 4516 145220 4522 145222
rect 4214 145211 4522 145220
rect 34934 145276 35242 145285
rect 34934 145274 34940 145276
rect 34996 145274 35020 145276
rect 35076 145274 35100 145276
rect 35156 145274 35180 145276
rect 35236 145274 35242 145276
rect 34996 145222 34998 145274
rect 35178 145222 35180 145274
rect 34934 145220 34940 145222
rect 34996 145220 35020 145222
rect 35076 145220 35100 145222
rect 35156 145220 35180 145222
rect 35236 145220 35242 145222
rect 34934 145211 35242 145220
rect 65654 145276 65962 145285
rect 65654 145274 65660 145276
rect 65716 145274 65740 145276
rect 65796 145274 65820 145276
rect 65876 145274 65900 145276
rect 65956 145274 65962 145276
rect 65716 145222 65718 145274
rect 65898 145222 65900 145274
rect 65654 145220 65660 145222
rect 65716 145220 65740 145222
rect 65796 145220 65820 145222
rect 65876 145220 65900 145222
rect 65956 145220 65962 145222
rect 65654 145211 65962 145220
rect 96374 145276 96682 145285
rect 96374 145274 96380 145276
rect 96436 145274 96460 145276
rect 96516 145274 96540 145276
rect 96596 145274 96620 145276
rect 96676 145274 96682 145276
rect 96436 145222 96438 145274
rect 96618 145222 96620 145274
rect 96374 145220 96380 145222
rect 96436 145220 96460 145222
rect 96516 145220 96540 145222
rect 96596 145220 96620 145222
rect 96676 145220 96682 145222
rect 96374 145211 96682 145220
rect 4874 144732 5182 144741
rect 4874 144730 4880 144732
rect 4936 144730 4960 144732
rect 5016 144730 5040 144732
rect 5096 144730 5120 144732
rect 5176 144730 5182 144732
rect 4936 144678 4938 144730
rect 5118 144678 5120 144730
rect 4874 144676 4880 144678
rect 4936 144676 4960 144678
rect 5016 144676 5040 144678
rect 5096 144676 5120 144678
rect 5176 144676 5182 144678
rect 4874 144667 5182 144676
rect 35594 144732 35902 144741
rect 35594 144730 35600 144732
rect 35656 144730 35680 144732
rect 35736 144730 35760 144732
rect 35816 144730 35840 144732
rect 35896 144730 35902 144732
rect 35656 144678 35658 144730
rect 35838 144678 35840 144730
rect 35594 144676 35600 144678
rect 35656 144676 35680 144678
rect 35736 144676 35760 144678
rect 35816 144676 35840 144678
rect 35896 144676 35902 144678
rect 35594 144667 35902 144676
rect 66314 144732 66622 144741
rect 66314 144730 66320 144732
rect 66376 144730 66400 144732
rect 66456 144730 66480 144732
rect 66536 144730 66560 144732
rect 66616 144730 66622 144732
rect 66376 144678 66378 144730
rect 66558 144678 66560 144730
rect 66314 144676 66320 144678
rect 66376 144676 66400 144678
rect 66456 144676 66480 144678
rect 66536 144676 66560 144678
rect 66616 144676 66622 144678
rect 66314 144667 66622 144676
rect 97034 144732 97342 144741
rect 97034 144730 97040 144732
rect 97096 144730 97120 144732
rect 97176 144730 97200 144732
rect 97256 144730 97280 144732
rect 97336 144730 97342 144732
rect 97096 144678 97098 144730
rect 97278 144678 97280 144730
rect 97034 144676 97040 144678
rect 97096 144676 97120 144678
rect 97176 144676 97200 144678
rect 97256 144676 97280 144678
rect 97336 144676 97342 144678
rect 97034 144667 97342 144676
rect 4214 144188 4522 144197
rect 4214 144186 4220 144188
rect 4276 144186 4300 144188
rect 4356 144186 4380 144188
rect 4436 144186 4460 144188
rect 4516 144186 4522 144188
rect 4276 144134 4278 144186
rect 4458 144134 4460 144186
rect 4214 144132 4220 144134
rect 4276 144132 4300 144134
rect 4356 144132 4380 144134
rect 4436 144132 4460 144134
rect 4516 144132 4522 144134
rect 4214 144123 4522 144132
rect 34934 144188 35242 144197
rect 34934 144186 34940 144188
rect 34996 144186 35020 144188
rect 35076 144186 35100 144188
rect 35156 144186 35180 144188
rect 35236 144186 35242 144188
rect 34996 144134 34998 144186
rect 35178 144134 35180 144186
rect 34934 144132 34940 144134
rect 34996 144132 35020 144134
rect 35076 144132 35100 144134
rect 35156 144132 35180 144134
rect 35236 144132 35242 144134
rect 34934 144123 35242 144132
rect 65654 144188 65962 144197
rect 65654 144186 65660 144188
rect 65716 144186 65740 144188
rect 65796 144186 65820 144188
rect 65876 144186 65900 144188
rect 65956 144186 65962 144188
rect 65716 144134 65718 144186
rect 65898 144134 65900 144186
rect 65654 144132 65660 144134
rect 65716 144132 65740 144134
rect 65796 144132 65820 144134
rect 65876 144132 65900 144134
rect 65956 144132 65962 144134
rect 65654 144123 65962 144132
rect 96374 144188 96682 144197
rect 96374 144186 96380 144188
rect 96436 144186 96460 144188
rect 96516 144186 96540 144188
rect 96596 144186 96620 144188
rect 96676 144186 96682 144188
rect 96436 144134 96438 144186
rect 96618 144134 96620 144186
rect 96374 144132 96380 144134
rect 96436 144132 96460 144134
rect 96516 144132 96540 144134
rect 96596 144132 96620 144134
rect 96676 144132 96682 144134
rect 96374 144123 96682 144132
rect 4874 143644 5182 143653
rect 4874 143642 4880 143644
rect 4936 143642 4960 143644
rect 5016 143642 5040 143644
rect 5096 143642 5120 143644
rect 5176 143642 5182 143644
rect 4936 143590 4938 143642
rect 5118 143590 5120 143642
rect 4874 143588 4880 143590
rect 4936 143588 4960 143590
rect 5016 143588 5040 143590
rect 5096 143588 5120 143590
rect 5176 143588 5182 143590
rect 4874 143579 5182 143588
rect 35594 143644 35902 143653
rect 35594 143642 35600 143644
rect 35656 143642 35680 143644
rect 35736 143642 35760 143644
rect 35816 143642 35840 143644
rect 35896 143642 35902 143644
rect 35656 143590 35658 143642
rect 35838 143590 35840 143642
rect 35594 143588 35600 143590
rect 35656 143588 35680 143590
rect 35736 143588 35760 143590
rect 35816 143588 35840 143590
rect 35896 143588 35902 143590
rect 35594 143579 35902 143588
rect 66314 143644 66622 143653
rect 66314 143642 66320 143644
rect 66376 143642 66400 143644
rect 66456 143642 66480 143644
rect 66536 143642 66560 143644
rect 66616 143642 66622 143644
rect 66376 143590 66378 143642
rect 66558 143590 66560 143642
rect 66314 143588 66320 143590
rect 66376 143588 66400 143590
rect 66456 143588 66480 143590
rect 66536 143588 66560 143590
rect 66616 143588 66622 143590
rect 66314 143579 66622 143588
rect 97034 143644 97342 143653
rect 97034 143642 97040 143644
rect 97096 143642 97120 143644
rect 97176 143642 97200 143644
rect 97256 143642 97280 143644
rect 97336 143642 97342 143644
rect 97096 143590 97098 143642
rect 97278 143590 97280 143642
rect 97034 143588 97040 143590
rect 97096 143588 97120 143590
rect 97176 143588 97200 143590
rect 97256 143588 97280 143590
rect 97336 143588 97342 143590
rect 97034 143579 97342 143588
rect 4214 143100 4522 143109
rect 4214 143098 4220 143100
rect 4276 143098 4300 143100
rect 4356 143098 4380 143100
rect 4436 143098 4460 143100
rect 4516 143098 4522 143100
rect 4276 143046 4278 143098
rect 4458 143046 4460 143098
rect 4214 143044 4220 143046
rect 4276 143044 4300 143046
rect 4356 143044 4380 143046
rect 4436 143044 4460 143046
rect 4516 143044 4522 143046
rect 4214 143035 4522 143044
rect 34934 143100 35242 143109
rect 34934 143098 34940 143100
rect 34996 143098 35020 143100
rect 35076 143098 35100 143100
rect 35156 143098 35180 143100
rect 35236 143098 35242 143100
rect 34996 143046 34998 143098
rect 35178 143046 35180 143098
rect 34934 143044 34940 143046
rect 34996 143044 35020 143046
rect 35076 143044 35100 143046
rect 35156 143044 35180 143046
rect 35236 143044 35242 143046
rect 34934 143035 35242 143044
rect 65654 143100 65962 143109
rect 65654 143098 65660 143100
rect 65716 143098 65740 143100
rect 65796 143098 65820 143100
rect 65876 143098 65900 143100
rect 65956 143098 65962 143100
rect 65716 143046 65718 143098
rect 65898 143046 65900 143098
rect 65654 143044 65660 143046
rect 65716 143044 65740 143046
rect 65796 143044 65820 143046
rect 65876 143044 65900 143046
rect 65956 143044 65962 143046
rect 65654 143035 65962 143044
rect 96374 143100 96682 143109
rect 96374 143098 96380 143100
rect 96436 143098 96460 143100
rect 96516 143098 96540 143100
rect 96596 143098 96620 143100
rect 96676 143098 96682 143100
rect 96436 143046 96438 143098
rect 96618 143046 96620 143098
rect 96374 143044 96380 143046
rect 96436 143044 96460 143046
rect 96516 143044 96540 143046
rect 96596 143044 96620 143046
rect 96676 143044 96682 143046
rect 96374 143035 96682 143044
rect 4874 142556 5182 142565
rect 4874 142554 4880 142556
rect 4936 142554 4960 142556
rect 5016 142554 5040 142556
rect 5096 142554 5120 142556
rect 5176 142554 5182 142556
rect 4936 142502 4938 142554
rect 5118 142502 5120 142554
rect 4874 142500 4880 142502
rect 4936 142500 4960 142502
rect 5016 142500 5040 142502
rect 5096 142500 5120 142502
rect 5176 142500 5182 142502
rect 4874 142491 5182 142500
rect 35594 142556 35902 142565
rect 35594 142554 35600 142556
rect 35656 142554 35680 142556
rect 35736 142554 35760 142556
rect 35816 142554 35840 142556
rect 35896 142554 35902 142556
rect 35656 142502 35658 142554
rect 35838 142502 35840 142554
rect 35594 142500 35600 142502
rect 35656 142500 35680 142502
rect 35736 142500 35760 142502
rect 35816 142500 35840 142502
rect 35896 142500 35902 142502
rect 35594 142491 35902 142500
rect 66314 142556 66622 142565
rect 66314 142554 66320 142556
rect 66376 142554 66400 142556
rect 66456 142554 66480 142556
rect 66536 142554 66560 142556
rect 66616 142554 66622 142556
rect 66376 142502 66378 142554
rect 66558 142502 66560 142554
rect 66314 142500 66320 142502
rect 66376 142500 66400 142502
rect 66456 142500 66480 142502
rect 66536 142500 66560 142502
rect 66616 142500 66622 142502
rect 66314 142491 66622 142500
rect 97034 142556 97342 142565
rect 97034 142554 97040 142556
rect 97096 142554 97120 142556
rect 97176 142554 97200 142556
rect 97256 142554 97280 142556
rect 97336 142554 97342 142556
rect 97096 142502 97098 142554
rect 97278 142502 97280 142554
rect 97034 142500 97040 142502
rect 97096 142500 97120 142502
rect 97176 142500 97200 142502
rect 97256 142500 97280 142502
rect 97336 142500 97342 142502
rect 97034 142491 97342 142500
rect 4214 142012 4522 142021
rect 4214 142010 4220 142012
rect 4276 142010 4300 142012
rect 4356 142010 4380 142012
rect 4436 142010 4460 142012
rect 4516 142010 4522 142012
rect 4276 141958 4278 142010
rect 4458 141958 4460 142010
rect 4214 141956 4220 141958
rect 4276 141956 4300 141958
rect 4356 141956 4380 141958
rect 4436 141956 4460 141958
rect 4516 141956 4522 141958
rect 4214 141947 4522 141956
rect 34934 142012 35242 142021
rect 34934 142010 34940 142012
rect 34996 142010 35020 142012
rect 35076 142010 35100 142012
rect 35156 142010 35180 142012
rect 35236 142010 35242 142012
rect 34996 141958 34998 142010
rect 35178 141958 35180 142010
rect 34934 141956 34940 141958
rect 34996 141956 35020 141958
rect 35076 141956 35100 141958
rect 35156 141956 35180 141958
rect 35236 141956 35242 141958
rect 34934 141947 35242 141956
rect 65654 142012 65962 142021
rect 65654 142010 65660 142012
rect 65716 142010 65740 142012
rect 65796 142010 65820 142012
rect 65876 142010 65900 142012
rect 65956 142010 65962 142012
rect 65716 141958 65718 142010
rect 65898 141958 65900 142010
rect 65654 141956 65660 141958
rect 65716 141956 65740 141958
rect 65796 141956 65820 141958
rect 65876 141956 65900 141958
rect 65956 141956 65962 141958
rect 65654 141947 65962 141956
rect 96374 142012 96682 142021
rect 96374 142010 96380 142012
rect 96436 142010 96460 142012
rect 96516 142010 96540 142012
rect 96596 142010 96620 142012
rect 96676 142010 96682 142012
rect 96436 141958 96438 142010
rect 96618 141958 96620 142010
rect 96374 141956 96380 141958
rect 96436 141956 96460 141958
rect 96516 141956 96540 141958
rect 96596 141956 96620 141958
rect 96676 141956 96682 141958
rect 96374 141947 96682 141956
rect 4874 141468 5182 141477
rect 4874 141466 4880 141468
rect 4936 141466 4960 141468
rect 5016 141466 5040 141468
rect 5096 141466 5120 141468
rect 5176 141466 5182 141468
rect 4936 141414 4938 141466
rect 5118 141414 5120 141466
rect 4874 141412 4880 141414
rect 4936 141412 4960 141414
rect 5016 141412 5040 141414
rect 5096 141412 5120 141414
rect 5176 141412 5182 141414
rect 4874 141403 5182 141412
rect 35594 141468 35902 141477
rect 35594 141466 35600 141468
rect 35656 141466 35680 141468
rect 35736 141466 35760 141468
rect 35816 141466 35840 141468
rect 35896 141466 35902 141468
rect 35656 141414 35658 141466
rect 35838 141414 35840 141466
rect 35594 141412 35600 141414
rect 35656 141412 35680 141414
rect 35736 141412 35760 141414
rect 35816 141412 35840 141414
rect 35896 141412 35902 141414
rect 35594 141403 35902 141412
rect 66314 141468 66622 141477
rect 66314 141466 66320 141468
rect 66376 141466 66400 141468
rect 66456 141466 66480 141468
rect 66536 141466 66560 141468
rect 66616 141466 66622 141468
rect 66376 141414 66378 141466
rect 66558 141414 66560 141466
rect 66314 141412 66320 141414
rect 66376 141412 66400 141414
rect 66456 141412 66480 141414
rect 66536 141412 66560 141414
rect 66616 141412 66622 141414
rect 66314 141403 66622 141412
rect 97034 141468 97342 141477
rect 97034 141466 97040 141468
rect 97096 141466 97120 141468
rect 97176 141466 97200 141468
rect 97256 141466 97280 141468
rect 97336 141466 97342 141468
rect 97096 141414 97098 141466
rect 97278 141414 97280 141466
rect 97034 141412 97040 141414
rect 97096 141412 97120 141414
rect 97176 141412 97200 141414
rect 97256 141412 97280 141414
rect 97336 141412 97342 141414
rect 97034 141403 97342 141412
rect 4214 140924 4522 140933
rect 4214 140922 4220 140924
rect 4276 140922 4300 140924
rect 4356 140922 4380 140924
rect 4436 140922 4460 140924
rect 4516 140922 4522 140924
rect 4276 140870 4278 140922
rect 4458 140870 4460 140922
rect 4214 140868 4220 140870
rect 4276 140868 4300 140870
rect 4356 140868 4380 140870
rect 4436 140868 4460 140870
rect 4516 140868 4522 140870
rect 4214 140859 4522 140868
rect 34934 140924 35242 140933
rect 34934 140922 34940 140924
rect 34996 140922 35020 140924
rect 35076 140922 35100 140924
rect 35156 140922 35180 140924
rect 35236 140922 35242 140924
rect 34996 140870 34998 140922
rect 35178 140870 35180 140922
rect 34934 140868 34940 140870
rect 34996 140868 35020 140870
rect 35076 140868 35100 140870
rect 35156 140868 35180 140870
rect 35236 140868 35242 140870
rect 34934 140859 35242 140868
rect 65654 140924 65962 140933
rect 65654 140922 65660 140924
rect 65716 140922 65740 140924
rect 65796 140922 65820 140924
rect 65876 140922 65900 140924
rect 65956 140922 65962 140924
rect 65716 140870 65718 140922
rect 65898 140870 65900 140922
rect 65654 140868 65660 140870
rect 65716 140868 65740 140870
rect 65796 140868 65820 140870
rect 65876 140868 65900 140870
rect 65956 140868 65962 140870
rect 65654 140859 65962 140868
rect 96374 140924 96682 140933
rect 96374 140922 96380 140924
rect 96436 140922 96460 140924
rect 96516 140922 96540 140924
rect 96596 140922 96620 140924
rect 96676 140922 96682 140924
rect 96436 140870 96438 140922
rect 96618 140870 96620 140922
rect 96374 140868 96380 140870
rect 96436 140868 96460 140870
rect 96516 140868 96540 140870
rect 96596 140868 96620 140870
rect 96676 140868 96682 140870
rect 96374 140859 96682 140868
rect 4874 140380 5182 140389
rect 4874 140378 4880 140380
rect 4936 140378 4960 140380
rect 5016 140378 5040 140380
rect 5096 140378 5120 140380
rect 5176 140378 5182 140380
rect 4936 140326 4938 140378
rect 5118 140326 5120 140378
rect 4874 140324 4880 140326
rect 4936 140324 4960 140326
rect 5016 140324 5040 140326
rect 5096 140324 5120 140326
rect 5176 140324 5182 140326
rect 4874 140315 5182 140324
rect 35594 140380 35902 140389
rect 35594 140378 35600 140380
rect 35656 140378 35680 140380
rect 35736 140378 35760 140380
rect 35816 140378 35840 140380
rect 35896 140378 35902 140380
rect 35656 140326 35658 140378
rect 35838 140326 35840 140378
rect 35594 140324 35600 140326
rect 35656 140324 35680 140326
rect 35736 140324 35760 140326
rect 35816 140324 35840 140326
rect 35896 140324 35902 140326
rect 35594 140315 35902 140324
rect 66314 140380 66622 140389
rect 66314 140378 66320 140380
rect 66376 140378 66400 140380
rect 66456 140378 66480 140380
rect 66536 140378 66560 140380
rect 66616 140378 66622 140380
rect 66376 140326 66378 140378
rect 66558 140326 66560 140378
rect 66314 140324 66320 140326
rect 66376 140324 66400 140326
rect 66456 140324 66480 140326
rect 66536 140324 66560 140326
rect 66616 140324 66622 140326
rect 66314 140315 66622 140324
rect 97034 140380 97342 140389
rect 97034 140378 97040 140380
rect 97096 140378 97120 140380
rect 97176 140378 97200 140380
rect 97256 140378 97280 140380
rect 97336 140378 97342 140380
rect 97096 140326 97098 140378
rect 97278 140326 97280 140378
rect 97034 140324 97040 140326
rect 97096 140324 97120 140326
rect 97176 140324 97200 140326
rect 97256 140324 97280 140326
rect 97336 140324 97342 140326
rect 97034 140315 97342 140324
rect 4214 139836 4522 139845
rect 4214 139834 4220 139836
rect 4276 139834 4300 139836
rect 4356 139834 4380 139836
rect 4436 139834 4460 139836
rect 4516 139834 4522 139836
rect 4276 139782 4278 139834
rect 4458 139782 4460 139834
rect 4214 139780 4220 139782
rect 4276 139780 4300 139782
rect 4356 139780 4380 139782
rect 4436 139780 4460 139782
rect 4516 139780 4522 139782
rect 4214 139771 4522 139780
rect 34934 139836 35242 139845
rect 34934 139834 34940 139836
rect 34996 139834 35020 139836
rect 35076 139834 35100 139836
rect 35156 139834 35180 139836
rect 35236 139834 35242 139836
rect 34996 139782 34998 139834
rect 35178 139782 35180 139834
rect 34934 139780 34940 139782
rect 34996 139780 35020 139782
rect 35076 139780 35100 139782
rect 35156 139780 35180 139782
rect 35236 139780 35242 139782
rect 34934 139771 35242 139780
rect 65654 139836 65962 139845
rect 65654 139834 65660 139836
rect 65716 139834 65740 139836
rect 65796 139834 65820 139836
rect 65876 139834 65900 139836
rect 65956 139834 65962 139836
rect 65716 139782 65718 139834
rect 65898 139782 65900 139834
rect 65654 139780 65660 139782
rect 65716 139780 65740 139782
rect 65796 139780 65820 139782
rect 65876 139780 65900 139782
rect 65956 139780 65962 139782
rect 65654 139771 65962 139780
rect 96374 139836 96682 139845
rect 96374 139834 96380 139836
rect 96436 139834 96460 139836
rect 96516 139834 96540 139836
rect 96596 139834 96620 139836
rect 96676 139834 96682 139836
rect 96436 139782 96438 139834
rect 96618 139782 96620 139834
rect 96374 139780 96380 139782
rect 96436 139780 96460 139782
rect 96516 139780 96540 139782
rect 96596 139780 96620 139782
rect 96676 139780 96682 139782
rect 96374 139771 96682 139780
rect 4874 139292 5182 139301
rect 4874 139290 4880 139292
rect 4936 139290 4960 139292
rect 5016 139290 5040 139292
rect 5096 139290 5120 139292
rect 5176 139290 5182 139292
rect 4936 139238 4938 139290
rect 5118 139238 5120 139290
rect 4874 139236 4880 139238
rect 4936 139236 4960 139238
rect 5016 139236 5040 139238
rect 5096 139236 5120 139238
rect 5176 139236 5182 139238
rect 4874 139227 5182 139236
rect 35594 139292 35902 139301
rect 35594 139290 35600 139292
rect 35656 139290 35680 139292
rect 35736 139290 35760 139292
rect 35816 139290 35840 139292
rect 35896 139290 35902 139292
rect 35656 139238 35658 139290
rect 35838 139238 35840 139290
rect 35594 139236 35600 139238
rect 35656 139236 35680 139238
rect 35736 139236 35760 139238
rect 35816 139236 35840 139238
rect 35896 139236 35902 139238
rect 35594 139227 35902 139236
rect 66314 139292 66622 139301
rect 66314 139290 66320 139292
rect 66376 139290 66400 139292
rect 66456 139290 66480 139292
rect 66536 139290 66560 139292
rect 66616 139290 66622 139292
rect 66376 139238 66378 139290
rect 66558 139238 66560 139290
rect 66314 139236 66320 139238
rect 66376 139236 66400 139238
rect 66456 139236 66480 139238
rect 66536 139236 66560 139238
rect 66616 139236 66622 139238
rect 66314 139227 66622 139236
rect 97034 139292 97342 139301
rect 97034 139290 97040 139292
rect 97096 139290 97120 139292
rect 97176 139290 97200 139292
rect 97256 139290 97280 139292
rect 97336 139290 97342 139292
rect 97096 139238 97098 139290
rect 97278 139238 97280 139290
rect 97034 139236 97040 139238
rect 97096 139236 97120 139238
rect 97176 139236 97200 139238
rect 97256 139236 97280 139238
rect 97336 139236 97342 139238
rect 97034 139227 97342 139236
rect 4214 138748 4522 138757
rect 4214 138746 4220 138748
rect 4276 138746 4300 138748
rect 4356 138746 4380 138748
rect 4436 138746 4460 138748
rect 4516 138746 4522 138748
rect 4276 138694 4278 138746
rect 4458 138694 4460 138746
rect 4214 138692 4220 138694
rect 4276 138692 4300 138694
rect 4356 138692 4380 138694
rect 4436 138692 4460 138694
rect 4516 138692 4522 138694
rect 4214 138683 4522 138692
rect 34934 138748 35242 138757
rect 34934 138746 34940 138748
rect 34996 138746 35020 138748
rect 35076 138746 35100 138748
rect 35156 138746 35180 138748
rect 35236 138746 35242 138748
rect 34996 138694 34998 138746
rect 35178 138694 35180 138746
rect 34934 138692 34940 138694
rect 34996 138692 35020 138694
rect 35076 138692 35100 138694
rect 35156 138692 35180 138694
rect 35236 138692 35242 138694
rect 34934 138683 35242 138692
rect 65654 138748 65962 138757
rect 65654 138746 65660 138748
rect 65716 138746 65740 138748
rect 65796 138746 65820 138748
rect 65876 138746 65900 138748
rect 65956 138746 65962 138748
rect 65716 138694 65718 138746
rect 65898 138694 65900 138746
rect 65654 138692 65660 138694
rect 65716 138692 65740 138694
rect 65796 138692 65820 138694
rect 65876 138692 65900 138694
rect 65956 138692 65962 138694
rect 65654 138683 65962 138692
rect 96374 138748 96682 138757
rect 96374 138746 96380 138748
rect 96436 138746 96460 138748
rect 96516 138746 96540 138748
rect 96596 138746 96620 138748
rect 96676 138746 96682 138748
rect 96436 138694 96438 138746
rect 96618 138694 96620 138746
rect 96374 138692 96380 138694
rect 96436 138692 96460 138694
rect 96516 138692 96540 138694
rect 96596 138692 96620 138694
rect 96676 138692 96682 138694
rect 96374 138683 96682 138692
rect 4874 138204 5182 138213
rect 4874 138202 4880 138204
rect 4936 138202 4960 138204
rect 5016 138202 5040 138204
rect 5096 138202 5120 138204
rect 5176 138202 5182 138204
rect 4936 138150 4938 138202
rect 5118 138150 5120 138202
rect 4874 138148 4880 138150
rect 4936 138148 4960 138150
rect 5016 138148 5040 138150
rect 5096 138148 5120 138150
rect 5176 138148 5182 138150
rect 4874 138139 5182 138148
rect 35594 138204 35902 138213
rect 35594 138202 35600 138204
rect 35656 138202 35680 138204
rect 35736 138202 35760 138204
rect 35816 138202 35840 138204
rect 35896 138202 35902 138204
rect 35656 138150 35658 138202
rect 35838 138150 35840 138202
rect 35594 138148 35600 138150
rect 35656 138148 35680 138150
rect 35736 138148 35760 138150
rect 35816 138148 35840 138150
rect 35896 138148 35902 138150
rect 35594 138139 35902 138148
rect 66314 138204 66622 138213
rect 66314 138202 66320 138204
rect 66376 138202 66400 138204
rect 66456 138202 66480 138204
rect 66536 138202 66560 138204
rect 66616 138202 66622 138204
rect 66376 138150 66378 138202
rect 66558 138150 66560 138202
rect 66314 138148 66320 138150
rect 66376 138148 66400 138150
rect 66456 138148 66480 138150
rect 66536 138148 66560 138150
rect 66616 138148 66622 138150
rect 66314 138139 66622 138148
rect 97034 138204 97342 138213
rect 97034 138202 97040 138204
rect 97096 138202 97120 138204
rect 97176 138202 97200 138204
rect 97256 138202 97280 138204
rect 97336 138202 97342 138204
rect 97096 138150 97098 138202
rect 97278 138150 97280 138202
rect 97034 138148 97040 138150
rect 97096 138148 97120 138150
rect 97176 138148 97200 138150
rect 97256 138148 97280 138150
rect 97336 138148 97342 138150
rect 97034 138139 97342 138148
rect 4214 137660 4522 137669
rect 4214 137658 4220 137660
rect 4276 137658 4300 137660
rect 4356 137658 4380 137660
rect 4436 137658 4460 137660
rect 4516 137658 4522 137660
rect 4276 137606 4278 137658
rect 4458 137606 4460 137658
rect 4214 137604 4220 137606
rect 4276 137604 4300 137606
rect 4356 137604 4380 137606
rect 4436 137604 4460 137606
rect 4516 137604 4522 137606
rect 4214 137595 4522 137604
rect 34934 137660 35242 137669
rect 34934 137658 34940 137660
rect 34996 137658 35020 137660
rect 35076 137658 35100 137660
rect 35156 137658 35180 137660
rect 35236 137658 35242 137660
rect 34996 137606 34998 137658
rect 35178 137606 35180 137658
rect 34934 137604 34940 137606
rect 34996 137604 35020 137606
rect 35076 137604 35100 137606
rect 35156 137604 35180 137606
rect 35236 137604 35242 137606
rect 34934 137595 35242 137604
rect 65654 137660 65962 137669
rect 65654 137658 65660 137660
rect 65716 137658 65740 137660
rect 65796 137658 65820 137660
rect 65876 137658 65900 137660
rect 65956 137658 65962 137660
rect 65716 137606 65718 137658
rect 65898 137606 65900 137658
rect 65654 137604 65660 137606
rect 65716 137604 65740 137606
rect 65796 137604 65820 137606
rect 65876 137604 65900 137606
rect 65956 137604 65962 137606
rect 65654 137595 65962 137604
rect 96374 137660 96682 137669
rect 96374 137658 96380 137660
rect 96436 137658 96460 137660
rect 96516 137658 96540 137660
rect 96596 137658 96620 137660
rect 96676 137658 96682 137660
rect 96436 137606 96438 137658
rect 96618 137606 96620 137658
rect 96374 137604 96380 137606
rect 96436 137604 96460 137606
rect 96516 137604 96540 137606
rect 96596 137604 96620 137606
rect 96676 137604 96682 137606
rect 96374 137595 96682 137604
rect 4874 137116 5182 137125
rect 4874 137114 4880 137116
rect 4936 137114 4960 137116
rect 5016 137114 5040 137116
rect 5096 137114 5120 137116
rect 5176 137114 5182 137116
rect 4936 137062 4938 137114
rect 5118 137062 5120 137114
rect 4874 137060 4880 137062
rect 4936 137060 4960 137062
rect 5016 137060 5040 137062
rect 5096 137060 5120 137062
rect 5176 137060 5182 137062
rect 4874 137051 5182 137060
rect 35594 137116 35902 137125
rect 35594 137114 35600 137116
rect 35656 137114 35680 137116
rect 35736 137114 35760 137116
rect 35816 137114 35840 137116
rect 35896 137114 35902 137116
rect 35656 137062 35658 137114
rect 35838 137062 35840 137114
rect 35594 137060 35600 137062
rect 35656 137060 35680 137062
rect 35736 137060 35760 137062
rect 35816 137060 35840 137062
rect 35896 137060 35902 137062
rect 35594 137051 35902 137060
rect 66314 137116 66622 137125
rect 66314 137114 66320 137116
rect 66376 137114 66400 137116
rect 66456 137114 66480 137116
rect 66536 137114 66560 137116
rect 66616 137114 66622 137116
rect 66376 137062 66378 137114
rect 66558 137062 66560 137114
rect 66314 137060 66320 137062
rect 66376 137060 66400 137062
rect 66456 137060 66480 137062
rect 66536 137060 66560 137062
rect 66616 137060 66622 137062
rect 66314 137051 66622 137060
rect 97034 137116 97342 137125
rect 97034 137114 97040 137116
rect 97096 137114 97120 137116
rect 97176 137114 97200 137116
rect 97256 137114 97280 137116
rect 97336 137114 97342 137116
rect 97096 137062 97098 137114
rect 97278 137062 97280 137114
rect 97034 137060 97040 137062
rect 97096 137060 97120 137062
rect 97176 137060 97200 137062
rect 97256 137060 97280 137062
rect 97336 137060 97342 137062
rect 97034 137051 97342 137060
rect 4214 136572 4522 136581
rect 4214 136570 4220 136572
rect 4276 136570 4300 136572
rect 4356 136570 4380 136572
rect 4436 136570 4460 136572
rect 4516 136570 4522 136572
rect 4276 136518 4278 136570
rect 4458 136518 4460 136570
rect 4214 136516 4220 136518
rect 4276 136516 4300 136518
rect 4356 136516 4380 136518
rect 4436 136516 4460 136518
rect 4516 136516 4522 136518
rect 4214 136507 4522 136516
rect 34934 136572 35242 136581
rect 34934 136570 34940 136572
rect 34996 136570 35020 136572
rect 35076 136570 35100 136572
rect 35156 136570 35180 136572
rect 35236 136570 35242 136572
rect 34996 136518 34998 136570
rect 35178 136518 35180 136570
rect 34934 136516 34940 136518
rect 34996 136516 35020 136518
rect 35076 136516 35100 136518
rect 35156 136516 35180 136518
rect 35236 136516 35242 136518
rect 34934 136507 35242 136516
rect 65654 136572 65962 136581
rect 65654 136570 65660 136572
rect 65716 136570 65740 136572
rect 65796 136570 65820 136572
rect 65876 136570 65900 136572
rect 65956 136570 65962 136572
rect 65716 136518 65718 136570
rect 65898 136518 65900 136570
rect 65654 136516 65660 136518
rect 65716 136516 65740 136518
rect 65796 136516 65820 136518
rect 65876 136516 65900 136518
rect 65956 136516 65962 136518
rect 65654 136507 65962 136516
rect 96374 136572 96682 136581
rect 96374 136570 96380 136572
rect 96436 136570 96460 136572
rect 96516 136570 96540 136572
rect 96596 136570 96620 136572
rect 96676 136570 96682 136572
rect 96436 136518 96438 136570
rect 96618 136518 96620 136570
rect 96374 136516 96380 136518
rect 96436 136516 96460 136518
rect 96516 136516 96540 136518
rect 96596 136516 96620 136518
rect 96676 136516 96682 136518
rect 96374 136507 96682 136516
rect 105922 136572 106230 136581
rect 105922 136570 105928 136572
rect 105984 136570 106008 136572
rect 106064 136570 106088 136572
rect 106144 136570 106168 136572
rect 106224 136570 106230 136572
rect 105984 136518 105986 136570
rect 106166 136518 106168 136570
rect 105922 136516 105928 136518
rect 105984 136516 106008 136518
rect 106064 136516 106088 136518
rect 106144 136516 106168 136518
rect 106224 136516 106230 136518
rect 105922 136507 106230 136516
rect 101956 136264 102008 136270
rect 101956 136206 102008 136212
rect 38200 136196 38252 136202
rect 38200 136138 38252 136144
rect 40684 136196 40736 136202
rect 40684 136138 40736 136144
rect 42984 136196 43036 136202
rect 42984 136138 43036 136144
rect 46020 136196 46072 136202
rect 46020 136138 46072 136144
rect 48504 136196 48556 136202
rect 48504 136138 48556 136144
rect 52368 136196 52420 136202
rect 52368 136138 52420 136144
rect 55772 136196 55824 136202
rect 55772 136138 55824 136144
rect 58164 136196 58216 136202
rect 58164 136138 58216 136144
rect 60648 136196 60700 136202
rect 60648 136138 60700 136144
rect 63132 136196 63184 136202
rect 63132 136138 63184 136144
rect 64420 136196 64472 136202
rect 64420 136138 64472 136144
rect 67548 136196 67600 136202
rect 67548 136138 67600 136144
rect 69756 136196 69808 136202
rect 69756 136138 69808 136144
rect 72148 136196 72200 136202
rect 72148 136138 72200 136144
rect 74172 136196 74224 136202
rect 74172 136138 74224 136144
rect 9496 136128 9548 136134
rect 9496 136070 9548 136076
rect 36084 136128 36136 136134
rect 36084 136070 36136 136076
rect 38108 136128 38160 136134
rect 38108 136070 38160 136076
rect 4874 136028 5182 136037
rect 4874 136026 4880 136028
rect 4936 136026 4960 136028
rect 5016 136026 5040 136028
rect 5096 136026 5120 136028
rect 5176 136026 5182 136028
rect 4936 135974 4938 136026
rect 5118 135974 5120 136026
rect 4874 135972 4880 135974
rect 4936 135972 4960 135974
rect 5016 135972 5040 135974
rect 5096 135972 5120 135974
rect 5176 135972 5182 135974
rect 4874 135963 5182 135972
rect 8116 135924 8168 135930
rect 8116 135866 8168 135872
rect 8024 135720 8076 135726
rect 8024 135662 8076 135668
rect 4214 135484 4522 135493
rect 4214 135482 4220 135484
rect 4276 135482 4300 135484
rect 4356 135482 4380 135484
rect 4436 135482 4460 135484
rect 4516 135482 4522 135484
rect 4276 135430 4278 135482
rect 4458 135430 4460 135482
rect 4214 135428 4220 135430
rect 4276 135428 4300 135430
rect 4356 135428 4380 135430
rect 4436 135428 4460 135430
rect 4516 135428 4522 135430
rect 4214 135419 4522 135428
rect 4874 134940 5182 134949
rect 4874 134938 4880 134940
rect 4936 134938 4960 134940
rect 5016 134938 5040 134940
rect 5096 134938 5120 134940
rect 5176 134938 5182 134940
rect 4936 134886 4938 134938
rect 5118 134886 5120 134938
rect 4874 134884 4880 134886
rect 4936 134884 4960 134886
rect 5016 134884 5040 134886
rect 5096 134884 5120 134886
rect 5176 134884 5182 134886
rect 4874 134875 5182 134884
rect 4214 134396 4522 134405
rect 4214 134394 4220 134396
rect 4276 134394 4300 134396
rect 4356 134394 4380 134396
rect 4436 134394 4460 134396
rect 4516 134394 4522 134396
rect 4276 134342 4278 134394
rect 4458 134342 4460 134394
rect 4214 134340 4220 134342
rect 4276 134340 4300 134342
rect 4356 134340 4380 134342
rect 4436 134340 4460 134342
rect 4516 134340 4522 134342
rect 4214 134331 4522 134340
rect 7932 133952 7984 133958
rect 7932 133894 7984 133900
rect 4874 133852 5182 133861
rect 4874 133850 4880 133852
rect 4936 133850 4960 133852
rect 5016 133850 5040 133852
rect 5096 133850 5120 133852
rect 5176 133850 5182 133852
rect 4936 133798 4938 133850
rect 5118 133798 5120 133850
rect 4874 133796 4880 133798
rect 4936 133796 4960 133798
rect 5016 133796 5040 133798
rect 5096 133796 5120 133798
rect 5176 133796 5182 133798
rect 4874 133787 5182 133796
rect 4214 133308 4522 133317
rect 4214 133306 4220 133308
rect 4276 133306 4300 133308
rect 4356 133306 4380 133308
rect 4436 133306 4460 133308
rect 4516 133306 4522 133308
rect 4276 133254 4278 133306
rect 4458 133254 4460 133306
rect 4214 133252 4220 133254
rect 4276 133252 4300 133254
rect 4356 133252 4380 133254
rect 4436 133252 4460 133254
rect 4516 133252 4522 133254
rect 4214 133243 4522 133252
rect 4874 132764 5182 132773
rect 4874 132762 4880 132764
rect 4936 132762 4960 132764
rect 5016 132762 5040 132764
rect 5096 132762 5120 132764
rect 5176 132762 5182 132764
rect 4936 132710 4938 132762
rect 5118 132710 5120 132762
rect 4874 132708 4880 132710
rect 4936 132708 4960 132710
rect 5016 132708 5040 132710
rect 5096 132708 5120 132710
rect 5176 132708 5182 132710
rect 4874 132699 5182 132708
rect 4214 132220 4522 132229
rect 4214 132218 4220 132220
rect 4276 132218 4300 132220
rect 4356 132218 4380 132220
rect 4436 132218 4460 132220
rect 4516 132218 4522 132220
rect 4276 132166 4278 132218
rect 4458 132166 4460 132218
rect 4214 132164 4220 132166
rect 4276 132164 4300 132166
rect 4356 132164 4380 132166
rect 4436 132164 4460 132166
rect 4516 132164 4522 132166
rect 4214 132155 4522 132164
rect 4874 131676 5182 131685
rect 4874 131674 4880 131676
rect 4936 131674 4960 131676
rect 5016 131674 5040 131676
rect 5096 131674 5120 131676
rect 5176 131674 5182 131676
rect 4936 131622 4938 131674
rect 5118 131622 5120 131674
rect 4874 131620 4880 131622
rect 4936 131620 4960 131622
rect 5016 131620 5040 131622
rect 5096 131620 5120 131622
rect 5176 131620 5182 131622
rect 4874 131611 5182 131620
rect 4214 131132 4522 131141
rect 4214 131130 4220 131132
rect 4276 131130 4300 131132
rect 4356 131130 4380 131132
rect 4436 131130 4460 131132
rect 4516 131130 4522 131132
rect 4276 131078 4278 131130
rect 4458 131078 4460 131130
rect 4214 131076 4220 131078
rect 4276 131076 4300 131078
rect 4356 131076 4380 131078
rect 4436 131076 4460 131078
rect 4516 131076 4522 131078
rect 4214 131067 4522 131076
rect 4874 130588 5182 130597
rect 4874 130586 4880 130588
rect 4936 130586 4960 130588
rect 5016 130586 5040 130588
rect 5096 130586 5120 130588
rect 5176 130586 5182 130588
rect 4936 130534 4938 130586
rect 5118 130534 5120 130586
rect 4874 130532 4880 130534
rect 4936 130532 4960 130534
rect 5016 130532 5040 130534
rect 5096 130532 5120 130534
rect 5176 130532 5182 130534
rect 4874 130523 5182 130532
rect 4214 130044 4522 130053
rect 4214 130042 4220 130044
rect 4276 130042 4300 130044
rect 4356 130042 4380 130044
rect 4436 130042 4460 130044
rect 4516 130042 4522 130044
rect 4276 129990 4278 130042
rect 4458 129990 4460 130042
rect 4214 129988 4220 129990
rect 4276 129988 4300 129990
rect 4356 129988 4380 129990
rect 4436 129988 4460 129990
rect 4516 129988 4522 129990
rect 4214 129979 4522 129988
rect 4874 129500 5182 129509
rect 4874 129498 4880 129500
rect 4936 129498 4960 129500
rect 5016 129498 5040 129500
rect 5096 129498 5120 129500
rect 5176 129498 5182 129500
rect 4936 129446 4938 129498
rect 5118 129446 5120 129498
rect 4874 129444 4880 129446
rect 4936 129444 4960 129446
rect 5016 129444 5040 129446
rect 5096 129444 5120 129446
rect 5176 129444 5182 129446
rect 4874 129435 5182 129444
rect 4214 128956 4522 128965
rect 4214 128954 4220 128956
rect 4276 128954 4300 128956
rect 4356 128954 4380 128956
rect 4436 128954 4460 128956
rect 4516 128954 4522 128956
rect 4276 128902 4278 128954
rect 4458 128902 4460 128954
rect 4214 128900 4220 128902
rect 4276 128900 4300 128902
rect 4356 128900 4380 128902
rect 4436 128900 4460 128902
rect 4516 128900 4522 128902
rect 4214 128891 4522 128900
rect 4874 128412 5182 128421
rect 4874 128410 4880 128412
rect 4936 128410 4960 128412
rect 5016 128410 5040 128412
rect 5096 128410 5120 128412
rect 5176 128410 5182 128412
rect 4936 128358 4938 128410
rect 5118 128358 5120 128410
rect 4874 128356 4880 128358
rect 4936 128356 4960 128358
rect 5016 128356 5040 128358
rect 5096 128356 5120 128358
rect 5176 128356 5182 128358
rect 4874 128347 5182 128356
rect 4214 127868 4522 127877
rect 4214 127866 4220 127868
rect 4276 127866 4300 127868
rect 4356 127866 4380 127868
rect 4436 127866 4460 127868
rect 4516 127866 4522 127868
rect 4276 127814 4278 127866
rect 4458 127814 4460 127866
rect 4214 127812 4220 127814
rect 4276 127812 4300 127814
rect 4356 127812 4380 127814
rect 4436 127812 4460 127814
rect 4516 127812 4522 127814
rect 4214 127803 4522 127812
rect 4874 127324 5182 127333
rect 4874 127322 4880 127324
rect 4936 127322 4960 127324
rect 5016 127322 5040 127324
rect 5096 127322 5120 127324
rect 5176 127322 5182 127324
rect 4936 127270 4938 127322
rect 5118 127270 5120 127322
rect 4874 127268 4880 127270
rect 4936 127268 4960 127270
rect 5016 127268 5040 127270
rect 5096 127268 5120 127270
rect 5176 127268 5182 127270
rect 4874 127259 5182 127268
rect 4214 126780 4522 126789
rect 4214 126778 4220 126780
rect 4276 126778 4300 126780
rect 4356 126778 4380 126780
rect 4436 126778 4460 126780
rect 4516 126778 4522 126780
rect 4276 126726 4278 126778
rect 4458 126726 4460 126778
rect 4214 126724 4220 126726
rect 4276 126724 4300 126726
rect 4356 126724 4380 126726
rect 4436 126724 4460 126726
rect 4516 126724 4522 126726
rect 4214 126715 4522 126724
rect 4874 126236 5182 126245
rect 4874 126234 4880 126236
rect 4936 126234 4960 126236
rect 5016 126234 5040 126236
rect 5096 126234 5120 126236
rect 5176 126234 5182 126236
rect 4936 126182 4938 126234
rect 5118 126182 5120 126234
rect 4874 126180 4880 126182
rect 4936 126180 4960 126182
rect 5016 126180 5040 126182
rect 5096 126180 5120 126182
rect 5176 126180 5182 126182
rect 4874 126171 5182 126180
rect 4214 125692 4522 125701
rect 4214 125690 4220 125692
rect 4276 125690 4300 125692
rect 4356 125690 4380 125692
rect 4436 125690 4460 125692
rect 4516 125690 4522 125692
rect 4276 125638 4278 125690
rect 4458 125638 4460 125690
rect 4214 125636 4220 125638
rect 4276 125636 4300 125638
rect 4356 125636 4380 125638
rect 4436 125636 4460 125638
rect 4516 125636 4522 125638
rect 4214 125627 4522 125636
rect 4874 125148 5182 125157
rect 4874 125146 4880 125148
rect 4936 125146 4960 125148
rect 5016 125146 5040 125148
rect 5096 125146 5120 125148
rect 5176 125146 5182 125148
rect 4936 125094 4938 125146
rect 5118 125094 5120 125146
rect 4874 125092 4880 125094
rect 4936 125092 4960 125094
rect 5016 125092 5040 125094
rect 5096 125092 5120 125094
rect 5176 125092 5182 125094
rect 4874 125083 5182 125092
rect 4214 124604 4522 124613
rect 4214 124602 4220 124604
rect 4276 124602 4300 124604
rect 4356 124602 4380 124604
rect 4436 124602 4460 124604
rect 4516 124602 4522 124604
rect 4276 124550 4278 124602
rect 4458 124550 4460 124602
rect 4214 124548 4220 124550
rect 4276 124548 4300 124550
rect 4356 124548 4380 124550
rect 4436 124548 4460 124550
rect 4516 124548 4522 124550
rect 4214 124539 4522 124548
rect 4874 124060 5182 124069
rect 4874 124058 4880 124060
rect 4936 124058 4960 124060
rect 5016 124058 5040 124060
rect 5096 124058 5120 124060
rect 5176 124058 5182 124060
rect 4936 124006 4938 124058
rect 5118 124006 5120 124058
rect 4874 124004 4880 124006
rect 4936 124004 4960 124006
rect 5016 124004 5040 124006
rect 5096 124004 5120 124006
rect 5176 124004 5182 124006
rect 4874 123995 5182 124004
rect 4214 123516 4522 123525
rect 4214 123514 4220 123516
rect 4276 123514 4300 123516
rect 4356 123514 4380 123516
rect 4436 123514 4460 123516
rect 4516 123514 4522 123516
rect 4276 123462 4278 123514
rect 4458 123462 4460 123514
rect 4214 123460 4220 123462
rect 4276 123460 4300 123462
rect 4356 123460 4380 123462
rect 4436 123460 4460 123462
rect 4516 123460 4522 123462
rect 4214 123451 4522 123460
rect 4874 122972 5182 122981
rect 4874 122970 4880 122972
rect 4936 122970 4960 122972
rect 5016 122970 5040 122972
rect 5096 122970 5120 122972
rect 5176 122970 5182 122972
rect 4936 122918 4938 122970
rect 5118 122918 5120 122970
rect 4874 122916 4880 122918
rect 4936 122916 4960 122918
rect 5016 122916 5040 122918
rect 5096 122916 5120 122918
rect 5176 122916 5182 122918
rect 4874 122907 5182 122916
rect 4214 122428 4522 122437
rect 4214 122426 4220 122428
rect 4276 122426 4300 122428
rect 4356 122426 4380 122428
rect 4436 122426 4460 122428
rect 4516 122426 4522 122428
rect 4276 122374 4278 122426
rect 4458 122374 4460 122426
rect 4214 122372 4220 122374
rect 4276 122372 4300 122374
rect 4356 122372 4380 122374
rect 4436 122372 4460 122374
rect 4516 122372 4522 122374
rect 4214 122363 4522 122372
rect 4874 121884 5182 121893
rect 4874 121882 4880 121884
rect 4936 121882 4960 121884
rect 5016 121882 5040 121884
rect 5096 121882 5120 121884
rect 5176 121882 5182 121884
rect 4936 121830 4938 121882
rect 5118 121830 5120 121882
rect 4874 121828 4880 121830
rect 4936 121828 4960 121830
rect 5016 121828 5040 121830
rect 5096 121828 5120 121830
rect 5176 121828 5182 121830
rect 4874 121819 5182 121828
rect 4214 121340 4522 121349
rect 4214 121338 4220 121340
rect 4276 121338 4300 121340
rect 4356 121338 4380 121340
rect 4436 121338 4460 121340
rect 4516 121338 4522 121340
rect 4276 121286 4278 121338
rect 4458 121286 4460 121338
rect 4214 121284 4220 121286
rect 4276 121284 4300 121286
rect 4356 121284 4380 121286
rect 4436 121284 4460 121286
rect 4516 121284 4522 121286
rect 4214 121275 4522 121284
rect 4874 120796 5182 120805
rect 4874 120794 4880 120796
rect 4936 120794 4960 120796
rect 5016 120794 5040 120796
rect 5096 120794 5120 120796
rect 5176 120794 5182 120796
rect 4936 120742 4938 120794
rect 5118 120742 5120 120794
rect 4874 120740 4880 120742
rect 4936 120740 4960 120742
rect 5016 120740 5040 120742
rect 5096 120740 5120 120742
rect 5176 120740 5182 120742
rect 4874 120731 5182 120740
rect 4214 120252 4522 120261
rect 4214 120250 4220 120252
rect 4276 120250 4300 120252
rect 4356 120250 4380 120252
rect 4436 120250 4460 120252
rect 4516 120250 4522 120252
rect 4276 120198 4278 120250
rect 4458 120198 4460 120250
rect 4214 120196 4220 120198
rect 4276 120196 4300 120198
rect 4356 120196 4380 120198
rect 4436 120196 4460 120198
rect 4516 120196 4522 120198
rect 4214 120187 4522 120196
rect 4874 119708 5182 119717
rect 4874 119706 4880 119708
rect 4936 119706 4960 119708
rect 5016 119706 5040 119708
rect 5096 119706 5120 119708
rect 5176 119706 5182 119708
rect 4936 119654 4938 119706
rect 5118 119654 5120 119706
rect 4874 119652 4880 119654
rect 4936 119652 4960 119654
rect 5016 119652 5040 119654
rect 5096 119652 5120 119654
rect 5176 119652 5182 119654
rect 4874 119643 5182 119652
rect 4214 119164 4522 119173
rect 4214 119162 4220 119164
rect 4276 119162 4300 119164
rect 4356 119162 4380 119164
rect 4436 119162 4460 119164
rect 4516 119162 4522 119164
rect 4276 119110 4278 119162
rect 4458 119110 4460 119162
rect 4214 119108 4220 119110
rect 4276 119108 4300 119110
rect 4356 119108 4380 119110
rect 4436 119108 4460 119110
rect 4516 119108 4522 119110
rect 4214 119099 4522 119108
rect 4874 118620 5182 118629
rect 4874 118618 4880 118620
rect 4936 118618 4960 118620
rect 5016 118618 5040 118620
rect 5096 118618 5120 118620
rect 5176 118618 5182 118620
rect 4936 118566 4938 118618
rect 5118 118566 5120 118618
rect 4874 118564 4880 118566
rect 4936 118564 4960 118566
rect 5016 118564 5040 118566
rect 5096 118564 5120 118566
rect 5176 118564 5182 118566
rect 4874 118555 5182 118564
rect 4214 118076 4522 118085
rect 4214 118074 4220 118076
rect 4276 118074 4300 118076
rect 4356 118074 4380 118076
rect 4436 118074 4460 118076
rect 4516 118074 4522 118076
rect 4276 118022 4278 118074
rect 4458 118022 4460 118074
rect 4214 118020 4220 118022
rect 4276 118020 4300 118022
rect 4356 118020 4380 118022
rect 4436 118020 4460 118022
rect 4516 118020 4522 118022
rect 4214 118011 4522 118020
rect 4874 117532 5182 117541
rect 4874 117530 4880 117532
rect 4936 117530 4960 117532
rect 5016 117530 5040 117532
rect 5096 117530 5120 117532
rect 5176 117530 5182 117532
rect 4936 117478 4938 117530
rect 5118 117478 5120 117530
rect 4874 117476 4880 117478
rect 4936 117476 4960 117478
rect 5016 117476 5040 117478
rect 5096 117476 5120 117478
rect 5176 117476 5182 117478
rect 4874 117467 5182 117476
rect 4214 116988 4522 116997
rect 4214 116986 4220 116988
rect 4276 116986 4300 116988
rect 4356 116986 4380 116988
rect 4436 116986 4460 116988
rect 4516 116986 4522 116988
rect 4276 116934 4278 116986
rect 4458 116934 4460 116986
rect 4214 116932 4220 116934
rect 4276 116932 4300 116934
rect 4356 116932 4380 116934
rect 4436 116932 4460 116934
rect 4516 116932 4522 116934
rect 4214 116923 4522 116932
rect 4874 116444 5182 116453
rect 4874 116442 4880 116444
rect 4936 116442 4960 116444
rect 5016 116442 5040 116444
rect 5096 116442 5120 116444
rect 5176 116442 5182 116444
rect 4936 116390 4938 116442
rect 5118 116390 5120 116442
rect 4874 116388 4880 116390
rect 4936 116388 4960 116390
rect 5016 116388 5040 116390
rect 5096 116388 5120 116390
rect 5176 116388 5182 116390
rect 4874 116379 5182 116388
rect 4214 115900 4522 115909
rect 4214 115898 4220 115900
rect 4276 115898 4300 115900
rect 4356 115898 4380 115900
rect 4436 115898 4460 115900
rect 4516 115898 4522 115900
rect 4276 115846 4278 115898
rect 4458 115846 4460 115898
rect 4214 115844 4220 115846
rect 4276 115844 4300 115846
rect 4356 115844 4380 115846
rect 4436 115844 4460 115846
rect 4516 115844 4522 115846
rect 4214 115835 4522 115844
rect 4874 115356 5182 115365
rect 4874 115354 4880 115356
rect 4936 115354 4960 115356
rect 5016 115354 5040 115356
rect 5096 115354 5120 115356
rect 5176 115354 5182 115356
rect 4936 115302 4938 115354
rect 5118 115302 5120 115354
rect 4874 115300 4880 115302
rect 4936 115300 4960 115302
rect 5016 115300 5040 115302
rect 5096 115300 5120 115302
rect 5176 115300 5182 115302
rect 4874 115291 5182 115300
rect 4214 114812 4522 114821
rect 4214 114810 4220 114812
rect 4276 114810 4300 114812
rect 4356 114810 4380 114812
rect 4436 114810 4460 114812
rect 4516 114810 4522 114812
rect 4276 114758 4278 114810
rect 4458 114758 4460 114810
rect 4214 114756 4220 114758
rect 4276 114756 4300 114758
rect 4356 114756 4380 114758
rect 4436 114756 4460 114758
rect 4516 114756 4522 114758
rect 4214 114747 4522 114756
rect 4874 114268 5182 114277
rect 4874 114266 4880 114268
rect 4936 114266 4960 114268
rect 5016 114266 5040 114268
rect 5096 114266 5120 114268
rect 5176 114266 5182 114268
rect 4936 114214 4938 114266
rect 5118 114214 5120 114266
rect 4874 114212 4880 114214
rect 4936 114212 4960 114214
rect 5016 114212 5040 114214
rect 5096 114212 5120 114214
rect 5176 114212 5182 114214
rect 4874 114203 5182 114212
rect 4214 113724 4522 113733
rect 4214 113722 4220 113724
rect 4276 113722 4300 113724
rect 4356 113722 4380 113724
rect 4436 113722 4460 113724
rect 4516 113722 4522 113724
rect 4276 113670 4278 113722
rect 4458 113670 4460 113722
rect 4214 113668 4220 113670
rect 4276 113668 4300 113670
rect 4356 113668 4380 113670
rect 4436 113668 4460 113670
rect 4516 113668 4522 113670
rect 4214 113659 4522 113668
rect 4874 113180 5182 113189
rect 4874 113178 4880 113180
rect 4936 113178 4960 113180
rect 5016 113178 5040 113180
rect 5096 113178 5120 113180
rect 5176 113178 5182 113180
rect 4936 113126 4938 113178
rect 5118 113126 5120 113178
rect 4874 113124 4880 113126
rect 4936 113124 4960 113126
rect 5016 113124 5040 113126
rect 5096 113124 5120 113126
rect 5176 113124 5182 113126
rect 4874 113115 5182 113124
rect 4214 112636 4522 112645
rect 4214 112634 4220 112636
rect 4276 112634 4300 112636
rect 4356 112634 4380 112636
rect 4436 112634 4460 112636
rect 4516 112634 4522 112636
rect 4276 112582 4278 112634
rect 4458 112582 4460 112634
rect 4214 112580 4220 112582
rect 4276 112580 4300 112582
rect 4356 112580 4380 112582
rect 4436 112580 4460 112582
rect 4516 112580 4522 112582
rect 4214 112571 4522 112580
rect 4874 112092 5182 112101
rect 4874 112090 4880 112092
rect 4936 112090 4960 112092
rect 5016 112090 5040 112092
rect 5096 112090 5120 112092
rect 5176 112090 5182 112092
rect 4936 112038 4938 112090
rect 5118 112038 5120 112090
rect 4874 112036 4880 112038
rect 4936 112036 4960 112038
rect 5016 112036 5040 112038
rect 5096 112036 5120 112038
rect 5176 112036 5182 112038
rect 4874 112027 5182 112036
rect 4214 111548 4522 111557
rect 4214 111546 4220 111548
rect 4276 111546 4300 111548
rect 4356 111546 4380 111548
rect 4436 111546 4460 111548
rect 4516 111546 4522 111548
rect 4276 111494 4278 111546
rect 4458 111494 4460 111546
rect 4214 111492 4220 111494
rect 4276 111492 4300 111494
rect 4356 111492 4380 111494
rect 4436 111492 4460 111494
rect 4516 111492 4522 111494
rect 4214 111483 4522 111492
rect 1308 111240 1360 111246
rect 1308 111182 1360 111188
rect 1320 110945 1348 111182
rect 4874 111004 5182 111013
rect 4874 111002 4880 111004
rect 4936 111002 4960 111004
rect 5016 111002 5040 111004
rect 5096 111002 5120 111004
rect 5176 111002 5182 111004
rect 4936 110950 4938 111002
rect 5118 110950 5120 111002
rect 4874 110948 4880 110950
rect 4936 110948 4960 110950
rect 5016 110948 5040 110950
rect 5096 110948 5120 110950
rect 5176 110948 5182 110950
rect 1306 110936 1362 110945
rect 4874 110939 5182 110948
rect 1306 110871 1362 110880
rect 4214 110460 4522 110469
rect 4214 110458 4220 110460
rect 4276 110458 4300 110460
rect 4356 110458 4380 110460
rect 4436 110458 4460 110460
rect 4516 110458 4522 110460
rect 4276 110406 4278 110458
rect 4458 110406 4460 110458
rect 4214 110404 4220 110406
rect 4276 110404 4300 110406
rect 4356 110404 4380 110406
rect 4436 110404 4460 110406
rect 4516 110404 4522 110406
rect 4214 110395 4522 110404
rect 4874 109916 5182 109925
rect 4874 109914 4880 109916
rect 4936 109914 4960 109916
rect 5016 109914 5040 109916
rect 5096 109914 5120 109916
rect 5176 109914 5182 109916
rect 4936 109862 4938 109914
rect 5118 109862 5120 109914
rect 4874 109860 4880 109862
rect 4936 109860 4960 109862
rect 5016 109860 5040 109862
rect 5096 109860 5120 109862
rect 5176 109860 5182 109862
rect 4874 109851 5182 109860
rect 1308 109676 1360 109682
rect 1308 109618 1360 109624
rect 1320 109585 1348 109618
rect 1306 109576 1362 109585
rect 1306 109511 1362 109520
rect 4214 109372 4522 109381
rect 4214 109370 4220 109372
rect 4276 109370 4300 109372
rect 4356 109370 4380 109372
rect 4436 109370 4460 109372
rect 4516 109370 4522 109372
rect 4276 109318 4278 109370
rect 4458 109318 4460 109370
rect 4214 109316 4220 109318
rect 4276 109316 4300 109318
rect 4356 109316 4380 109318
rect 4436 109316 4460 109318
rect 4516 109316 4522 109318
rect 4214 109307 4522 109316
rect 4874 108828 5182 108837
rect 4874 108826 4880 108828
rect 4936 108826 4960 108828
rect 5016 108826 5040 108828
rect 5096 108826 5120 108828
rect 5176 108826 5182 108828
rect 4936 108774 4938 108826
rect 5118 108774 5120 108826
rect 4874 108772 4880 108774
rect 4936 108772 4960 108774
rect 5016 108772 5040 108774
rect 5096 108772 5120 108774
rect 5176 108772 5182 108774
rect 4874 108763 5182 108772
rect 1308 108588 1360 108594
rect 1308 108530 1360 108536
rect 1320 108225 1348 108530
rect 4214 108284 4522 108293
rect 4214 108282 4220 108284
rect 4276 108282 4300 108284
rect 4356 108282 4380 108284
rect 4436 108282 4460 108284
rect 4516 108282 4522 108284
rect 4276 108230 4278 108282
rect 4458 108230 4460 108282
rect 4214 108228 4220 108230
rect 4276 108228 4300 108230
rect 4356 108228 4380 108230
rect 4436 108228 4460 108230
rect 4516 108228 4522 108230
rect 1306 108216 1362 108225
rect 4214 108219 4522 108228
rect 1306 108151 1362 108160
rect 4874 107740 5182 107749
rect 4874 107738 4880 107740
rect 4936 107738 4960 107740
rect 5016 107738 5040 107740
rect 5096 107738 5120 107740
rect 5176 107738 5182 107740
rect 4936 107686 4938 107738
rect 5118 107686 5120 107738
rect 4874 107684 4880 107686
rect 4936 107684 4960 107686
rect 5016 107684 5040 107686
rect 5096 107684 5120 107686
rect 5176 107684 5182 107686
rect 4874 107675 5182 107684
rect 4214 107196 4522 107205
rect 4214 107194 4220 107196
rect 4276 107194 4300 107196
rect 4356 107194 4380 107196
rect 4436 107194 4460 107196
rect 4516 107194 4522 107196
rect 4276 107142 4278 107194
rect 4458 107142 4460 107194
rect 4214 107140 4220 107142
rect 4276 107140 4300 107142
rect 4356 107140 4380 107142
rect 4436 107140 4460 107142
rect 4516 107140 4522 107142
rect 4214 107131 4522 107140
rect 1216 106888 1268 106894
rect 1214 106856 1216 106865
rect 1268 106856 1270 106865
rect 1214 106791 1270 106800
rect 4874 106652 5182 106661
rect 4874 106650 4880 106652
rect 4936 106650 4960 106652
rect 5016 106650 5040 106652
rect 5096 106650 5120 106652
rect 5176 106650 5182 106652
rect 4936 106598 4938 106650
rect 5118 106598 5120 106650
rect 4874 106596 4880 106598
rect 4936 106596 4960 106598
rect 5016 106596 5040 106598
rect 5096 106596 5120 106598
rect 5176 106596 5182 106598
rect 4874 106587 5182 106596
rect 4214 106108 4522 106117
rect 4214 106106 4220 106108
rect 4276 106106 4300 106108
rect 4356 106106 4380 106108
rect 4436 106106 4460 106108
rect 4516 106106 4522 106108
rect 4276 106054 4278 106106
rect 4458 106054 4460 106106
rect 4214 106052 4220 106054
rect 4276 106052 4300 106054
rect 4356 106052 4380 106054
rect 4436 106052 4460 106054
rect 4516 106052 4522 106054
rect 4214 106043 4522 106052
rect 1308 105800 1360 105806
rect 1308 105742 1360 105748
rect 1320 105505 1348 105742
rect 4874 105564 5182 105573
rect 4874 105562 4880 105564
rect 4936 105562 4960 105564
rect 5016 105562 5040 105564
rect 5096 105562 5120 105564
rect 5176 105562 5182 105564
rect 4936 105510 4938 105562
rect 5118 105510 5120 105562
rect 4874 105508 4880 105510
rect 4936 105508 4960 105510
rect 5016 105508 5040 105510
rect 5096 105508 5120 105510
rect 5176 105508 5182 105510
rect 1306 105496 1362 105505
rect 4874 105499 5182 105508
rect 1306 105431 1362 105440
rect 4214 105020 4522 105029
rect 4214 105018 4220 105020
rect 4276 105018 4300 105020
rect 4356 105018 4380 105020
rect 4436 105018 4460 105020
rect 4516 105018 4522 105020
rect 4276 104966 4278 105018
rect 4458 104966 4460 105018
rect 4214 104964 4220 104966
rect 4276 104964 4300 104966
rect 4356 104964 4380 104966
rect 4436 104964 4460 104966
rect 4516 104964 4522 104966
rect 4214 104955 4522 104964
rect 4874 104476 5182 104485
rect 4874 104474 4880 104476
rect 4936 104474 4960 104476
rect 5016 104474 5040 104476
rect 5096 104474 5120 104476
rect 5176 104474 5182 104476
rect 4936 104422 4938 104474
rect 5118 104422 5120 104474
rect 4874 104420 4880 104422
rect 4936 104420 4960 104422
rect 5016 104420 5040 104422
rect 5096 104420 5120 104422
rect 5176 104420 5182 104422
rect 4874 104411 5182 104420
rect 1308 104236 1360 104242
rect 1308 104178 1360 104184
rect 1320 104145 1348 104178
rect 1306 104136 1362 104145
rect 1306 104071 1362 104080
rect 4214 103932 4522 103941
rect 4214 103930 4220 103932
rect 4276 103930 4300 103932
rect 4356 103930 4380 103932
rect 4436 103930 4460 103932
rect 4516 103930 4522 103932
rect 4276 103878 4278 103930
rect 4458 103878 4460 103930
rect 4214 103876 4220 103878
rect 4276 103876 4300 103878
rect 4356 103876 4380 103878
rect 4436 103876 4460 103878
rect 4516 103876 4522 103878
rect 4214 103867 4522 103876
rect 4874 103388 5182 103397
rect 4874 103386 4880 103388
rect 4936 103386 4960 103388
rect 5016 103386 5040 103388
rect 5096 103386 5120 103388
rect 5176 103386 5182 103388
rect 4936 103334 4938 103386
rect 5118 103334 5120 103386
rect 4874 103332 4880 103334
rect 4936 103332 4960 103334
rect 5016 103332 5040 103334
rect 5096 103332 5120 103334
rect 5176 103332 5182 103334
rect 4874 103323 5182 103332
rect 4214 102844 4522 102853
rect 4214 102842 4220 102844
rect 4276 102842 4300 102844
rect 4356 102842 4380 102844
rect 4436 102842 4460 102844
rect 4516 102842 4522 102844
rect 4276 102790 4278 102842
rect 4458 102790 4460 102842
rect 4214 102788 4220 102790
rect 4276 102788 4300 102790
rect 4356 102788 4380 102790
rect 4436 102788 4460 102790
rect 4516 102788 4522 102790
rect 4214 102779 4522 102788
rect 4874 102300 5182 102309
rect 4874 102298 4880 102300
rect 4936 102298 4960 102300
rect 5016 102298 5040 102300
rect 5096 102298 5120 102300
rect 5176 102298 5182 102300
rect 4936 102246 4938 102298
rect 5118 102246 5120 102298
rect 4874 102244 4880 102246
rect 4936 102244 4960 102246
rect 5016 102244 5040 102246
rect 5096 102244 5120 102246
rect 5176 102244 5182 102246
rect 4874 102235 5182 102244
rect 4214 101756 4522 101765
rect 4214 101754 4220 101756
rect 4276 101754 4300 101756
rect 4356 101754 4380 101756
rect 4436 101754 4460 101756
rect 4516 101754 4522 101756
rect 4276 101702 4278 101754
rect 4458 101702 4460 101754
rect 4214 101700 4220 101702
rect 4276 101700 4300 101702
rect 4356 101700 4380 101702
rect 4436 101700 4460 101702
rect 4516 101700 4522 101702
rect 4214 101691 4522 101700
rect 4874 101212 5182 101221
rect 4874 101210 4880 101212
rect 4936 101210 4960 101212
rect 5016 101210 5040 101212
rect 5096 101210 5120 101212
rect 5176 101210 5182 101212
rect 4936 101158 4938 101210
rect 5118 101158 5120 101210
rect 4874 101156 4880 101158
rect 4936 101156 4960 101158
rect 5016 101156 5040 101158
rect 5096 101156 5120 101158
rect 5176 101156 5182 101158
rect 4874 101147 5182 101156
rect 4214 100668 4522 100677
rect 4214 100666 4220 100668
rect 4276 100666 4300 100668
rect 4356 100666 4380 100668
rect 4436 100666 4460 100668
rect 4516 100666 4522 100668
rect 4276 100614 4278 100666
rect 4458 100614 4460 100666
rect 4214 100612 4220 100614
rect 4276 100612 4300 100614
rect 4356 100612 4380 100614
rect 4436 100612 4460 100614
rect 4516 100612 4522 100614
rect 4214 100603 4522 100612
rect 4874 100124 5182 100133
rect 4874 100122 4880 100124
rect 4936 100122 4960 100124
rect 5016 100122 5040 100124
rect 5096 100122 5120 100124
rect 5176 100122 5182 100124
rect 4936 100070 4938 100122
rect 5118 100070 5120 100122
rect 4874 100068 4880 100070
rect 4936 100068 4960 100070
rect 5016 100068 5040 100070
rect 5096 100068 5120 100070
rect 5176 100068 5182 100070
rect 4874 100059 5182 100068
rect 4214 99580 4522 99589
rect 4214 99578 4220 99580
rect 4276 99578 4300 99580
rect 4356 99578 4380 99580
rect 4436 99578 4460 99580
rect 4516 99578 4522 99580
rect 4276 99526 4278 99578
rect 4458 99526 4460 99578
rect 4214 99524 4220 99526
rect 4276 99524 4300 99526
rect 4356 99524 4380 99526
rect 4436 99524 4460 99526
rect 4516 99524 4522 99526
rect 4214 99515 4522 99524
rect 4874 99036 5182 99045
rect 4874 99034 4880 99036
rect 4936 99034 4960 99036
rect 5016 99034 5040 99036
rect 5096 99034 5120 99036
rect 5176 99034 5182 99036
rect 4936 98982 4938 99034
rect 5118 98982 5120 99034
rect 4874 98980 4880 98982
rect 4936 98980 4960 98982
rect 5016 98980 5040 98982
rect 5096 98980 5120 98982
rect 5176 98980 5182 98982
rect 4874 98971 5182 98980
rect 4214 98492 4522 98501
rect 4214 98490 4220 98492
rect 4276 98490 4300 98492
rect 4356 98490 4380 98492
rect 4436 98490 4460 98492
rect 4516 98490 4522 98492
rect 4276 98438 4278 98490
rect 4458 98438 4460 98490
rect 4214 98436 4220 98438
rect 4276 98436 4300 98438
rect 4356 98436 4380 98438
rect 4436 98436 4460 98438
rect 4516 98436 4522 98438
rect 4214 98427 4522 98436
rect 4874 97948 5182 97957
rect 4874 97946 4880 97948
rect 4936 97946 4960 97948
rect 5016 97946 5040 97948
rect 5096 97946 5120 97948
rect 5176 97946 5182 97948
rect 4936 97894 4938 97946
rect 5118 97894 5120 97946
rect 4874 97892 4880 97894
rect 4936 97892 4960 97894
rect 5016 97892 5040 97894
rect 5096 97892 5120 97894
rect 5176 97892 5182 97894
rect 4874 97883 5182 97892
rect 4214 97404 4522 97413
rect 4214 97402 4220 97404
rect 4276 97402 4300 97404
rect 4356 97402 4380 97404
rect 4436 97402 4460 97404
rect 4516 97402 4522 97404
rect 4276 97350 4278 97402
rect 4458 97350 4460 97402
rect 4214 97348 4220 97350
rect 4276 97348 4300 97350
rect 4356 97348 4380 97350
rect 4436 97348 4460 97350
rect 4516 97348 4522 97350
rect 4214 97339 4522 97348
rect 4874 96860 5182 96869
rect 4874 96858 4880 96860
rect 4936 96858 4960 96860
rect 5016 96858 5040 96860
rect 5096 96858 5120 96860
rect 5176 96858 5182 96860
rect 4936 96806 4938 96858
rect 5118 96806 5120 96858
rect 4874 96804 4880 96806
rect 4936 96804 4960 96806
rect 5016 96804 5040 96806
rect 5096 96804 5120 96806
rect 5176 96804 5182 96806
rect 4874 96795 5182 96804
rect 4214 96316 4522 96325
rect 4214 96314 4220 96316
rect 4276 96314 4300 96316
rect 4356 96314 4380 96316
rect 4436 96314 4460 96316
rect 4516 96314 4522 96316
rect 4276 96262 4278 96314
rect 4458 96262 4460 96314
rect 4214 96260 4220 96262
rect 4276 96260 4300 96262
rect 4356 96260 4380 96262
rect 4436 96260 4460 96262
rect 4516 96260 4522 96262
rect 4214 96251 4522 96260
rect 4874 95772 5182 95781
rect 4874 95770 4880 95772
rect 4936 95770 4960 95772
rect 5016 95770 5040 95772
rect 5096 95770 5120 95772
rect 5176 95770 5182 95772
rect 4936 95718 4938 95770
rect 5118 95718 5120 95770
rect 4874 95716 4880 95718
rect 4936 95716 4960 95718
rect 5016 95716 5040 95718
rect 5096 95716 5120 95718
rect 5176 95716 5182 95718
rect 4874 95707 5182 95716
rect 4214 95228 4522 95237
rect 4214 95226 4220 95228
rect 4276 95226 4300 95228
rect 4356 95226 4380 95228
rect 4436 95226 4460 95228
rect 4516 95226 4522 95228
rect 4276 95174 4278 95226
rect 4458 95174 4460 95226
rect 4214 95172 4220 95174
rect 4276 95172 4300 95174
rect 4356 95172 4380 95174
rect 4436 95172 4460 95174
rect 4516 95172 4522 95174
rect 4214 95163 4522 95172
rect 4874 94684 5182 94693
rect 4874 94682 4880 94684
rect 4936 94682 4960 94684
rect 5016 94682 5040 94684
rect 5096 94682 5120 94684
rect 5176 94682 5182 94684
rect 4936 94630 4938 94682
rect 5118 94630 5120 94682
rect 4874 94628 4880 94630
rect 4936 94628 4960 94630
rect 5016 94628 5040 94630
rect 5096 94628 5120 94630
rect 5176 94628 5182 94630
rect 4874 94619 5182 94628
rect 4214 94140 4522 94149
rect 4214 94138 4220 94140
rect 4276 94138 4300 94140
rect 4356 94138 4380 94140
rect 4436 94138 4460 94140
rect 4516 94138 4522 94140
rect 4276 94086 4278 94138
rect 4458 94086 4460 94138
rect 4214 94084 4220 94086
rect 4276 94084 4300 94086
rect 4356 94084 4380 94086
rect 4436 94084 4460 94086
rect 4516 94084 4522 94086
rect 4214 94075 4522 94084
rect 4874 93596 5182 93605
rect 4874 93594 4880 93596
rect 4936 93594 4960 93596
rect 5016 93594 5040 93596
rect 5096 93594 5120 93596
rect 5176 93594 5182 93596
rect 4936 93542 4938 93594
rect 5118 93542 5120 93594
rect 4874 93540 4880 93542
rect 4936 93540 4960 93542
rect 5016 93540 5040 93542
rect 5096 93540 5120 93542
rect 5176 93540 5182 93542
rect 4874 93531 5182 93540
rect 4214 93052 4522 93061
rect 4214 93050 4220 93052
rect 4276 93050 4300 93052
rect 4356 93050 4380 93052
rect 4436 93050 4460 93052
rect 4516 93050 4522 93052
rect 4276 92998 4278 93050
rect 4458 92998 4460 93050
rect 4214 92996 4220 92998
rect 4276 92996 4300 92998
rect 4356 92996 4380 92998
rect 4436 92996 4460 92998
rect 4516 92996 4522 92998
rect 4214 92987 4522 92996
rect 4874 92508 5182 92517
rect 4874 92506 4880 92508
rect 4936 92506 4960 92508
rect 5016 92506 5040 92508
rect 5096 92506 5120 92508
rect 5176 92506 5182 92508
rect 4936 92454 4938 92506
rect 5118 92454 5120 92506
rect 4874 92452 4880 92454
rect 4936 92452 4960 92454
rect 5016 92452 5040 92454
rect 5096 92452 5120 92454
rect 5176 92452 5182 92454
rect 4874 92443 5182 92452
rect 4214 91964 4522 91973
rect 4214 91962 4220 91964
rect 4276 91962 4300 91964
rect 4356 91962 4380 91964
rect 4436 91962 4460 91964
rect 4516 91962 4522 91964
rect 4276 91910 4278 91962
rect 4458 91910 4460 91962
rect 4214 91908 4220 91910
rect 4276 91908 4300 91910
rect 4356 91908 4380 91910
rect 4436 91908 4460 91910
rect 4516 91908 4522 91910
rect 4214 91899 4522 91908
rect 4874 91420 5182 91429
rect 4874 91418 4880 91420
rect 4936 91418 4960 91420
rect 5016 91418 5040 91420
rect 5096 91418 5120 91420
rect 5176 91418 5182 91420
rect 4936 91366 4938 91418
rect 5118 91366 5120 91418
rect 4874 91364 4880 91366
rect 4936 91364 4960 91366
rect 5016 91364 5040 91366
rect 5096 91364 5120 91366
rect 5176 91364 5182 91366
rect 4874 91355 5182 91364
rect 4214 90876 4522 90885
rect 4214 90874 4220 90876
rect 4276 90874 4300 90876
rect 4356 90874 4380 90876
rect 4436 90874 4460 90876
rect 4516 90874 4522 90876
rect 4276 90822 4278 90874
rect 4458 90822 4460 90874
rect 4214 90820 4220 90822
rect 4276 90820 4300 90822
rect 4356 90820 4380 90822
rect 4436 90820 4460 90822
rect 4516 90820 4522 90822
rect 4214 90811 4522 90820
rect 4874 90332 5182 90341
rect 4874 90330 4880 90332
rect 4936 90330 4960 90332
rect 5016 90330 5040 90332
rect 5096 90330 5120 90332
rect 5176 90330 5182 90332
rect 4936 90278 4938 90330
rect 5118 90278 5120 90330
rect 4874 90276 4880 90278
rect 4936 90276 4960 90278
rect 5016 90276 5040 90278
rect 5096 90276 5120 90278
rect 5176 90276 5182 90278
rect 4874 90267 5182 90276
rect 4214 89788 4522 89797
rect 4214 89786 4220 89788
rect 4276 89786 4300 89788
rect 4356 89786 4380 89788
rect 4436 89786 4460 89788
rect 4516 89786 4522 89788
rect 4276 89734 4278 89786
rect 4458 89734 4460 89786
rect 4214 89732 4220 89734
rect 4276 89732 4300 89734
rect 4356 89732 4380 89734
rect 4436 89732 4460 89734
rect 4516 89732 4522 89734
rect 4214 89723 4522 89732
rect 4874 89244 5182 89253
rect 4874 89242 4880 89244
rect 4936 89242 4960 89244
rect 5016 89242 5040 89244
rect 5096 89242 5120 89244
rect 5176 89242 5182 89244
rect 4936 89190 4938 89242
rect 5118 89190 5120 89242
rect 4874 89188 4880 89190
rect 4936 89188 4960 89190
rect 5016 89188 5040 89190
rect 5096 89188 5120 89190
rect 5176 89188 5182 89190
rect 4874 89179 5182 89188
rect 1308 89004 1360 89010
rect 1308 88946 1360 88952
rect 1320 88505 1348 88946
rect 7564 88868 7616 88874
rect 7564 88810 7616 88816
rect 4214 88700 4522 88709
rect 4214 88698 4220 88700
rect 4276 88698 4300 88700
rect 4356 88698 4380 88700
rect 4436 88698 4460 88700
rect 4516 88698 4522 88700
rect 4276 88646 4278 88698
rect 4458 88646 4460 88698
rect 4214 88644 4220 88646
rect 4276 88644 4300 88646
rect 4356 88644 4380 88646
rect 4436 88644 4460 88646
rect 4516 88644 4522 88646
rect 4214 88635 4522 88644
rect 1306 88496 1362 88505
rect 1306 88431 1362 88440
rect 4874 88156 5182 88165
rect 4874 88154 4880 88156
rect 4936 88154 4960 88156
rect 5016 88154 5040 88156
rect 5096 88154 5120 88156
rect 5176 88154 5182 88156
rect 4936 88102 4938 88154
rect 5118 88102 5120 88154
rect 4874 88100 4880 88102
rect 4936 88100 4960 88102
rect 5016 88100 5040 88102
rect 5096 88100 5120 88102
rect 5176 88100 5182 88102
rect 4874 88091 5182 88100
rect 1216 87916 1268 87922
rect 1216 87858 1268 87864
rect 1228 87825 1256 87858
rect 1214 87816 1270 87825
rect 1214 87751 1270 87760
rect 4214 87612 4522 87621
rect 4214 87610 4220 87612
rect 4276 87610 4300 87612
rect 4356 87610 4380 87612
rect 4436 87610 4460 87612
rect 4516 87610 4522 87612
rect 4276 87558 4278 87610
rect 4458 87558 4460 87610
rect 4214 87556 4220 87558
rect 4276 87556 4300 87558
rect 4356 87556 4380 87558
rect 4436 87556 4460 87558
rect 4516 87556 4522 87558
rect 4214 87547 4522 87556
rect 1216 87236 1268 87242
rect 1216 87178 1268 87184
rect 1228 87145 1256 87178
rect 1860 87168 1912 87174
rect 1214 87136 1270 87145
rect 1860 87110 1912 87116
rect 1214 87071 1270 87080
rect 1308 86828 1360 86834
rect 1308 86770 1360 86776
rect 1320 86465 1348 86770
rect 1306 86456 1362 86465
rect 1306 86391 1362 86400
rect 1308 86216 1360 86222
rect 1308 86158 1360 86164
rect 1320 85785 1348 86158
rect 1872 86154 1900 87110
rect 4874 87068 5182 87077
rect 4874 87066 4880 87068
rect 4936 87066 4960 87068
rect 5016 87066 5040 87068
rect 5096 87066 5120 87068
rect 5176 87066 5182 87068
rect 4936 87014 4938 87066
rect 5118 87014 5120 87066
rect 4874 87012 4880 87014
rect 4936 87012 4960 87014
rect 5016 87012 5040 87014
rect 5096 87012 5120 87014
rect 5176 87012 5182 87014
rect 4874 87003 5182 87012
rect 4214 86524 4522 86533
rect 4214 86522 4220 86524
rect 4276 86522 4300 86524
rect 4356 86522 4380 86524
rect 4436 86522 4460 86524
rect 4516 86522 4522 86524
rect 4276 86470 4278 86522
rect 4458 86470 4460 86522
rect 4214 86468 4220 86470
rect 4276 86468 4300 86470
rect 4356 86468 4380 86470
rect 4436 86468 4460 86470
rect 4516 86468 4522 86470
rect 4214 86459 4522 86468
rect 1860 86148 1912 86154
rect 1860 86090 1912 86096
rect 6000 86080 6052 86086
rect 6000 86022 6052 86028
rect 4874 85980 5182 85989
rect 4874 85978 4880 85980
rect 4936 85978 4960 85980
rect 5016 85978 5040 85980
rect 5096 85978 5120 85980
rect 5176 85978 5182 85980
rect 4936 85926 4938 85978
rect 5118 85926 5120 85978
rect 4874 85924 4880 85926
rect 4936 85924 4960 85926
rect 5016 85924 5040 85926
rect 5096 85924 5120 85926
rect 5176 85924 5182 85926
rect 4874 85915 5182 85924
rect 1306 85776 1362 85785
rect 1306 85711 1362 85720
rect 6012 85513 6040 86022
rect 5998 85504 6054 85513
rect 4214 85436 4522 85445
rect 5998 85439 6054 85448
rect 4214 85434 4220 85436
rect 4276 85434 4300 85436
rect 4356 85434 4380 85436
rect 4436 85434 4460 85436
rect 4516 85434 4522 85436
rect 4276 85382 4278 85434
rect 4458 85382 4460 85434
rect 4214 85380 4220 85382
rect 4276 85380 4300 85382
rect 4356 85380 4380 85382
rect 4436 85380 4460 85382
rect 4516 85380 4522 85382
rect 4214 85371 4522 85380
rect 1214 85096 1270 85105
rect 1214 85031 1216 85040
rect 1268 85031 1270 85040
rect 1216 85002 1268 85008
rect 1768 84992 1820 84998
rect 1768 84934 1820 84940
rect 1308 84652 1360 84658
rect 1308 84594 1360 84600
rect 1320 84425 1348 84594
rect 1306 84416 1362 84425
rect 1306 84351 1362 84360
rect 1780 84194 1808 84934
rect 4874 84892 5182 84901
rect 4874 84890 4880 84892
rect 4936 84890 4960 84892
rect 5016 84890 5040 84892
rect 5096 84890 5120 84892
rect 5176 84890 5182 84892
rect 4936 84838 4938 84890
rect 5118 84838 5120 84890
rect 4874 84836 4880 84838
rect 4936 84836 4960 84838
rect 5016 84836 5040 84838
rect 5096 84836 5120 84838
rect 5176 84836 5182 84838
rect 4874 84827 5182 84836
rect 1860 84516 1912 84522
rect 1860 84458 1912 84464
rect 1872 84402 1900 84458
rect 1872 84374 1992 84402
rect 1780 84166 1900 84194
rect 1964 84182 1992 84374
rect 4214 84348 4522 84357
rect 4214 84346 4220 84348
rect 4276 84346 4300 84348
rect 4356 84346 4380 84348
rect 4436 84346 4460 84348
rect 4516 84346 4522 84348
rect 4276 84294 4278 84346
rect 4458 84294 4460 84346
rect 4214 84292 4220 84294
rect 4276 84292 4300 84294
rect 4356 84292 4380 84294
rect 4436 84292 4460 84294
rect 4516 84292 4522 84294
rect 4214 84283 4522 84292
rect 1308 83972 1360 83978
rect 1308 83914 1360 83920
rect 1320 83745 1348 83914
rect 1306 83736 1362 83745
rect 1306 83671 1362 83680
rect 1308 83564 1360 83570
rect 1308 83506 1360 83512
rect 1320 83065 1348 83506
rect 1306 83056 1362 83065
rect 1306 82991 1362 83000
rect 1872 82822 1900 84166
rect 1952 84176 2004 84182
rect 1952 84118 2004 84124
rect 4874 83804 5182 83813
rect 4874 83802 4880 83804
rect 4936 83802 4960 83804
rect 5016 83802 5040 83804
rect 5096 83802 5120 83804
rect 5176 83802 5182 83804
rect 4936 83750 4938 83802
rect 5118 83750 5120 83802
rect 4874 83748 4880 83750
rect 4936 83748 4960 83750
rect 5016 83748 5040 83750
rect 5096 83748 5120 83750
rect 5176 83748 5182 83750
rect 4874 83739 5182 83748
rect 2504 83360 2556 83366
rect 2504 83302 2556 83308
rect 1860 82816 1912 82822
rect 1860 82758 1912 82764
rect 1216 82476 1268 82482
rect 1216 82418 1268 82424
rect 1228 82385 1256 82418
rect 1214 82376 1270 82385
rect 1214 82311 1270 82320
rect 2412 82272 2464 82278
rect 2412 82214 2464 82220
rect 1216 81796 1268 81802
rect 1216 81738 1268 81744
rect 1228 81705 1256 81738
rect 1860 81728 1912 81734
rect 1214 81696 1270 81705
rect 1860 81670 1912 81676
rect 1214 81631 1270 81640
rect 1308 81388 1360 81394
rect 1308 81330 1360 81336
rect 1320 81025 1348 81330
rect 1872 81258 1900 81670
rect 1860 81252 1912 81258
rect 1860 81194 1912 81200
rect 1306 81016 1362 81025
rect 1306 80951 1362 80960
rect 2424 80850 2452 82214
rect 2412 80844 2464 80850
rect 2412 80786 2464 80792
rect 1308 80776 1360 80782
rect 1308 80718 1360 80724
rect 1320 80374 1348 80718
rect 2516 80714 2544 83302
rect 4214 83260 4522 83269
rect 4214 83258 4220 83260
rect 4276 83258 4300 83260
rect 4356 83258 4380 83260
rect 4436 83258 4460 83260
rect 4516 83258 4522 83260
rect 4276 83206 4278 83258
rect 4458 83206 4460 83258
rect 4214 83204 4220 83206
rect 4276 83204 4300 83206
rect 4356 83204 4380 83206
rect 4436 83204 4460 83206
rect 4516 83204 4522 83206
rect 4214 83195 4522 83204
rect 4874 82716 5182 82725
rect 4874 82714 4880 82716
rect 4936 82714 4960 82716
rect 5016 82714 5040 82716
rect 5096 82714 5120 82716
rect 5176 82714 5182 82716
rect 4936 82662 4938 82714
rect 5118 82662 5120 82714
rect 4874 82660 4880 82662
rect 4936 82660 4960 82662
rect 5016 82660 5040 82662
rect 5096 82660 5120 82662
rect 5176 82660 5182 82662
rect 4874 82651 5182 82660
rect 4214 82172 4522 82181
rect 4214 82170 4220 82172
rect 4276 82170 4300 82172
rect 4356 82170 4380 82172
rect 4436 82170 4460 82172
rect 4516 82170 4522 82172
rect 4276 82118 4278 82170
rect 4458 82118 4460 82170
rect 4214 82116 4220 82118
rect 4276 82116 4300 82118
rect 4356 82116 4380 82118
rect 4436 82116 4460 82118
rect 4516 82116 4522 82118
rect 4214 82107 4522 82116
rect 4874 81628 5182 81637
rect 4874 81626 4880 81628
rect 4936 81626 4960 81628
rect 5016 81626 5040 81628
rect 5096 81626 5120 81628
rect 5176 81626 5182 81628
rect 4936 81574 4938 81626
rect 5118 81574 5120 81626
rect 4874 81572 4880 81574
rect 4936 81572 4960 81574
rect 5016 81572 5040 81574
rect 5096 81572 5120 81574
rect 5176 81572 5182 81574
rect 4874 81563 5182 81572
rect 5632 81184 5684 81190
rect 5632 81126 5684 81132
rect 4214 81084 4522 81093
rect 4214 81082 4220 81084
rect 4276 81082 4300 81084
rect 4356 81082 4380 81084
rect 4436 81082 4460 81084
rect 4516 81082 4522 81084
rect 4276 81030 4278 81082
rect 4458 81030 4460 81082
rect 4214 81028 4220 81030
rect 4276 81028 4300 81030
rect 4356 81028 4380 81030
rect 4436 81028 4460 81030
rect 4516 81028 4522 81030
rect 4214 81019 4522 81028
rect 2504 80708 2556 80714
rect 2504 80650 2556 80656
rect 5540 80640 5592 80646
rect 5540 80582 5592 80588
rect 4874 80540 5182 80549
rect 4874 80538 4880 80540
rect 4936 80538 4960 80540
rect 5016 80538 5040 80540
rect 5096 80538 5120 80540
rect 5176 80538 5182 80540
rect 4936 80486 4938 80538
rect 5118 80486 5120 80538
rect 4874 80484 4880 80486
rect 4936 80484 4960 80486
rect 5016 80484 5040 80486
rect 5096 80484 5120 80486
rect 5176 80484 5182 80486
rect 4874 80475 5182 80484
rect 1308 80368 1360 80374
rect 1306 80336 1308 80345
rect 1360 80336 1362 80345
rect 1306 80271 1362 80280
rect 4214 79996 4522 80005
rect 4214 79994 4220 79996
rect 4276 79994 4300 79996
rect 4356 79994 4380 79996
rect 4436 79994 4460 79996
rect 4516 79994 4522 79996
rect 4276 79942 4278 79994
rect 4458 79942 4460 79994
rect 4214 79940 4220 79942
rect 4276 79940 4300 79942
rect 4356 79940 4380 79942
rect 4436 79940 4460 79942
rect 4516 79940 4522 79942
rect 4214 79931 4522 79940
rect 1214 79656 1270 79665
rect 1214 79591 1216 79600
rect 1268 79591 1270 79600
rect 1216 79562 1268 79568
rect 5552 79529 5580 80582
rect 5644 79665 5672 81126
rect 5630 79656 5686 79665
rect 5630 79591 5686 79600
rect 5538 79520 5594 79529
rect 4874 79452 5182 79461
rect 5538 79455 5594 79464
rect 4874 79450 4880 79452
rect 4936 79450 4960 79452
rect 5016 79450 5040 79452
rect 5096 79450 5120 79452
rect 5176 79450 5182 79452
rect 4936 79398 4938 79450
rect 5118 79398 5120 79450
rect 4874 79396 4880 79398
rect 4936 79396 4960 79398
rect 5016 79396 5040 79398
rect 5096 79396 5120 79398
rect 5176 79396 5182 79398
rect 4874 79387 5182 79396
rect 7576 79257 7604 88810
rect 7562 79248 7618 79257
rect 1308 79212 1360 79218
rect 7562 79183 7618 79192
rect 1308 79154 1360 79160
rect 1320 78985 1348 79154
rect 1306 78976 1362 78985
rect 1306 78911 1362 78920
rect 4214 78908 4522 78917
rect 4214 78906 4220 78908
rect 4276 78906 4300 78908
rect 4356 78906 4380 78908
rect 4436 78906 4460 78908
rect 4516 78906 4522 78908
rect 4276 78854 4278 78906
rect 4458 78854 4460 78906
rect 4214 78852 4220 78854
rect 4276 78852 4300 78854
rect 4356 78852 4380 78854
rect 4436 78852 4460 78854
rect 4516 78852 4522 78854
rect 4214 78843 4522 78852
rect 1308 78532 1360 78538
rect 1308 78474 1360 78480
rect 1320 78305 1348 78474
rect 4874 78364 5182 78373
rect 4874 78362 4880 78364
rect 4936 78362 4960 78364
rect 5016 78362 5040 78364
rect 5096 78362 5120 78364
rect 5176 78362 5182 78364
rect 4936 78310 4938 78362
rect 5118 78310 5120 78362
rect 4874 78308 4880 78310
rect 4936 78308 4960 78310
rect 5016 78308 5040 78310
rect 5096 78308 5120 78310
rect 5176 78308 5182 78310
rect 1306 78296 1362 78305
rect 4874 78299 5182 78308
rect 1306 78231 1362 78240
rect 2320 78192 2372 78198
rect 2320 78134 2372 78140
rect 1308 78124 1360 78130
rect 1308 78066 1360 78072
rect 1320 77625 1348 78066
rect 1306 77616 1362 77625
rect 1306 77551 1362 77560
rect 1768 77172 1820 77178
rect 1768 77114 1820 77120
rect 1216 77036 1268 77042
rect 1216 76978 1268 76984
rect 1228 76945 1256 76978
rect 1214 76936 1270 76945
rect 1214 76871 1270 76880
rect 846 76392 902 76401
rect 846 76327 902 76336
rect 860 76294 888 76327
rect 848 76288 900 76294
rect 848 76230 900 76236
rect 1400 75744 1452 75750
rect 1400 75686 1452 75692
rect 1412 75585 1440 75686
rect 1398 75576 1454 75585
rect 1398 75511 1454 75520
rect 848 75200 900 75206
rect 848 75142 900 75148
rect 860 75041 888 75142
rect 846 75032 902 75041
rect 846 74967 902 74976
rect 848 74384 900 74390
rect 846 74352 848 74361
rect 900 74352 902 74361
rect 846 74287 902 74296
rect 846 73672 902 73681
rect 846 73607 848 73616
rect 900 73607 902 73616
rect 848 73578 900 73584
rect 1780 73370 1808 77114
rect 2332 76090 2360 78134
rect 4214 77820 4522 77829
rect 4214 77818 4220 77820
rect 4276 77818 4300 77820
rect 4356 77818 4380 77820
rect 4436 77818 4460 77820
rect 4516 77818 4522 77820
rect 4276 77766 4278 77818
rect 4458 77766 4460 77818
rect 4214 77764 4220 77766
rect 4276 77764 4300 77766
rect 4356 77764 4380 77766
rect 4436 77764 4460 77766
rect 4516 77764 4522 77766
rect 4214 77755 4522 77764
rect 7944 77761 7972 133894
rect 8036 78577 8064 135662
rect 8022 78568 8078 78577
rect 8022 78503 8078 78512
rect 8128 77897 8156 135866
rect 8208 135856 8260 135862
rect 8208 135798 8260 135804
rect 8220 78169 8248 135798
rect 8392 111376 8444 111382
rect 8392 111318 8444 111324
rect 8404 111217 8432 111318
rect 8390 111208 8446 111217
rect 8390 111143 8446 111152
rect 8390 109576 8446 109585
rect 8390 109511 8392 109520
rect 8444 109511 8446 109520
rect 8392 109482 8444 109488
rect 8390 108488 8446 108497
rect 8390 108423 8392 108432
rect 8444 108423 8446 108432
rect 8392 108394 8444 108400
rect 8392 107024 8444 107030
rect 8392 106966 8444 106972
rect 8404 106729 8432 106966
rect 8390 106720 8446 106729
rect 8390 106655 8446 106664
rect 8392 105936 8444 105942
rect 8392 105878 8444 105884
rect 8404 105641 8432 105878
rect 8390 105632 8446 105641
rect 8390 105567 8446 105576
rect 8392 104100 8444 104106
rect 8392 104042 8444 104048
rect 8404 104009 8432 104042
rect 8390 104000 8446 104009
rect 8390 103935 8446 103944
rect 8944 87780 8996 87786
rect 8944 87722 8996 87728
rect 8668 86692 8720 86698
rect 8668 86634 8720 86640
rect 8576 86148 8628 86154
rect 8576 86090 8628 86096
rect 8484 83972 8536 83978
rect 8484 83914 8536 83920
rect 8496 79937 8524 83914
rect 8482 79928 8538 79937
rect 8482 79863 8538 79872
rect 8588 79762 8616 86090
rect 8680 79801 8708 86634
rect 8956 79830 8984 87722
rect 9404 84176 9456 84182
rect 9404 84118 9456 84124
rect 9220 82816 9272 82822
rect 9220 82758 9272 82764
rect 8944 79824 8996 79830
rect 8666 79792 8722 79801
rect 8576 79756 8628 79762
rect 8944 79766 8996 79772
rect 8666 79727 8722 79736
rect 8576 79698 8628 79704
rect 9232 79694 9260 82758
rect 9220 79688 9272 79694
rect 9220 79630 9272 79636
rect 9416 79393 9444 84118
rect 9402 79384 9458 79393
rect 9402 79319 9458 79328
rect 8206 78160 8262 78169
rect 8206 78095 8262 78104
rect 8114 77888 8170 77897
rect 8114 77823 8170 77832
rect 7930 77752 7986 77761
rect 7930 77687 7986 77696
rect 9508 77625 9536 136070
rect 35594 136028 35902 136037
rect 35594 136026 35600 136028
rect 35656 136026 35680 136028
rect 35736 136026 35760 136028
rect 35816 136026 35840 136028
rect 35896 136026 35902 136028
rect 35656 135974 35658 136026
rect 35838 135974 35840 136026
rect 35594 135972 35600 135974
rect 35656 135972 35680 135974
rect 35736 135972 35760 135974
rect 35816 135972 35840 135974
rect 35896 135972 35902 135974
rect 35594 135963 35902 135972
rect 9588 135788 9640 135794
rect 9588 135730 9640 135736
rect 9600 78305 9628 135730
rect 36096 133958 36124 136070
rect 38120 135726 38148 136070
rect 38108 135720 38160 135726
rect 38108 135662 38160 135668
rect 38212 134201 38240 136138
rect 40592 136128 40644 136134
rect 40592 136070 40644 136076
rect 40604 135794 40632 136070
rect 40592 135788 40644 135794
rect 40592 135730 40644 135736
rect 40696 134201 40724 136138
rect 42892 136128 42944 136134
rect 42892 136070 42944 136076
rect 42904 135862 42932 136070
rect 42892 135856 42944 135862
rect 42892 135798 42944 135804
rect 38198 134192 38254 134201
rect 38198 134127 38254 134136
rect 40682 134192 40738 134201
rect 40682 134127 40738 134136
rect 36084 133952 36136 133958
rect 36082 133920 36084 133929
rect 42996 133929 43024 136138
rect 45192 136128 45244 136134
rect 45192 136070 45244 136076
rect 45204 135930 45232 136070
rect 45192 135924 45244 135930
rect 45192 135866 45244 135872
rect 46032 133929 46060 136138
rect 48516 133929 48544 136138
rect 52380 134201 52408 136138
rect 52366 134192 52422 134201
rect 52366 134127 52422 134136
rect 55784 134065 55812 136138
rect 56140 136128 56192 136134
rect 56140 136070 56192 136076
rect 56152 135930 56180 136070
rect 56140 135924 56192 135930
rect 56140 135866 56192 135872
rect 58176 134201 58204 136138
rect 58532 136128 58584 136134
rect 58532 136070 58584 136076
rect 58544 135862 58572 136070
rect 58532 135856 58584 135862
rect 58532 135798 58584 135804
rect 60660 135289 60688 136138
rect 61016 136128 61068 136134
rect 61016 136070 61068 136076
rect 61028 135794 61056 136070
rect 61016 135788 61068 135794
rect 61016 135730 61068 135736
rect 63144 135289 63172 136138
rect 63500 136128 63552 136134
rect 63500 136070 63552 136076
rect 63512 135726 63540 136070
rect 63500 135720 63552 135726
rect 63500 135662 63552 135668
rect 60646 135280 60702 135289
rect 60646 135215 60702 135224
rect 63130 135280 63186 135289
rect 63130 135215 63186 135224
rect 64432 135153 64460 136138
rect 65340 136128 65392 136134
rect 65340 136070 65392 136076
rect 65352 135658 65380 136070
rect 66314 136028 66622 136037
rect 66314 136026 66320 136028
rect 66376 136026 66400 136028
rect 66456 136026 66480 136028
rect 66536 136026 66560 136028
rect 66616 136026 66622 136028
rect 66376 135974 66378 136026
rect 66558 135974 66560 136026
rect 66314 135972 66320 135974
rect 66376 135972 66400 135974
rect 66456 135972 66480 135974
rect 66536 135972 66560 135974
rect 66616 135972 66622 135974
rect 66314 135963 66622 135972
rect 65340 135652 65392 135658
rect 65340 135594 65392 135600
rect 67560 135289 67588 136138
rect 67916 136128 67968 136134
rect 67916 136070 67968 136076
rect 67928 135590 67956 136070
rect 67916 135584 67968 135590
rect 67916 135526 67968 135532
rect 69768 135289 69796 136138
rect 70124 136128 70176 136134
rect 70124 136070 70176 136076
rect 70136 135522 70164 136070
rect 70124 135516 70176 135522
rect 70124 135458 70176 135464
rect 72160 135289 72188 136138
rect 72516 136128 72568 136134
rect 72516 136070 72568 136076
rect 72528 135454 72556 136070
rect 72516 135448 72568 135454
rect 72516 135390 72568 135396
rect 67546 135280 67602 135289
rect 67546 135215 67602 135224
rect 69754 135280 69810 135289
rect 69754 135215 69810 135224
rect 72146 135280 72202 135289
rect 72146 135215 72202 135224
rect 64418 135144 64474 135153
rect 64418 135079 64474 135088
rect 74184 134201 74212 136138
rect 77760 136128 77812 136134
rect 77760 136070 77812 136076
rect 86132 136128 86184 136134
rect 86132 136070 86184 136076
rect 87328 136128 87380 136134
rect 87328 136070 87380 136076
rect 95976 136128 96028 136134
rect 95976 136070 96028 136076
rect 77772 135386 77800 136070
rect 77760 135380 77812 135386
rect 77760 135322 77812 135328
rect 58162 134192 58218 134201
rect 58162 134127 58218 134136
rect 74170 134192 74226 134201
rect 74170 134127 74226 134136
rect 55770 134056 55826 134065
rect 55770 133991 55826 134000
rect 86144 133958 86172 136070
rect 87340 134026 87368 136070
rect 95988 134570 96016 136070
rect 97034 136028 97342 136037
rect 97034 136026 97040 136028
rect 97096 136026 97120 136028
rect 97176 136026 97200 136028
rect 97256 136026 97280 136028
rect 97336 136026 97342 136028
rect 97096 135974 97098 136026
rect 97278 135974 97280 136026
rect 97034 135972 97040 135974
rect 97096 135972 97120 135974
rect 97176 135972 97200 135974
rect 97256 135972 97280 135974
rect 97336 135972 97342 135974
rect 97034 135963 97342 135972
rect 95976 134564 96028 134570
rect 95976 134506 96028 134512
rect 95988 134473 96016 134506
rect 95974 134464 96030 134473
rect 95974 134399 96030 134408
rect 87328 134020 87380 134026
rect 87328 133962 87380 133968
rect 86132 133952 86184 133958
rect 36136 133920 36138 133929
rect 36082 133855 36138 133864
rect 42982 133920 43038 133929
rect 42982 133855 43038 133864
rect 46018 133920 46074 133929
rect 46018 133855 46074 133864
rect 48502 133920 48558 133929
rect 48502 133855 48558 133864
rect 86130 133920 86132 133929
rect 87340 133929 87368 133962
rect 86184 133920 86186 133929
rect 86130 133855 86186 133864
rect 87326 133920 87382 133929
rect 87326 133855 87382 133864
rect 9772 81252 9824 81258
rect 9772 81194 9824 81200
rect 9784 79898 9812 81194
rect 9864 80844 9916 80850
rect 9864 80786 9916 80792
rect 9876 79966 9904 80786
rect 9956 80708 10008 80714
rect 9956 80650 10008 80656
rect 9968 80034 9996 80650
rect 9956 80028 10008 80034
rect 9956 79970 10008 79976
rect 40960 80028 41012 80034
rect 40960 79970 41012 79976
rect 9864 79960 9916 79966
rect 39764 79960 39816 79966
rect 9864 79902 9916 79908
rect 36266 79928 36322 79937
rect 9772 79892 9824 79898
rect 36266 79863 36322 79872
rect 38658 79928 38714 79937
rect 38658 79863 38660 79872
rect 9772 79834 9824 79840
rect 36280 79830 36308 79863
rect 38712 79863 38714 79872
rect 39762 79928 39764 79937
rect 40972 79937 41000 79970
rect 39816 79928 39818 79937
rect 39762 79863 39818 79872
rect 40958 79928 41014 79937
rect 40958 79863 41014 79872
rect 90638 79928 90694 79937
rect 90638 79863 90694 79872
rect 38660 79834 38712 79840
rect 36268 79824 36320 79830
rect 32310 79792 32366 79801
rect 36268 79766 36320 79772
rect 32310 79727 32366 79736
rect 34704 79756 34756 79762
rect 32324 79694 32352 79727
rect 34704 79698 34756 79704
rect 32312 79688 32364 79694
rect 27618 79656 27674 79665
rect 32312 79630 32364 79636
rect 27618 79591 27674 79600
rect 24674 79520 24730 79529
rect 24674 79455 24730 79464
rect 22744 78328 22796 78334
rect 9586 78296 9642 78305
rect 22744 78270 22796 78276
rect 9586 78231 9642 78240
rect 22100 78260 22152 78266
rect 22100 78202 22152 78208
rect 20812 78056 20864 78062
rect 16026 78024 16082 78033
rect 20812 77998 20864 78004
rect 16026 77959 16082 77968
rect 9494 77616 9550 77625
rect 9494 77551 9550 77560
rect 16040 77382 16068 77959
rect 17868 77648 17920 77654
rect 17868 77590 17920 77596
rect 6828 77376 6880 77382
rect 6828 77318 6880 77324
rect 16028 77376 16080 77382
rect 16028 77318 16080 77324
rect 4874 77276 5182 77285
rect 4874 77274 4880 77276
rect 4936 77274 4960 77276
rect 5016 77274 5040 77276
rect 5096 77274 5120 77276
rect 5176 77274 5182 77276
rect 4936 77222 4938 77274
rect 5118 77222 5120 77274
rect 4874 77220 4880 77222
rect 4936 77220 4960 77222
rect 5016 77220 5040 77222
rect 5096 77220 5120 77222
rect 5176 77220 5182 77222
rect 4874 77211 5182 77220
rect 4214 76732 4522 76741
rect 4214 76730 4220 76732
rect 4276 76730 4300 76732
rect 4356 76730 4380 76732
rect 4436 76730 4460 76732
rect 4516 76730 4522 76732
rect 4276 76678 4278 76730
rect 4458 76678 4460 76730
rect 4214 76676 4220 76678
rect 4276 76676 4300 76678
rect 4356 76676 4380 76678
rect 4436 76676 4460 76678
rect 4516 76676 4522 76678
rect 4214 76667 4522 76676
rect 4874 76188 5182 76197
rect 4874 76186 4880 76188
rect 4936 76186 4960 76188
rect 5016 76186 5040 76188
rect 5096 76186 5120 76188
rect 5176 76186 5182 76188
rect 4936 76134 4938 76186
rect 5118 76134 5120 76186
rect 4874 76132 4880 76134
rect 4936 76132 4960 76134
rect 5016 76132 5040 76134
rect 5096 76132 5120 76134
rect 5176 76132 5182 76134
rect 4874 76123 5182 76132
rect 2320 76084 2372 76090
rect 2320 76026 2372 76032
rect 4214 75644 4522 75653
rect 4214 75642 4220 75644
rect 4276 75642 4300 75644
rect 4356 75642 4380 75644
rect 4436 75642 4460 75644
rect 4516 75642 4522 75644
rect 4276 75590 4278 75642
rect 4458 75590 4460 75642
rect 4214 75588 4220 75590
rect 4276 75588 4300 75590
rect 4356 75588 4380 75590
rect 4436 75588 4460 75590
rect 4516 75588 4522 75590
rect 4214 75579 4522 75588
rect 4874 75100 5182 75109
rect 4874 75098 4880 75100
rect 4936 75098 4960 75100
rect 5016 75098 5040 75100
rect 5096 75098 5120 75100
rect 5176 75098 5182 75100
rect 4936 75046 4938 75098
rect 5118 75046 5120 75098
rect 4874 75044 4880 75046
rect 4936 75044 4960 75046
rect 5016 75044 5040 75046
rect 5096 75044 5120 75046
rect 5176 75044 5182 75046
rect 4874 75035 5182 75044
rect 4214 74556 4522 74565
rect 4214 74554 4220 74556
rect 4276 74554 4300 74556
rect 4356 74554 4380 74556
rect 4436 74554 4460 74556
rect 4516 74554 4522 74556
rect 4276 74502 4278 74554
rect 4458 74502 4460 74554
rect 4214 74500 4220 74502
rect 4276 74500 4300 74502
rect 4356 74500 4380 74502
rect 4436 74500 4460 74502
rect 4516 74500 4522 74502
rect 4214 74491 4522 74500
rect 4874 74012 5182 74021
rect 4874 74010 4880 74012
rect 4936 74010 4960 74012
rect 5016 74010 5040 74012
rect 5096 74010 5120 74012
rect 5176 74010 5182 74012
rect 4936 73958 4938 74010
rect 5118 73958 5120 74010
rect 4874 73956 4880 73958
rect 4936 73956 4960 73958
rect 5016 73956 5040 73958
rect 5096 73956 5120 73958
rect 5176 73956 5182 73958
rect 4874 73947 5182 73956
rect 4214 73468 4522 73477
rect 4214 73466 4220 73468
rect 4276 73466 4300 73468
rect 4356 73466 4380 73468
rect 4436 73466 4460 73468
rect 4516 73466 4522 73468
rect 4276 73414 4278 73466
rect 4458 73414 4460 73466
rect 4214 73412 4220 73414
rect 4276 73412 4300 73414
rect 4356 73412 4380 73414
rect 4436 73412 4460 73414
rect 4516 73412 4522 73414
rect 4214 73403 4522 73412
rect 1768 73364 1820 73370
rect 1768 73306 1820 73312
rect 1780 73166 1808 73306
rect 1768 73160 1820 73166
rect 1768 73102 1820 73108
rect 848 73024 900 73030
rect 846 72992 848 73001
rect 900 72992 902 73001
rect 846 72927 902 72936
rect 4874 72924 5182 72933
rect 4874 72922 4880 72924
rect 4936 72922 4960 72924
rect 5016 72922 5040 72924
rect 5096 72922 5120 72924
rect 5176 72922 5182 72924
rect 4936 72870 4938 72922
rect 5118 72870 5120 72922
rect 4874 72868 4880 72870
rect 4936 72868 4960 72870
rect 5016 72868 5040 72870
rect 5096 72868 5120 72870
rect 5176 72868 5182 72870
rect 4874 72859 5182 72868
rect 1124 72684 1176 72690
rect 1124 72626 1176 72632
rect 1136 72185 1164 72626
rect 4214 72380 4522 72389
rect 4214 72378 4220 72380
rect 4276 72378 4300 72380
rect 4356 72378 4380 72380
rect 4436 72378 4460 72380
rect 4516 72378 4522 72380
rect 4276 72326 4278 72378
rect 4458 72326 4460 72378
rect 4214 72324 4220 72326
rect 4276 72324 4300 72326
rect 4356 72324 4380 72326
rect 4436 72324 4460 72326
rect 4516 72324 4522 72326
rect 4214 72315 4522 72324
rect 1122 72176 1178 72185
rect 1122 72111 1178 72120
rect 4874 71836 5182 71845
rect 4874 71834 4880 71836
rect 4936 71834 4960 71836
rect 5016 71834 5040 71836
rect 5096 71834 5120 71836
rect 5176 71834 5182 71836
rect 4936 71782 4938 71834
rect 5118 71782 5120 71834
rect 4874 71780 4880 71782
rect 4936 71780 4960 71782
rect 5016 71780 5040 71782
rect 5096 71780 5120 71782
rect 5176 71780 5182 71782
rect 4874 71771 5182 71780
rect 4214 71292 4522 71301
rect 4214 71290 4220 71292
rect 4276 71290 4300 71292
rect 4356 71290 4380 71292
rect 4436 71290 4460 71292
rect 4516 71290 4522 71292
rect 4276 71238 4278 71290
rect 4458 71238 4460 71290
rect 4214 71236 4220 71238
rect 4276 71236 4300 71238
rect 4356 71236 4380 71238
rect 4436 71236 4460 71238
rect 4516 71236 4522 71238
rect 4214 71227 4522 71236
rect 4874 70748 5182 70757
rect 4874 70746 4880 70748
rect 4936 70746 4960 70748
rect 5016 70746 5040 70748
rect 5096 70746 5120 70748
rect 5176 70746 5182 70748
rect 4936 70694 4938 70746
rect 5118 70694 5120 70746
rect 4874 70692 4880 70694
rect 4936 70692 4960 70694
rect 5016 70692 5040 70694
rect 5096 70692 5120 70694
rect 5176 70692 5182 70694
rect 4874 70683 5182 70692
rect 4214 70204 4522 70213
rect 4214 70202 4220 70204
rect 4276 70202 4300 70204
rect 4356 70202 4380 70204
rect 4436 70202 4460 70204
rect 4516 70202 4522 70204
rect 4276 70150 4278 70202
rect 4458 70150 4460 70202
rect 4214 70148 4220 70150
rect 4276 70148 4300 70150
rect 4356 70148 4380 70150
rect 4436 70148 4460 70150
rect 4516 70148 4522 70150
rect 4214 70139 4522 70148
rect 4874 69660 5182 69669
rect 4874 69658 4880 69660
rect 4936 69658 4960 69660
rect 5016 69658 5040 69660
rect 5096 69658 5120 69660
rect 5176 69658 5182 69660
rect 4936 69606 4938 69658
rect 5118 69606 5120 69658
rect 4874 69604 4880 69606
rect 4936 69604 4960 69606
rect 5016 69604 5040 69606
rect 5096 69604 5120 69606
rect 5176 69604 5182 69606
rect 4874 69595 5182 69604
rect 4214 69116 4522 69125
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69051 4522 69060
rect 4874 68572 5182 68581
rect 4874 68570 4880 68572
rect 4936 68570 4960 68572
rect 5016 68570 5040 68572
rect 5096 68570 5120 68572
rect 5176 68570 5182 68572
rect 4936 68518 4938 68570
rect 5118 68518 5120 68570
rect 4874 68516 4880 68518
rect 4936 68516 4960 68518
rect 5016 68516 5040 68518
rect 5096 68516 5120 68518
rect 5176 68516 5182 68518
rect 4874 68507 5182 68516
rect 4214 68028 4522 68037
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67963 4522 67972
rect 4874 67484 5182 67493
rect 4874 67482 4880 67484
rect 4936 67482 4960 67484
rect 5016 67482 5040 67484
rect 5096 67482 5120 67484
rect 5176 67482 5182 67484
rect 4936 67430 4938 67482
rect 5118 67430 5120 67482
rect 4874 67428 4880 67430
rect 4936 67428 4960 67430
rect 5016 67428 5040 67430
rect 5096 67428 5120 67430
rect 5176 67428 5182 67430
rect 4874 67419 5182 67428
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 4874 66396 5182 66405
rect 4874 66394 4880 66396
rect 4936 66394 4960 66396
rect 5016 66394 5040 66396
rect 5096 66394 5120 66396
rect 5176 66394 5182 66396
rect 4936 66342 4938 66394
rect 5118 66342 5120 66394
rect 4874 66340 4880 66342
rect 4936 66340 4960 66342
rect 5016 66340 5040 66342
rect 5096 66340 5120 66342
rect 5176 66340 5182 66342
rect 4874 66331 5182 66340
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 4874 65308 5182 65317
rect 4874 65306 4880 65308
rect 4936 65306 4960 65308
rect 5016 65306 5040 65308
rect 5096 65306 5120 65308
rect 5176 65306 5182 65308
rect 4936 65254 4938 65306
rect 5118 65254 5120 65306
rect 4874 65252 4880 65254
rect 4936 65252 4960 65254
rect 5016 65252 5040 65254
rect 5096 65252 5120 65254
rect 5176 65252 5182 65254
rect 4874 65243 5182 65252
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 4874 64220 5182 64229
rect 4874 64218 4880 64220
rect 4936 64218 4960 64220
rect 5016 64218 5040 64220
rect 5096 64218 5120 64220
rect 5176 64218 5182 64220
rect 4936 64166 4938 64218
rect 5118 64166 5120 64218
rect 4874 64164 4880 64166
rect 4936 64164 4960 64166
rect 5016 64164 5040 64166
rect 5096 64164 5120 64166
rect 5176 64164 5182 64166
rect 4874 64155 5182 64164
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 4874 63132 5182 63141
rect 4874 63130 4880 63132
rect 4936 63130 4960 63132
rect 5016 63130 5040 63132
rect 5096 63130 5120 63132
rect 5176 63130 5182 63132
rect 4936 63078 4938 63130
rect 5118 63078 5120 63130
rect 4874 63076 4880 63078
rect 4936 63076 4960 63078
rect 5016 63076 5040 63078
rect 5096 63076 5120 63078
rect 5176 63076 5182 63078
rect 4874 63067 5182 63076
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 4874 62044 5182 62053
rect 4874 62042 4880 62044
rect 4936 62042 4960 62044
rect 5016 62042 5040 62044
rect 5096 62042 5120 62044
rect 5176 62042 5182 62044
rect 4936 61990 4938 62042
rect 5118 61990 5120 62042
rect 4874 61988 4880 61990
rect 4936 61988 4960 61990
rect 5016 61988 5040 61990
rect 5096 61988 5120 61990
rect 5176 61988 5182 61990
rect 4874 61979 5182 61988
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 4874 60956 5182 60965
rect 4874 60954 4880 60956
rect 4936 60954 4960 60956
rect 5016 60954 5040 60956
rect 5096 60954 5120 60956
rect 5176 60954 5182 60956
rect 4936 60902 4938 60954
rect 5118 60902 5120 60954
rect 4874 60900 4880 60902
rect 4936 60900 4960 60902
rect 5016 60900 5040 60902
rect 5096 60900 5120 60902
rect 5176 60900 5182 60902
rect 4874 60891 5182 60900
rect 6840 60654 6868 77318
rect 17880 76430 17908 77590
rect 20824 77450 20852 77998
rect 21272 77988 21324 77994
rect 21272 77930 21324 77936
rect 21284 77450 21312 77930
rect 21548 77580 21600 77586
rect 21548 77522 21600 77528
rect 20812 77444 20864 77450
rect 20812 77386 20864 77392
rect 21272 77444 21324 77450
rect 21272 77386 21324 77392
rect 21364 77376 21416 77382
rect 21364 77318 21416 77324
rect 17868 76424 17920 76430
rect 17868 76366 17920 76372
rect 21376 73778 21404 77318
rect 21560 76634 21588 77522
rect 22008 76900 22060 76906
rect 22008 76842 22060 76848
rect 21548 76628 21600 76634
rect 21548 76570 21600 76576
rect 22020 75206 22048 76842
rect 22112 76838 22140 78202
rect 22756 77586 22784 78270
rect 24688 77654 24716 79455
rect 26790 79384 26846 79393
rect 26790 79319 26846 79328
rect 24766 78840 24822 78849
rect 24766 78775 24822 78784
rect 24780 77654 24808 78775
rect 26056 78260 26108 78266
rect 26056 78202 26108 78208
rect 25044 78124 25096 78130
rect 25044 78066 25096 78072
rect 25056 77654 25084 78066
rect 24676 77648 24728 77654
rect 24676 77590 24728 77596
rect 24768 77648 24820 77654
rect 24768 77590 24820 77596
rect 25044 77648 25096 77654
rect 25044 77590 25096 77596
rect 22744 77580 22796 77586
rect 22744 77522 22796 77528
rect 26068 77450 26096 78202
rect 26804 77654 26832 79319
rect 27252 78056 27304 78062
rect 27252 77998 27304 78004
rect 26792 77648 26844 77654
rect 26792 77590 26844 77596
rect 26792 77512 26844 77518
rect 26792 77454 26844 77460
rect 26056 77444 26108 77450
rect 26056 77386 26108 77392
rect 23480 77172 23532 77178
rect 23480 77114 23532 77120
rect 22100 76832 22152 76838
rect 22100 76774 22152 76780
rect 22836 76832 22888 76838
rect 22836 76774 22888 76780
rect 22848 76514 22876 76774
rect 23492 76634 23520 77114
rect 24768 77104 24820 77110
rect 24768 77046 24820 77052
rect 24308 76968 24360 76974
rect 24308 76910 24360 76916
rect 24584 76968 24636 76974
rect 24584 76910 24636 76916
rect 23480 76628 23532 76634
rect 23480 76570 23532 76576
rect 23020 76560 23072 76566
rect 22848 76508 23020 76514
rect 22848 76502 23072 76508
rect 22848 76486 23060 76502
rect 22008 75200 22060 75206
rect 22008 75142 22060 75148
rect 22848 74254 22876 76486
rect 24320 76022 24348 76910
rect 24596 76634 24624 76910
rect 24584 76628 24636 76634
rect 24584 76570 24636 76576
rect 24780 76566 24808 77046
rect 26804 77042 26832 77454
rect 27264 77178 27292 77998
rect 27632 77722 27660 79591
rect 29550 79520 29606 79529
rect 29550 79455 29606 79464
rect 30470 79520 30526 79529
rect 30470 79455 30526 79464
rect 31574 79520 31630 79529
rect 31574 79455 31630 79464
rect 29564 78470 29592 79455
rect 29552 78464 29604 78470
rect 29552 78406 29604 78412
rect 28170 77752 28226 77761
rect 27528 77716 27580 77722
rect 27528 77658 27580 77664
rect 27620 77716 27672 77722
rect 29564 77722 29592 78406
rect 30288 78260 30340 78266
rect 30288 78202 30340 78208
rect 28170 77687 28172 77696
rect 27620 77658 27672 77664
rect 28224 77687 28226 77696
rect 29552 77716 29604 77722
rect 28172 77658 28224 77664
rect 29552 77658 29604 77664
rect 27252 77172 27304 77178
rect 27252 77114 27304 77120
rect 27540 77110 27568 77658
rect 27436 77104 27488 77110
rect 27436 77046 27488 77052
rect 27528 77104 27580 77110
rect 27528 77046 27580 77052
rect 26792 77036 26844 77042
rect 26792 76978 26844 76984
rect 26804 76838 26832 76978
rect 26792 76832 26844 76838
rect 26792 76774 26844 76780
rect 26804 76634 26832 76774
rect 27448 76634 27476 77046
rect 26792 76628 26844 76634
rect 26792 76570 26844 76576
rect 27436 76628 27488 76634
rect 27436 76570 27488 76576
rect 24768 76560 24820 76566
rect 24768 76502 24820 76508
rect 24308 76016 24360 76022
rect 24308 75958 24360 75964
rect 22836 74248 22888 74254
rect 22836 74190 22888 74196
rect 21364 73772 21416 73778
rect 21364 73714 21416 73720
rect 26804 72758 26832 76570
rect 26792 72752 26844 72758
rect 26792 72694 26844 72700
rect 7288 72684 7340 72690
rect 7288 72626 7340 72632
rect 7300 60722 7328 72626
rect 28184 72486 28212 77658
rect 30300 76362 30328 78202
rect 30484 77722 30512 79455
rect 31484 78124 31536 78130
rect 31484 78066 31536 78072
rect 30748 78056 30800 78062
rect 30748 77998 30800 78004
rect 30564 77988 30616 77994
rect 30564 77930 30616 77936
rect 30576 77722 30604 77930
rect 30472 77716 30524 77722
rect 30472 77658 30524 77664
rect 30564 77716 30616 77722
rect 30564 77658 30616 77664
rect 30760 77058 30788 77998
rect 31496 77926 31524 78066
rect 31484 77920 31536 77926
rect 31206 77888 31262 77897
rect 31484 77862 31536 77868
rect 31206 77823 31262 77832
rect 31220 77586 31248 77823
rect 31208 77580 31260 77586
rect 31208 77522 31260 77528
rect 31588 77382 31616 79455
rect 31668 77920 31720 77926
rect 31668 77862 31720 77868
rect 31680 77722 31708 77862
rect 32324 77722 32352 79630
rect 34716 79529 34744 79698
rect 33966 79520 34022 79529
rect 33966 79455 34022 79464
rect 34702 79520 34758 79529
rect 34702 79455 34758 79464
rect 32954 78568 33010 78577
rect 32954 78503 33010 78512
rect 32968 77722 32996 78503
rect 33980 78130 34008 79455
rect 33968 78124 34020 78130
rect 33968 78066 34020 78072
rect 33980 77722 34008 78066
rect 34716 77722 34744 79455
rect 35346 78296 35402 78305
rect 35346 78231 35402 78240
rect 34796 78192 34848 78198
rect 34796 78134 34848 78140
rect 34808 77722 34836 78134
rect 34934 77820 35242 77829
rect 34934 77818 34940 77820
rect 34996 77818 35020 77820
rect 35076 77818 35100 77820
rect 35156 77818 35180 77820
rect 35236 77818 35242 77820
rect 34996 77766 34998 77818
rect 35178 77766 35180 77818
rect 34934 77764 34940 77766
rect 34996 77764 35020 77766
rect 35076 77764 35100 77766
rect 35156 77764 35180 77766
rect 35236 77764 35242 77766
rect 34934 77755 35242 77764
rect 31668 77716 31720 77722
rect 31668 77658 31720 77664
rect 32312 77716 32364 77722
rect 32312 77658 32364 77664
rect 32956 77716 33008 77722
rect 32956 77658 33008 77664
rect 33968 77716 34020 77722
rect 33968 77658 34020 77664
rect 34704 77716 34756 77722
rect 34704 77658 34756 77664
rect 34796 77716 34848 77722
rect 34796 77658 34848 77664
rect 35256 77716 35308 77722
rect 35256 77658 35308 77664
rect 32968 77586 32996 77658
rect 32956 77580 33008 77586
rect 32956 77522 33008 77528
rect 35268 77518 35296 77658
rect 35360 77518 35388 78231
rect 36084 77920 36136 77926
rect 36084 77862 36136 77868
rect 35256 77512 35308 77518
rect 35256 77454 35308 77460
rect 35348 77512 35400 77518
rect 35348 77454 35400 77460
rect 31576 77376 31628 77382
rect 31576 77318 31628 77324
rect 32680 77376 32732 77382
rect 35992 77376 36044 77382
rect 32680 77318 32732 77324
rect 35990 77344 35992 77353
rect 36044 77344 36046 77353
rect 30484 77030 30788 77058
rect 30484 76974 30512 77030
rect 30472 76968 30524 76974
rect 30472 76910 30524 76916
rect 30564 76832 30616 76838
rect 30564 76774 30616 76780
rect 30576 76430 30604 76774
rect 32692 76498 32720 77318
rect 35594 77276 35902 77285
rect 35990 77279 36046 77288
rect 35594 77274 35600 77276
rect 35656 77274 35680 77276
rect 35736 77274 35760 77276
rect 35816 77274 35840 77276
rect 35896 77274 35902 77276
rect 35656 77222 35658 77274
rect 35838 77222 35840 77274
rect 35594 77220 35600 77222
rect 35656 77220 35680 77222
rect 35736 77220 35760 77222
rect 35816 77220 35840 77222
rect 35896 77220 35902 77222
rect 35594 77211 35902 77220
rect 34934 76732 35242 76741
rect 34934 76730 34940 76732
rect 34996 76730 35020 76732
rect 35076 76730 35100 76732
rect 35156 76730 35180 76732
rect 35236 76730 35242 76732
rect 34996 76678 34998 76730
rect 35178 76678 35180 76730
rect 34934 76676 34940 76678
rect 34996 76676 35020 76678
rect 35076 76676 35100 76678
rect 35156 76676 35180 76678
rect 35236 76676 35242 76678
rect 34934 76667 35242 76676
rect 32680 76492 32732 76498
rect 32680 76434 32732 76440
rect 30564 76424 30616 76430
rect 30564 76366 30616 76372
rect 30288 76356 30340 76362
rect 30288 76298 30340 76304
rect 35594 76188 35902 76197
rect 35594 76186 35600 76188
rect 35656 76186 35680 76188
rect 35736 76186 35760 76188
rect 35816 76186 35840 76188
rect 35896 76186 35902 76188
rect 35656 76134 35658 76186
rect 35838 76134 35840 76186
rect 35594 76132 35600 76134
rect 35656 76132 35680 76134
rect 35736 76132 35760 76134
rect 35816 76132 35840 76134
rect 35896 76132 35902 76134
rect 35594 76123 35902 76132
rect 34934 75644 35242 75653
rect 34934 75642 34940 75644
rect 34996 75642 35020 75644
rect 35076 75642 35100 75644
rect 35156 75642 35180 75644
rect 35236 75642 35242 75644
rect 34996 75590 34998 75642
rect 35178 75590 35180 75642
rect 34934 75588 34940 75590
rect 34996 75588 35020 75590
rect 35076 75588 35100 75590
rect 35156 75588 35180 75590
rect 35236 75588 35242 75590
rect 34934 75579 35242 75588
rect 35594 75100 35902 75109
rect 35594 75098 35600 75100
rect 35656 75098 35680 75100
rect 35736 75098 35760 75100
rect 35816 75098 35840 75100
rect 35896 75098 35902 75100
rect 35656 75046 35658 75098
rect 35838 75046 35840 75098
rect 35594 75044 35600 75046
rect 35656 75044 35680 75046
rect 35736 75044 35760 75046
rect 35816 75044 35840 75046
rect 35896 75044 35902 75046
rect 35594 75035 35902 75044
rect 34934 74556 35242 74565
rect 34934 74554 34940 74556
rect 34996 74554 35020 74556
rect 35076 74554 35100 74556
rect 35156 74554 35180 74556
rect 35236 74554 35242 74556
rect 34996 74502 34998 74554
rect 35178 74502 35180 74554
rect 34934 74500 34940 74502
rect 34996 74500 35020 74502
rect 35076 74500 35100 74502
rect 35156 74500 35180 74502
rect 35236 74500 35242 74502
rect 34934 74491 35242 74500
rect 35594 74012 35902 74021
rect 35594 74010 35600 74012
rect 35656 74010 35680 74012
rect 35736 74010 35760 74012
rect 35816 74010 35840 74012
rect 35896 74010 35902 74012
rect 35656 73958 35658 74010
rect 35838 73958 35840 74010
rect 35594 73956 35600 73958
rect 35656 73956 35680 73958
rect 35736 73956 35760 73958
rect 35816 73956 35840 73958
rect 35896 73956 35902 73958
rect 35594 73947 35902 73956
rect 34934 73468 35242 73477
rect 34934 73466 34940 73468
rect 34996 73466 35020 73468
rect 35076 73466 35100 73468
rect 35156 73466 35180 73468
rect 35236 73466 35242 73468
rect 34996 73414 34998 73466
rect 35178 73414 35180 73466
rect 34934 73412 34940 73414
rect 34996 73412 35020 73414
rect 35076 73412 35100 73414
rect 35156 73412 35180 73414
rect 35236 73412 35242 73414
rect 34934 73403 35242 73412
rect 35594 72924 35902 72933
rect 35594 72922 35600 72924
rect 35656 72922 35680 72924
rect 35736 72922 35760 72924
rect 35816 72922 35840 72924
rect 35896 72922 35902 72924
rect 35656 72870 35658 72922
rect 35838 72870 35840 72922
rect 35594 72868 35600 72870
rect 35656 72868 35680 72870
rect 35736 72868 35760 72870
rect 35816 72868 35840 72870
rect 35896 72868 35902 72870
rect 35594 72859 35902 72868
rect 28172 72480 28224 72486
rect 28172 72422 28224 72428
rect 34934 72380 35242 72389
rect 34934 72378 34940 72380
rect 34996 72378 35020 72380
rect 35076 72378 35100 72380
rect 35156 72378 35180 72380
rect 35236 72378 35242 72380
rect 34996 72326 34998 72378
rect 35178 72326 35180 72378
rect 34934 72324 34940 72326
rect 34996 72324 35020 72326
rect 35076 72324 35100 72326
rect 35156 72324 35180 72326
rect 35236 72324 35242 72326
rect 34934 72315 35242 72324
rect 9588 72004 9640 72010
rect 9588 71946 9640 71952
rect 7288 60716 7340 60722
rect 7288 60658 7340 60664
rect 6828 60648 6880 60654
rect 6828 60590 6880 60596
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 6840 60314 6868 60590
rect 6828 60308 6880 60314
rect 6828 60250 6880 60256
rect 4874 59868 5182 59877
rect 4874 59866 4880 59868
rect 4936 59866 4960 59868
rect 5016 59866 5040 59868
rect 5096 59866 5120 59868
rect 5176 59866 5182 59868
rect 4936 59814 4938 59866
rect 5118 59814 5120 59866
rect 4874 59812 4880 59814
rect 4936 59812 4960 59814
rect 5016 59812 5040 59814
rect 5096 59812 5120 59814
rect 5176 59812 5182 59814
rect 4874 59803 5182 59812
rect 6840 59770 6868 60250
rect 7300 60110 7328 60658
rect 7288 60104 7340 60110
rect 7288 60046 7340 60052
rect 6828 59764 6880 59770
rect 6828 59706 6880 59712
rect 6840 59650 6868 59706
rect 6840 59622 6960 59650
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 4874 58780 5182 58789
rect 4874 58778 4880 58780
rect 4936 58778 4960 58780
rect 5016 58778 5040 58780
rect 5096 58778 5120 58780
rect 5176 58778 5182 58780
rect 4936 58726 4938 58778
rect 5118 58726 5120 58778
rect 4874 58724 4880 58726
rect 4936 58724 4960 58726
rect 5016 58724 5040 58726
rect 5096 58724 5120 58726
rect 5176 58724 5182 58726
rect 4874 58715 5182 58724
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 4874 57692 5182 57701
rect 4874 57690 4880 57692
rect 4936 57690 4960 57692
rect 5016 57690 5040 57692
rect 5096 57690 5120 57692
rect 5176 57690 5182 57692
rect 4936 57638 4938 57690
rect 5118 57638 5120 57690
rect 4874 57636 4880 57638
rect 4936 57636 4960 57638
rect 5016 57636 5040 57638
rect 5096 57636 5120 57638
rect 5176 57636 5182 57638
rect 4874 57627 5182 57636
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4874 56604 5182 56613
rect 4874 56602 4880 56604
rect 4936 56602 4960 56604
rect 5016 56602 5040 56604
rect 5096 56602 5120 56604
rect 5176 56602 5182 56604
rect 4936 56550 4938 56602
rect 5118 56550 5120 56602
rect 4874 56548 4880 56550
rect 4936 56548 4960 56550
rect 5016 56548 5040 56550
rect 5096 56548 5120 56550
rect 5176 56548 5182 56550
rect 4874 56539 5182 56548
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4874 55516 5182 55525
rect 4874 55514 4880 55516
rect 4936 55514 4960 55516
rect 5016 55514 5040 55516
rect 5096 55514 5120 55516
rect 5176 55514 5182 55516
rect 4936 55462 4938 55514
rect 5118 55462 5120 55514
rect 4874 55460 4880 55462
rect 4936 55460 4960 55462
rect 5016 55460 5040 55462
rect 5096 55460 5120 55462
rect 5176 55460 5182 55462
rect 4874 55451 5182 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4874 54428 5182 54437
rect 4874 54426 4880 54428
rect 4936 54426 4960 54428
rect 5016 54426 5040 54428
rect 5096 54426 5120 54428
rect 5176 54426 5182 54428
rect 4936 54374 4938 54426
rect 5118 54374 5120 54426
rect 4874 54372 4880 54374
rect 4936 54372 4960 54374
rect 5016 54372 5040 54374
rect 5096 54372 5120 54374
rect 5176 54372 5182 54374
rect 4874 54363 5182 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4874 53340 5182 53349
rect 4874 53338 4880 53340
rect 4936 53338 4960 53340
rect 5016 53338 5040 53340
rect 5096 53338 5120 53340
rect 5176 53338 5182 53340
rect 4936 53286 4938 53338
rect 5118 53286 5120 53338
rect 4874 53284 4880 53286
rect 4936 53284 4960 53286
rect 5016 53284 5040 53286
rect 5096 53284 5120 53286
rect 5176 53284 5182 53286
rect 4874 53275 5182 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4874 52252 5182 52261
rect 4874 52250 4880 52252
rect 4936 52250 4960 52252
rect 5016 52250 5040 52252
rect 5096 52250 5120 52252
rect 5176 52250 5182 52252
rect 4936 52198 4938 52250
rect 5118 52198 5120 52250
rect 4874 52196 4880 52198
rect 4936 52196 4960 52198
rect 5016 52196 5040 52198
rect 5096 52196 5120 52198
rect 5176 52196 5182 52198
rect 4874 52187 5182 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4874 51164 5182 51173
rect 4874 51162 4880 51164
rect 4936 51162 4960 51164
rect 5016 51162 5040 51164
rect 5096 51162 5120 51164
rect 5176 51162 5182 51164
rect 4936 51110 4938 51162
rect 5118 51110 5120 51162
rect 4874 51108 4880 51110
rect 4936 51108 4960 51110
rect 5016 51108 5040 51110
rect 5096 51108 5120 51110
rect 5176 51108 5182 51110
rect 4874 51099 5182 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4874 50076 5182 50085
rect 4874 50074 4880 50076
rect 4936 50074 4960 50076
rect 5016 50074 5040 50076
rect 5096 50074 5120 50076
rect 5176 50074 5182 50076
rect 4936 50022 4938 50074
rect 5118 50022 5120 50074
rect 4874 50020 4880 50022
rect 4936 50020 4960 50022
rect 5016 50020 5040 50022
rect 5096 50020 5120 50022
rect 5176 50020 5182 50022
rect 4874 50011 5182 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4874 48988 5182 48997
rect 4874 48986 4880 48988
rect 4936 48986 4960 48988
rect 5016 48986 5040 48988
rect 5096 48986 5120 48988
rect 5176 48986 5182 48988
rect 4936 48934 4938 48986
rect 5118 48934 5120 48986
rect 4874 48932 4880 48934
rect 4936 48932 4960 48934
rect 5016 48932 5040 48934
rect 5096 48932 5120 48934
rect 5176 48932 5182 48934
rect 4874 48923 5182 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4874 47900 5182 47909
rect 4874 47898 4880 47900
rect 4936 47898 4960 47900
rect 5016 47898 5040 47900
rect 5096 47898 5120 47900
rect 5176 47898 5182 47900
rect 4936 47846 4938 47898
rect 5118 47846 5120 47898
rect 4874 47844 4880 47846
rect 4936 47844 4960 47846
rect 5016 47844 5040 47846
rect 5096 47844 5120 47846
rect 5176 47844 5182 47846
rect 4874 47835 5182 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 3424 40044 3476 40050
rect 3424 39986 3476 39992
rect 1768 33108 1820 33114
rect 1768 33050 1820 33056
rect 1584 30320 1636 30326
rect 1584 30262 1636 30268
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1504 13705 1532 13874
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 1308 13252 1360 13258
rect 1308 13194 1360 13200
rect 1320 13025 1348 13194
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 1492 12844 1544 12850
rect 1492 12786 1544 12792
rect 1504 12345 1532 12786
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 1596 11898 1624 30262
rect 1676 26308 1728 26314
rect 1676 26250 1728 26256
rect 1688 12918 1716 26250
rect 1676 12912 1728 12918
rect 1676 12854 1728 12860
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1216 11756 1268 11762
rect 1216 11698 1268 11704
rect 1228 11665 1256 11698
rect 1214 11656 1270 11665
rect 1214 11591 1270 11600
rect 1492 11076 1544 11082
rect 1492 11018 1544 11024
rect 1504 10985 1532 11018
rect 1490 10976 1546 10985
rect 1490 10911 1546 10920
rect 1780 10810 1808 33050
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 1872 13530 1900 23598
rect 3436 14074 3464 39986
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10305 1348 10610
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 1306 10296 1362 10305
rect 4214 10299 4522 10308
rect 1306 10231 1362 10240
rect 1492 9988 1544 9994
rect 1492 9930 1544 9936
rect 1504 9625 1532 9930
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 1490 9616 1546 9625
rect 6932 9586 6960 59622
rect 7564 41472 7616 41478
rect 7564 41414 7616 41420
rect 7576 41313 7604 41414
rect 7562 41304 7618 41313
rect 7562 41239 7618 41248
rect 7576 40050 7604 41239
rect 7564 40044 7616 40050
rect 7564 39986 7616 39992
rect 7288 39840 7340 39846
rect 7288 39782 7340 39788
rect 7300 39545 7328 39782
rect 7286 39536 7342 39545
rect 7286 39471 7342 39480
rect 7300 11354 7328 39471
rect 7564 38752 7616 38758
rect 7564 38694 7616 38700
rect 7576 38457 7604 38694
rect 7562 38448 7618 38457
rect 7618 38406 7696 38434
rect 7562 38383 7618 38392
rect 7562 36680 7618 36689
rect 7562 36615 7564 36624
rect 7616 36615 7618 36624
rect 7564 36586 7616 36592
rect 7576 36394 7604 36586
rect 7392 36366 7604 36394
rect 7392 26314 7420 36366
rect 7470 35592 7526 35601
rect 7470 35527 7526 35536
rect 7484 35494 7512 35527
rect 7472 35488 7524 35494
rect 7472 35430 7524 35436
rect 7484 30326 7512 35430
rect 7562 33960 7618 33969
rect 7562 33895 7564 33904
rect 7616 33895 7618 33904
rect 7564 33866 7616 33872
rect 7576 33114 7604 33866
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7472 30320 7524 30326
rect 7472 30262 7524 30268
rect 7380 26308 7432 26314
rect 7380 26250 7432 26256
rect 7668 26234 7696 38406
rect 7576 26206 7696 26234
rect 7576 23662 7604 26206
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7470 15464 7526 15473
rect 7470 15399 7526 15408
rect 7484 15366 7512 15399
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 1490 9551 1546 9560
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 1306 8936 1362 8945
rect 1306 8871 1308 8880
rect 1360 8871 1362 8880
rect 1308 8842 1360 8848
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1950 8256 2006 8265
rect 2056 8242 2084 8366
rect 2006 8214 2084 8242
rect 1950 8191 2006 8200
rect 1964 8090 1992 8191
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1308 7812 1360 7818
rect 1308 7754 1360 7760
rect 1320 7585 1348 7754
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 1306 7576 1362 7585
rect 4874 7579 5182 7588
rect 1306 7511 1362 7520
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1320 6905 1348 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 1306 6896 1362 6905
rect 1306 6831 1362 6840
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 1216 6316 1268 6322
rect 1216 6258 1268 6264
rect 1228 6225 1256 6258
rect 1214 6216 1270 6225
rect 1214 6151 1270 6160
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 7484 5914 7512 15302
rect 9600 9654 9628 71946
rect 35594 71836 35902 71845
rect 35594 71834 35600 71836
rect 35656 71834 35680 71836
rect 35736 71834 35760 71836
rect 35816 71834 35840 71836
rect 35896 71834 35902 71836
rect 35656 71782 35658 71834
rect 35838 71782 35840 71834
rect 35594 71780 35600 71782
rect 35656 71780 35680 71782
rect 35736 71780 35760 71782
rect 35816 71780 35840 71782
rect 35896 71780 35902 71782
rect 35594 71771 35902 71780
rect 34934 71292 35242 71301
rect 34934 71290 34940 71292
rect 34996 71290 35020 71292
rect 35076 71290 35100 71292
rect 35156 71290 35180 71292
rect 35236 71290 35242 71292
rect 34996 71238 34998 71290
rect 35178 71238 35180 71290
rect 34934 71236 34940 71238
rect 34996 71236 35020 71238
rect 35076 71236 35100 71238
rect 35156 71236 35180 71238
rect 35236 71236 35242 71238
rect 34934 71227 35242 71236
rect 35594 70748 35902 70757
rect 35594 70746 35600 70748
rect 35656 70746 35680 70748
rect 35736 70746 35760 70748
rect 35816 70746 35840 70748
rect 35896 70746 35902 70748
rect 35656 70694 35658 70746
rect 35838 70694 35840 70746
rect 35594 70692 35600 70694
rect 35656 70692 35680 70694
rect 35736 70692 35760 70694
rect 35816 70692 35840 70694
rect 35896 70692 35902 70694
rect 35594 70683 35902 70692
rect 34934 70204 35242 70213
rect 34934 70202 34940 70204
rect 34996 70202 35020 70204
rect 35076 70202 35100 70204
rect 35156 70202 35180 70204
rect 35236 70202 35242 70204
rect 34996 70150 34998 70202
rect 35178 70150 35180 70202
rect 34934 70148 34940 70150
rect 34996 70148 35020 70150
rect 35076 70148 35100 70150
rect 35156 70148 35180 70150
rect 35236 70148 35242 70150
rect 34934 70139 35242 70148
rect 35594 69660 35902 69669
rect 35594 69658 35600 69660
rect 35656 69658 35680 69660
rect 35736 69658 35760 69660
rect 35816 69658 35840 69660
rect 35896 69658 35902 69660
rect 35656 69606 35658 69658
rect 35838 69606 35840 69658
rect 35594 69604 35600 69606
rect 35656 69604 35680 69606
rect 35736 69604 35760 69606
rect 35816 69604 35840 69606
rect 35896 69604 35902 69606
rect 35594 69595 35902 69604
rect 34934 69116 35242 69125
rect 34934 69114 34940 69116
rect 34996 69114 35020 69116
rect 35076 69114 35100 69116
rect 35156 69114 35180 69116
rect 35236 69114 35242 69116
rect 34996 69062 34998 69114
rect 35178 69062 35180 69114
rect 34934 69060 34940 69062
rect 34996 69060 35020 69062
rect 35076 69060 35100 69062
rect 35156 69060 35180 69062
rect 35236 69060 35242 69062
rect 34934 69051 35242 69060
rect 35594 68572 35902 68581
rect 35594 68570 35600 68572
rect 35656 68570 35680 68572
rect 35736 68570 35760 68572
rect 35816 68570 35840 68572
rect 35896 68570 35902 68572
rect 35656 68518 35658 68570
rect 35838 68518 35840 68570
rect 35594 68516 35600 68518
rect 35656 68516 35680 68518
rect 35736 68516 35760 68518
rect 35816 68516 35840 68518
rect 35896 68516 35902 68518
rect 35594 68507 35902 68516
rect 34934 68028 35242 68037
rect 34934 68026 34940 68028
rect 34996 68026 35020 68028
rect 35076 68026 35100 68028
rect 35156 68026 35180 68028
rect 35236 68026 35242 68028
rect 34996 67974 34998 68026
rect 35178 67974 35180 68026
rect 34934 67972 34940 67974
rect 34996 67972 35020 67974
rect 35076 67972 35100 67974
rect 35156 67972 35180 67974
rect 35236 67972 35242 67974
rect 34934 67963 35242 67972
rect 35594 67484 35902 67493
rect 35594 67482 35600 67484
rect 35656 67482 35680 67484
rect 35736 67482 35760 67484
rect 35816 67482 35840 67484
rect 35896 67482 35902 67484
rect 35656 67430 35658 67482
rect 35838 67430 35840 67482
rect 35594 67428 35600 67430
rect 35656 67428 35680 67430
rect 35736 67428 35760 67430
rect 35816 67428 35840 67430
rect 35896 67428 35902 67430
rect 35594 67419 35902 67428
rect 34934 66940 35242 66949
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66875 35242 66884
rect 35594 66396 35902 66405
rect 35594 66394 35600 66396
rect 35656 66394 35680 66396
rect 35736 66394 35760 66396
rect 35816 66394 35840 66396
rect 35896 66394 35902 66396
rect 35656 66342 35658 66394
rect 35838 66342 35840 66394
rect 35594 66340 35600 66342
rect 35656 66340 35680 66342
rect 35736 66340 35760 66342
rect 35816 66340 35840 66342
rect 35896 66340 35902 66342
rect 35594 66331 35902 66340
rect 36096 66230 36124 77862
rect 36280 77518 36308 79766
rect 37002 79656 37058 79665
rect 37002 79591 37058 79600
rect 37016 79558 37044 79591
rect 37004 79552 37056 79558
rect 37004 79494 37056 79500
rect 37016 77518 37044 79494
rect 37738 78160 37794 78169
rect 37738 78095 37794 78104
rect 36268 77512 36320 77518
rect 36268 77454 36320 77460
rect 37004 77512 37056 77518
rect 37004 77454 37056 77460
rect 37752 77382 37780 78095
rect 38672 77654 38700 79834
rect 39776 77654 39804 79863
rect 39856 78056 39908 78062
rect 39856 77998 39908 78004
rect 40130 78024 40186 78033
rect 39868 77654 39896 77998
rect 40130 77959 40186 77968
rect 40866 78024 40922 78033
rect 40866 77959 40922 77968
rect 38660 77648 38712 77654
rect 38660 77590 38712 77596
rect 39764 77648 39816 77654
rect 39764 77590 39816 77596
rect 39856 77648 39908 77654
rect 39856 77590 39908 77596
rect 40040 77512 40092 77518
rect 40038 77480 40040 77489
rect 40092 77480 40094 77489
rect 39948 77444 40000 77450
rect 40038 77415 40094 77424
rect 39948 77386 40000 77392
rect 37280 77376 37332 77382
rect 37280 77318 37332 77324
rect 37740 77376 37792 77382
rect 39960 77353 39988 77386
rect 40144 77382 40172 77959
rect 40684 77716 40736 77722
rect 40684 77658 40736 77664
rect 40132 77376 40184 77382
rect 37740 77318 37792 77324
rect 37922 77344 37978 77353
rect 37292 76022 37320 77318
rect 37922 77279 37978 77288
rect 39946 77344 40002 77353
rect 40132 77318 40184 77324
rect 39946 77279 40002 77288
rect 37280 76016 37332 76022
rect 37280 75958 37332 75964
rect 37936 66230 37964 77279
rect 40696 70394 40724 77658
rect 40880 77654 40908 77959
rect 40972 77654 41000 79863
rect 42154 79520 42210 79529
rect 42154 79455 42210 79464
rect 43258 79520 43314 79529
rect 43258 79455 43314 79464
rect 42168 79014 42196 79455
rect 42156 79008 42208 79014
rect 42156 78950 42208 78956
rect 42168 77654 42196 78950
rect 43272 77994 43300 79455
rect 61108 79348 61160 79354
rect 61108 79290 61160 79296
rect 58624 78056 58676 78062
rect 58624 77998 58676 78004
rect 43260 77988 43312 77994
rect 43260 77930 43312 77936
rect 43812 77988 43864 77994
rect 43812 77930 43864 77936
rect 53564 77988 53616 77994
rect 53564 77930 53616 77936
rect 40868 77648 40920 77654
rect 40868 77590 40920 77596
rect 40960 77648 41012 77654
rect 40960 77590 41012 77596
rect 42156 77648 42208 77654
rect 42156 77590 42208 77596
rect 42890 77616 42946 77625
rect 43824 77586 43852 77930
rect 42890 77551 42946 77560
rect 43812 77580 43864 77586
rect 42904 77382 42932 77551
rect 43812 77522 43864 77528
rect 46112 77512 46164 77518
rect 43626 77480 43682 77489
rect 46112 77454 46164 77460
rect 43626 77415 43682 77424
rect 42432 77376 42484 77382
rect 42430 77344 42432 77353
rect 42892 77376 42944 77382
rect 42484 77344 42486 77353
rect 42892 77318 42944 77324
rect 42430 77279 42486 77288
rect 40696 70366 41184 70394
rect 41156 66230 41184 70366
rect 43640 66230 43668 77415
rect 44180 72684 44232 72690
rect 44180 72626 44232 72632
rect 44192 72282 44220 72626
rect 44180 72276 44232 72282
rect 44180 72218 44232 72224
rect 46124 66230 46152 77454
rect 48596 77444 48648 77450
rect 48596 77386 48648 77392
rect 51080 77444 51132 77450
rect 51080 77386 51132 77392
rect 48608 66230 48636 77386
rect 51092 66230 51120 77386
rect 53576 66230 53604 77930
rect 56140 77920 56192 77926
rect 56140 77862 56192 77868
rect 56152 66230 56180 77862
rect 57796 72548 57848 72554
rect 57796 72490 57848 72496
rect 57808 72010 57836 72490
rect 57796 72004 57848 72010
rect 57796 71946 57848 71952
rect 58636 66230 58664 77998
rect 61120 77518 61148 79290
rect 88892 79008 88944 79014
rect 88892 78950 88944 78956
rect 63314 78568 63370 78577
rect 63314 78503 63370 78512
rect 79232 78532 79284 78538
rect 62488 77988 62540 77994
rect 62488 77930 62540 77936
rect 62500 77654 62528 77930
rect 62488 77648 62540 77654
rect 62488 77590 62540 77596
rect 61108 77512 61160 77518
rect 61108 77454 61160 77460
rect 62500 77450 62528 77590
rect 63328 77518 63356 78503
rect 79232 78474 79284 78480
rect 76656 78464 76708 78470
rect 76656 78406 76708 78412
rect 78770 78432 78826 78441
rect 71964 78396 72016 78402
rect 71964 78338 72016 78344
rect 69756 78260 69808 78266
rect 69756 78202 69808 78208
rect 63960 78192 64012 78198
rect 63960 78134 64012 78140
rect 63592 78124 63644 78130
rect 63592 78066 63644 78072
rect 63316 77512 63368 77518
rect 63316 77454 63368 77460
rect 62488 77444 62540 77450
rect 62488 77386 62540 77392
rect 61108 76832 61160 76838
rect 61108 76774 61160 76780
rect 61120 66230 61148 76774
rect 63604 66230 63632 78066
rect 63972 77654 64000 78134
rect 69112 78056 69164 78062
rect 69112 77998 69164 78004
rect 66076 77988 66128 77994
rect 66076 77930 66128 77936
rect 64144 77920 64196 77926
rect 64144 77862 64196 77868
rect 63960 77648 64012 77654
rect 63960 77590 64012 77596
rect 64156 77586 64184 77862
rect 65654 77820 65962 77829
rect 65654 77818 65660 77820
rect 65716 77818 65740 77820
rect 65796 77818 65820 77820
rect 65876 77818 65900 77820
rect 65956 77818 65962 77820
rect 65716 77766 65718 77818
rect 65898 77766 65900 77818
rect 65654 77764 65660 77766
rect 65716 77764 65740 77766
rect 65796 77764 65820 77766
rect 65876 77764 65900 77766
rect 65956 77764 65962 77766
rect 65654 77755 65962 77764
rect 64972 77648 65024 77654
rect 64972 77590 65024 77596
rect 64052 77580 64104 77586
rect 64052 77522 64104 77528
rect 64144 77580 64196 77586
rect 64144 77522 64196 77528
rect 64064 77382 64092 77522
rect 64984 77382 65012 77590
rect 65892 77512 65944 77518
rect 65890 77480 65892 77489
rect 65944 77480 65946 77489
rect 65890 77415 65946 77424
rect 64052 77376 64104 77382
rect 64052 77318 64104 77324
rect 64972 77376 65024 77382
rect 64972 77318 65024 77324
rect 65654 76732 65962 76741
rect 65654 76730 65660 76732
rect 65716 76730 65740 76732
rect 65796 76730 65820 76732
rect 65876 76730 65900 76732
rect 65956 76730 65962 76732
rect 65716 76678 65718 76730
rect 65898 76678 65900 76730
rect 65654 76676 65660 76678
rect 65716 76676 65740 76678
rect 65796 76676 65820 76678
rect 65876 76676 65900 76678
rect 65956 76676 65962 76678
rect 65654 76667 65962 76676
rect 65654 75644 65962 75653
rect 65654 75642 65660 75644
rect 65716 75642 65740 75644
rect 65796 75642 65820 75644
rect 65876 75642 65900 75644
rect 65956 75642 65962 75644
rect 65716 75590 65718 75642
rect 65898 75590 65900 75642
rect 65654 75588 65660 75590
rect 65716 75588 65740 75590
rect 65796 75588 65820 75590
rect 65876 75588 65900 75590
rect 65956 75588 65962 75590
rect 65654 75579 65962 75588
rect 65654 74556 65962 74565
rect 65654 74554 65660 74556
rect 65716 74554 65740 74556
rect 65796 74554 65820 74556
rect 65876 74554 65900 74556
rect 65956 74554 65962 74556
rect 65716 74502 65718 74554
rect 65898 74502 65900 74554
rect 65654 74500 65660 74502
rect 65716 74500 65740 74502
rect 65796 74500 65820 74502
rect 65876 74500 65900 74502
rect 65956 74500 65962 74502
rect 65654 74491 65962 74500
rect 65654 73468 65962 73477
rect 65654 73466 65660 73468
rect 65716 73466 65740 73468
rect 65796 73466 65820 73468
rect 65876 73466 65900 73468
rect 65956 73466 65962 73468
rect 65716 73414 65718 73466
rect 65898 73414 65900 73466
rect 65654 73412 65660 73414
rect 65716 73412 65740 73414
rect 65796 73412 65820 73414
rect 65876 73412 65900 73414
rect 65956 73412 65962 73414
rect 65654 73403 65962 73412
rect 65654 72380 65962 72389
rect 65654 72378 65660 72380
rect 65716 72378 65740 72380
rect 65796 72378 65820 72380
rect 65876 72378 65900 72380
rect 65956 72378 65962 72380
rect 65716 72326 65718 72378
rect 65898 72326 65900 72378
rect 65654 72324 65660 72326
rect 65716 72324 65740 72326
rect 65796 72324 65820 72326
rect 65876 72324 65900 72326
rect 65956 72324 65962 72326
rect 65654 72315 65962 72324
rect 65654 71292 65962 71301
rect 65654 71290 65660 71292
rect 65716 71290 65740 71292
rect 65796 71290 65820 71292
rect 65876 71290 65900 71292
rect 65956 71290 65962 71292
rect 65716 71238 65718 71290
rect 65898 71238 65900 71290
rect 65654 71236 65660 71238
rect 65716 71236 65740 71238
rect 65796 71236 65820 71238
rect 65876 71236 65900 71238
rect 65956 71236 65962 71238
rect 65654 71227 65962 71236
rect 65654 70204 65962 70213
rect 65654 70202 65660 70204
rect 65716 70202 65740 70204
rect 65796 70202 65820 70204
rect 65876 70202 65900 70204
rect 65956 70202 65962 70204
rect 65716 70150 65718 70202
rect 65898 70150 65900 70202
rect 65654 70148 65660 70150
rect 65716 70148 65740 70150
rect 65796 70148 65820 70150
rect 65876 70148 65900 70150
rect 65956 70148 65962 70150
rect 65654 70139 65962 70148
rect 65654 69116 65962 69125
rect 65654 69114 65660 69116
rect 65716 69114 65740 69116
rect 65796 69114 65820 69116
rect 65876 69114 65900 69116
rect 65956 69114 65962 69116
rect 65716 69062 65718 69114
rect 65898 69062 65900 69114
rect 65654 69060 65660 69062
rect 65716 69060 65740 69062
rect 65796 69060 65820 69062
rect 65876 69060 65900 69062
rect 65956 69060 65962 69062
rect 65654 69051 65962 69060
rect 65654 68028 65962 68037
rect 65654 68026 65660 68028
rect 65716 68026 65740 68028
rect 65796 68026 65820 68028
rect 65876 68026 65900 68028
rect 65956 68026 65962 68028
rect 65716 67974 65718 68026
rect 65898 67974 65900 68026
rect 65654 67972 65660 67974
rect 65716 67972 65740 67974
rect 65796 67972 65820 67974
rect 65876 67972 65900 67974
rect 65956 67972 65962 67974
rect 65654 67963 65962 67972
rect 65654 66940 65962 66949
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66875 65962 66884
rect 66088 66230 66116 77930
rect 67640 77920 67692 77926
rect 67640 77862 67692 77868
rect 67652 77654 67680 77862
rect 69124 77654 69152 77998
rect 67640 77648 67692 77654
rect 69112 77648 69164 77654
rect 67640 77590 67692 77596
rect 68466 77616 68522 77625
rect 68284 77580 68336 77586
rect 69112 77590 69164 77596
rect 69768 77586 69796 78202
rect 71136 78124 71188 78130
rect 71136 78066 71188 78072
rect 70950 78024 71006 78033
rect 70950 77959 71006 77968
rect 70400 77920 70452 77926
rect 70400 77862 70452 77868
rect 70412 77722 70440 77862
rect 70964 77722 70992 77959
rect 70400 77716 70452 77722
rect 70400 77658 70452 77664
rect 70952 77716 71004 77722
rect 70952 77658 71004 77664
rect 71044 77716 71096 77722
rect 71044 77658 71096 77664
rect 68466 77551 68468 77560
rect 68284 77522 68336 77528
rect 68520 77551 68522 77560
rect 69204 77580 69256 77586
rect 68468 77522 68520 77528
rect 69204 77522 69256 77528
rect 69756 77580 69808 77586
rect 69756 77522 69808 77528
rect 67364 77512 67416 77518
rect 67364 77454 67416 77460
rect 66314 77276 66622 77285
rect 66314 77274 66320 77276
rect 66376 77274 66400 77276
rect 66456 77274 66480 77276
rect 66536 77274 66560 77276
rect 66616 77274 66622 77276
rect 66376 77222 66378 77274
rect 66558 77222 66560 77274
rect 66314 77220 66320 77222
rect 66376 77220 66400 77222
rect 66456 77220 66480 77222
rect 66536 77220 66560 77222
rect 66616 77220 66622 77222
rect 66314 77211 66622 77220
rect 66314 76188 66622 76197
rect 66314 76186 66320 76188
rect 66376 76186 66400 76188
rect 66456 76186 66480 76188
rect 66536 76186 66560 76188
rect 66616 76186 66622 76188
rect 66376 76134 66378 76186
rect 66558 76134 66560 76186
rect 66314 76132 66320 76134
rect 66376 76132 66400 76134
rect 66456 76132 66480 76134
rect 66536 76132 66560 76134
rect 66616 76132 66622 76134
rect 66314 76123 66622 76132
rect 67376 75274 67404 77454
rect 68296 77382 68324 77522
rect 69216 77382 69244 77522
rect 69768 77382 69796 77522
rect 68284 77376 68336 77382
rect 68284 77318 68336 77324
rect 69204 77376 69256 77382
rect 69204 77318 69256 77324
rect 69756 77376 69808 77382
rect 69756 77318 69808 77324
rect 69848 77376 69900 77382
rect 69848 77318 69900 77324
rect 68560 77172 68612 77178
rect 68560 77114 68612 77120
rect 67364 75268 67416 75274
rect 67364 75210 67416 75216
rect 66314 75100 66622 75109
rect 66314 75098 66320 75100
rect 66376 75098 66400 75100
rect 66456 75098 66480 75100
rect 66536 75098 66560 75100
rect 66616 75098 66622 75100
rect 66376 75046 66378 75098
rect 66558 75046 66560 75098
rect 66314 75044 66320 75046
rect 66376 75044 66400 75046
rect 66456 75044 66480 75046
rect 66536 75044 66560 75046
rect 66616 75044 66622 75046
rect 66314 75035 66622 75044
rect 66314 74012 66622 74021
rect 66314 74010 66320 74012
rect 66376 74010 66400 74012
rect 66456 74010 66480 74012
rect 66536 74010 66560 74012
rect 66616 74010 66622 74012
rect 66376 73958 66378 74010
rect 66558 73958 66560 74010
rect 66314 73956 66320 73958
rect 66376 73956 66400 73958
rect 66456 73956 66480 73958
rect 66536 73956 66560 73958
rect 66616 73956 66622 73958
rect 66314 73947 66622 73956
rect 66314 72924 66622 72933
rect 66314 72922 66320 72924
rect 66376 72922 66400 72924
rect 66456 72922 66480 72924
rect 66536 72922 66560 72924
rect 66616 72922 66622 72924
rect 66376 72870 66378 72922
rect 66558 72870 66560 72922
rect 66314 72868 66320 72870
rect 66376 72868 66400 72870
rect 66456 72868 66480 72870
rect 66536 72868 66560 72870
rect 66616 72868 66622 72870
rect 66314 72859 66622 72868
rect 66314 71836 66622 71845
rect 66314 71834 66320 71836
rect 66376 71834 66400 71836
rect 66456 71834 66480 71836
rect 66536 71834 66560 71836
rect 66616 71834 66622 71836
rect 66376 71782 66378 71834
rect 66558 71782 66560 71834
rect 66314 71780 66320 71782
rect 66376 71780 66400 71782
rect 66456 71780 66480 71782
rect 66536 71780 66560 71782
rect 66616 71780 66622 71782
rect 66314 71771 66622 71780
rect 66314 70748 66622 70757
rect 66314 70746 66320 70748
rect 66376 70746 66400 70748
rect 66456 70746 66480 70748
rect 66536 70746 66560 70748
rect 66616 70746 66622 70748
rect 66376 70694 66378 70746
rect 66558 70694 66560 70746
rect 66314 70692 66320 70694
rect 66376 70692 66400 70694
rect 66456 70692 66480 70694
rect 66536 70692 66560 70694
rect 66616 70692 66622 70694
rect 66314 70683 66622 70692
rect 66314 69660 66622 69669
rect 66314 69658 66320 69660
rect 66376 69658 66400 69660
rect 66456 69658 66480 69660
rect 66536 69658 66560 69660
rect 66616 69658 66622 69660
rect 66376 69606 66378 69658
rect 66558 69606 66560 69658
rect 66314 69604 66320 69606
rect 66376 69604 66400 69606
rect 66456 69604 66480 69606
rect 66536 69604 66560 69606
rect 66616 69604 66622 69606
rect 66314 69595 66622 69604
rect 66314 68572 66622 68581
rect 66314 68570 66320 68572
rect 66376 68570 66400 68572
rect 66456 68570 66480 68572
rect 66536 68570 66560 68572
rect 66616 68570 66622 68572
rect 66376 68518 66378 68570
rect 66558 68518 66560 68570
rect 66314 68516 66320 68518
rect 66376 68516 66400 68518
rect 66456 68516 66480 68518
rect 66536 68516 66560 68518
rect 66616 68516 66622 68518
rect 66314 68507 66622 68516
rect 66314 67484 66622 67493
rect 66314 67482 66320 67484
rect 66376 67482 66400 67484
rect 66456 67482 66480 67484
rect 66536 67482 66560 67484
rect 66616 67482 66622 67484
rect 66376 67430 66378 67482
rect 66558 67430 66560 67482
rect 66314 67428 66320 67430
rect 66376 67428 66400 67430
rect 66456 67428 66480 67430
rect 66536 67428 66560 67430
rect 66616 67428 66622 67430
rect 66314 67419 66622 67428
rect 66314 66396 66622 66405
rect 66314 66394 66320 66396
rect 66376 66394 66400 66396
rect 66456 66394 66480 66396
rect 66536 66394 66560 66396
rect 66616 66394 66622 66396
rect 66376 66342 66378 66394
rect 66558 66342 66560 66394
rect 66314 66340 66320 66342
rect 66376 66340 66400 66342
rect 66456 66340 66480 66342
rect 66536 66340 66560 66342
rect 66616 66340 66622 66342
rect 66314 66331 66622 66340
rect 68572 66230 68600 77114
rect 69216 77110 69244 77318
rect 69204 77104 69256 77110
rect 69204 77046 69256 77052
rect 69860 76906 69888 77318
rect 69848 76900 69900 76906
rect 69848 76842 69900 76848
rect 71056 66230 71084 77658
rect 71148 77654 71176 78066
rect 71686 78024 71742 78033
rect 71686 77959 71742 77968
rect 71136 77648 71188 77654
rect 71136 77590 71188 77596
rect 71148 77382 71176 77590
rect 71320 77444 71372 77450
rect 71320 77386 71372 77392
rect 71136 77376 71188 77382
rect 71136 77318 71188 77324
rect 71332 77194 71360 77386
rect 71700 77382 71728 77959
rect 71976 77722 72004 78338
rect 73528 78328 73580 78334
rect 73528 78270 73580 78276
rect 76194 78296 76250 78305
rect 73436 77988 73488 77994
rect 73436 77930 73488 77936
rect 71964 77716 72016 77722
rect 71964 77658 72016 77664
rect 73448 77450 73476 77930
rect 73436 77444 73488 77450
rect 73436 77386 73488 77392
rect 71688 77376 71740 77382
rect 71688 77318 71740 77324
rect 71332 77166 71820 77194
rect 71792 75886 71820 77166
rect 71780 75880 71832 75886
rect 71780 75822 71832 75828
rect 73540 66230 73568 78270
rect 76194 78231 76250 78240
rect 73986 78160 74042 78169
rect 73986 78095 74042 78104
rect 74448 78124 74500 78130
rect 74000 77586 74028 78095
rect 74448 78066 74500 78072
rect 74460 77722 74488 78066
rect 74448 77716 74500 77722
rect 74448 77658 74500 77664
rect 76208 77586 76236 78231
rect 76668 77722 76696 78406
rect 78770 78367 78826 78376
rect 78784 77722 78812 78367
rect 79244 77722 79272 78474
rect 85672 78396 85724 78402
rect 85672 78338 85724 78344
rect 80060 78328 80112 78334
rect 80060 78270 80112 78276
rect 80072 77722 80100 78270
rect 81348 78192 81400 78198
rect 81348 78134 81400 78140
rect 80888 77988 80940 77994
rect 80888 77930 80940 77936
rect 76656 77716 76708 77722
rect 76656 77658 76708 77664
rect 78772 77716 78824 77722
rect 78772 77658 78824 77664
rect 79232 77716 79284 77722
rect 79232 77658 79284 77664
rect 80060 77716 80112 77722
rect 80060 77658 80112 77664
rect 78784 77586 78812 77658
rect 73804 77580 73856 77586
rect 73804 77522 73856 77528
rect 73988 77580 74040 77586
rect 73988 77522 74040 77528
rect 76196 77580 76248 77586
rect 76196 77522 76248 77528
rect 78772 77580 78824 77586
rect 78772 77522 78824 77528
rect 73816 77382 73844 77522
rect 74632 77512 74684 77518
rect 74632 77454 74684 77460
rect 73804 77376 73856 77382
rect 73804 77318 73856 77324
rect 73988 76288 74040 76294
rect 73988 76230 74040 76236
rect 74000 72078 74028 76230
rect 74080 72752 74132 72758
rect 74080 72694 74132 72700
rect 74092 72282 74120 72694
rect 74080 72276 74132 72282
rect 74080 72218 74132 72224
rect 73988 72072 74040 72078
rect 73988 72014 74040 72020
rect 74356 72072 74408 72078
rect 74356 72014 74408 72020
rect 74368 71942 74396 72014
rect 74356 71936 74408 71942
rect 74356 71878 74408 71884
rect 74368 68746 74396 71878
rect 74644 71058 74672 77454
rect 76208 77382 76236 77522
rect 80072 77518 80100 77658
rect 80900 77654 80928 77930
rect 80888 77648 80940 77654
rect 80888 77590 80940 77596
rect 80060 77512 80112 77518
rect 80060 77454 80112 77460
rect 75644 77376 75696 77382
rect 75644 77318 75696 77324
rect 76196 77376 76248 77382
rect 76196 77318 76248 77324
rect 76288 77376 76340 77382
rect 76288 77318 76340 77324
rect 75656 77110 75684 77318
rect 76300 77178 76328 77318
rect 76288 77172 76340 77178
rect 76288 77114 76340 77120
rect 75644 77104 75696 77110
rect 75644 77046 75696 77052
rect 81360 76022 81388 78134
rect 83832 77512 83884 77518
rect 83832 77454 83884 77460
rect 81532 77444 81584 77450
rect 81532 77386 81584 77392
rect 83096 77444 83148 77450
rect 83096 77386 83148 77392
rect 81544 77178 81572 77386
rect 83108 77178 83136 77386
rect 83648 77376 83700 77382
rect 83648 77318 83700 77324
rect 81532 77172 81584 77178
rect 81532 77114 81584 77120
rect 83096 77172 83148 77178
rect 83096 77114 83148 77120
rect 82820 76832 82872 76838
rect 82820 76774 82872 76780
rect 82832 76430 82860 76774
rect 83660 76498 83688 77318
rect 83844 77042 83872 77454
rect 84292 77444 84344 77450
rect 84292 77386 84344 77392
rect 84016 77376 84068 77382
rect 84016 77318 84068 77324
rect 83832 77036 83884 77042
rect 83832 76978 83884 76984
rect 83924 76968 83976 76974
rect 83924 76910 83976 76916
rect 83648 76492 83700 76498
rect 83648 76434 83700 76440
rect 82820 76424 82872 76430
rect 82820 76366 82872 76372
rect 82832 76090 82860 76366
rect 83280 76356 83332 76362
rect 83280 76298 83332 76304
rect 82820 76084 82872 76090
rect 82820 76026 82872 76032
rect 81348 76016 81400 76022
rect 81348 75958 81400 75964
rect 82176 75336 82228 75342
rect 82176 75278 82228 75284
rect 82084 75200 82136 75206
rect 82084 75142 82136 75148
rect 77208 72752 77260 72758
rect 77208 72694 77260 72700
rect 75092 72616 75144 72622
rect 75092 72558 75144 72564
rect 74632 71052 74684 71058
rect 74632 70994 74684 71000
rect 75104 70990 75132 72558
rect 75092 70984 75144 70990
rect 75092 70926 75144 70932
rect 77220 70446 77248 72694
rect 82096 72622 82124 75142
rect 82188 75002 82216 75278
rect 82832 75002 82860 76026
rect 83292 76022 83320 76298
rect 83936 76090 83964 76910
rect 84028 76838 84056 77318
rect 84016 76832 84068 76838
rect 84016 76774 84068 76780
rect 84304 76634 84332 77386
rect 85580 77036 85632 77042
rect 85580 76978 85632 76984
rect 85592 76838 85620 76978
rect 85684 76974 85712 78338
rect 85948 78056 86000 78062
rect 85948 77998 86000 78004
rect 87328 78056 87380 78062
rect 87328 77998 87380 78004
rect 85764 77104 85816 77110
rect 85764 77046 85816 77052
rect 85672 76968 85724 76974
rect 85672 76910 85724 76916
rect 85580 76832 85632 76838
rect 85580 76774 85632 76780
rect 85776 76634 85804 77046
rect 85960 76634 85988 77998
rect 87052 77920 87104 77926
rect 87052 77862 87104 77868
rect 86592 77648 86644 77654
rect 86592 77590 86644 77596
rect 86500 77580 86552 77586
rect 86500 77522 86552 77528
rect 86408 77512 86460 77518
rect 86408 77454 86460 77460
rect 86420 77042 86448 77454
rect 86512 77382 86540 77522
rect 86500 77376 86552 77382
rect 86500 77318 86552 77324
rect 86512 77042 86540 77318
rect 86408 77036 86460 77042
rect 86408 76978 86460 76984
rect 86500 77036 86552 77042
rect 86500 76978 86552 76984
rect 86604 76838 86632 77590
rect 86868 77512 86920 77518
rect 86868 77454 86920 77460
rect 86880 77042 86908 77454
rect 86868 77036 86920 77042
rect 86868 76978 86920 76984
rect 86776 76900 86828 76906
rect 86776 76842 86828 76848
rect 86132 76832 86184 76838
rect 86132 76774 86184 76780
rect 86592 76832 86644 76838
rect 86592 76774 86644 76780
rect 86144 76634 86172 76774
rect 84292 76628 84344 76634
rect 84292 76570 84344 76576
rect 85764 76628 85816 76634
rect 85764 76570 85816 76576
rect 85948 76628 86000 76634
rect 85948 76570 86000 76576
rect 86132 76628 86184 76634
rect 86132 76570 86184 76576
rect 85960 76514 85988 76570
rect 85960 76486 86356 76514
rect 86328 76378 86356 76486
rect 86328 76362 86448 76378
rect 86328 76356 86460 76362
rect 86328 76350 86408 76356
rect 86408 76298 86460 76304
rect 85580 76288 85632 76294
rect 85580 76230 85632 76236
rect 83924 76084 83976 76090
rect 83924 76026 83976 76032
rect 84292 76084 84344 76090
rect 84292 76026 84344 76032
rect 83280 76016 83332 76022
rect 83280 75958 83332 75964
rect 84304 75954 84332 76026
rect 84292 75948 84344 75954
rect 84292 75890 84344 75896
rect 84384 75200 84436 75206
rect 84384 75142 84436 75148
rect 84396 75002 84424 75142
rect 82176 74996 82228 75002
rect 82176 74938 82228 74944
rect 82820 74996 82872 75002
rect 82820 74938 82872 74944
rect 84384 74996 84436 75002
rect 84384 74938 84436 74944
rect 85592 74254 85620 76230
rect 86788 76090 86816 76842
rect 86880 76498 86908 76978
rect 86868 76492 86920 76498
rect 86868 76434 86920 76440
rect 86960 76356 87012 76362
rect 86960 76298 87012 76304
rect 86684 76084 86736 76090
rect 86684 76026 86736 76032
rect 86776 76084 86828 76090
rect 86776 76026 86828 76032
rect 86696 75886 86724 76026
rect 86684 75880 86736 75886
rect 86684 75822 86736 75828
rect 86592 75812 86644 75818
rect 86592 75754 86644 75760
rect 86316 75744 86368 75750
rect 86316 75686 86368 75692
rect 85580 74248 85632 74254
rect 85580 74190 85632 74196
rect 82084 72616 82136 72622
rect 82084 72558 82136 72564
rect 78036 71052 78088 71058
rect 78036 70994 78088 71000
rect 78048 70650 78076 70994
rect 78036 70644 78088 70650
rect 78036 70586 78088 70592
rect 77208 70440 77260 70446
rect 77208 70382 77260 70388
rect 74356 68740 74408 68746
rect 74356 68682 74408 68688
rect 82096 66842 82124 72558
rect 85672 70440 85724 70446
rect 85672 70382 85724 70388
rect 85488 68332 85540 68338
rect 85488 68274 85540 68280
rect 85500 67726 85528 68274
rect 84384 67720 84436 67726
rect 84384 67662 84436 67668
rect 85488 67720 85540 67726
rect 85488 67662 85540 67668
rect 84396 67250 84424 67662
rect 84384 67244 84436 67250
rect 84384 67186 84436 67192
rect 84384 67040 84436 67046
rect 84384 66982 84436 66988
rect 85580 67040 85632 67046
rect 85580 66982 85632 66988
rect 82084 66836 82136 66842
rect 82084 66778 82136 66784
rect 84396 66570 84424 66982
rect 84292 66564 84344 66570
rect 84292 66506 84344 66512
rect 84384 66564 84436 66570
rect 84384 66506 84436 66512
rect 84304 66298 84332 66506
rect 84292 66292 84344 66298
rect 84292 66234 84344 66240
rect 85592 66230 85620 66982
rect 36084 66224 36136 66230
rect 36082 66192 36084 66201
rect 37924 66224 37976 66230
rect 36136 66192 36138 66201
rect 38476 66224 38528 66230
rect 37924 66166 37976 66172
rect 38474 66192 38476 66201
rect 41144 66224 41196 66230
rect 38528 66192 38530 66201
rect 36082 66127 36138 66136
rect 38474 66127 38530 66136
rect 41142 66192 41144 66201
rect 43628 66224 43680 66230
rect 41196 66192 41198 66201
rect 41142 66127 41198 66136
rect 43626 66192 43628 66201
rect 46112 66224 46164 66230
rect 43680 66192 43682 66201
rect 43626 66127 43682 66136
rect 46110 66192 46112 66201
rect 48596 66224 48648 66230
rect 46164 66192 46166 66201
rect 46110 66127 46166 66136
rect 48594 66192 48596 66201
rect 51080 66224 51132 66230
rect 48648 66192 48650 66201
rect 48594 66127 48650 66136
rect 51078 66192 51080 66201
rect 53564 66224 53616 66230
rect 51132 66192 51134 66201
rect 51078 66127 51134 66136
rect 53562 66192 53564 66201
rect 56140 66224 56192 66230
rect 53616 66192 53618 66201
rect 53562 66127 53618 66136
rect 56138 66192 56140 66201
rect 58624 66224 58676 66230
rect 56192 66192 56194 66201
rect 56138 66127 56194 66136
rect 58622 66192 58624 66201
rect 61108 66224 61160 66230
rect 58676 66192 58678 66201
rect 58622 66127 58678 66136
rect 61106 66192 61108 66201
rect 63592 66224 63644 66230
rect 61160 66192 61162 66201
rect 61106 66127 61162 66136
rect 63590 66192 63592 66201
rect 66076 66224 66128 66230
rect 63644 66192 63646 66201
rect 63590 66127 63646 66136
rect 66074 66192 66076 66201
rect 68560 66224 68612 66230
rect 66128 66192 66130 66201
rect 66074 66127 66130 66136
rect 68558 66192 68560 66201
rect 71044 66224 71096 66230
rect 68612 66192 68614 66201
rect 68558 66127 68614 66136
rect 71042 66192 71044 66201
rect 73528 66224 73580 66230
rect 71096 66192 71098 66201
rect 71042 66127 71098 66136
rect 73526 66192 73528 66201
rect 85580 66224 85632 66230
rect 73580 66192 73582 66201
rect 85580 66166 85632 66172
rect 85684 66162 85712 70382
rect 86328 66201 86356 75686
rect 86604 75342 86632 75754
rect 86696 75546 86724 75822
rect 86684 75540 86736 75546
rect 86684 75482 86736 75488
rect 86972 75410 87000 76298
rect 87064 75886 87092 77862
rect 87340 77654 87368 77998
rect 87328 77648 87380 77654
rect 87328 77590 87380 77596
rect 87236 77444 87288 77450
rect 87236 77386 87288 77392
rect 87248 76838 87276 77386
rect 88904 77178 88932 78950
rect 89812 78464 89864 78470
rect 89812 78406 89864 78412
rect 88984 78124 89036 78130
rect 88984 78066 89036 78072
rect 88996 77450 89024 78066
rect 89076 77580 89128 77586
rect 89076 77522 89128 77528
rect 88984 77444 89036 77450
rect 88984 77386 89036 77392
rect 88432 77172 88484 77178
rect 88432 77114 88484 77120
rect 88892 77172 88944 77178
rect 88892 77114 88944 77120
rect 87236 76832 87288 76838
rect 87236 76774 87288 76780
rect 87144 76288 87196 76294
rect 87144 76230 87196 76236
rect 87052 75880 87104 75886
rect 87052 75822 87104 75828
rect 86960 75404 87012 75410
rect 86960 75346 87012 75352
rect 86592 75336 86644 75342
rect 86592 75278 86644 75284
rect 87064 75206 87092 75822
rect 87156 75274 87184 76230
rect 87248 76022 87276 76774
rect 88444 76430 88472 77114
rect 88524 77104 88576 77110
rect 88524 77046 88576 77052
rect 88536 76634 88564 77046
rect 88984 77036 89036 77042
rect 88984 76978 89036 76984
rect 88996 76634 89024 76978
rect 88524 76628 88576 76634
rect 88524 76570 88576 76576
rect 88984 76628 89036 76634
rect 88984 76570 89036 76576
rect 88432 76424 88484 76430
rect 88432 76366 88484 76372
rect 87236 76016 87288 76022
rect 87236 75958 87288 75964
rect 87420 76016 87472 76022
rect 87420 75958 87472 75964
rect 87432 75478 87460 75958
rect 89088 75886 89116 77522
rect 89720 77444 89772 77450
rect 89720 77386 89772 77392
rect 89444 77376 89496 77382
rect 89444 77318 89496 77324
rect 89456 77042 89484 77318
rect 89444 77036 89496 77042
rect 89444 76978 89496 76984
rect 89732 76566 89760 77386
rect 89824 76974 89852 78406
rect 90546 77208 90602 77217
rect 90546 77143 90602 77152
rect 89812 76968 89864 76974
rect 89812 76910 89864 76916
rect 89904 76832 89956 76838
rect 89904 76774 89956 76780
rect 89720 76560 89772 76566
rect 89720 76502 89772 76508
rect 89168 76424 89220 76430
rect 89168 76366 89220 76372
rect 89720 76424 89772 76430
rect 89720 76366 89772 76372
rect 89180 76294 89208 76366
rect 89732 76294 89760 76366
rect 89168 76288 89220 76294
rect 89168 76230 89220 76236
rect 89720 76288 89772 76294
rect 89720 76230 89772 76236
rect 88708 75880 88760 75886
rect 88708 75822 88760 75828
rect 89076 75880 89128 75886
rect 89076 75822 89128 75828
rect 88720 75546 88748 75822
rect 88708 75540 88760 75546
rect 88708 75482 88760 75488
rect 87420 75472 87472 75478
rect 87420 75414 87472 75420
rect 87144 75268 87196 75274
rect 87144 75210 87196 75216
rect 87052 75200 87104 75206
rect 87052 75142 87104 75148
rect 87156 70990 87184 75210
rect 87696 71936 87748 71942
rect 87696 71878 87748 71884
rect 87144 70984 87196 70990
rect 87144 70926 87196 70932
rect 87708 69057 87736 71878
rect 88720 71058 88748 75482
rect 88984 73296 89036 73302
rect 88984 73238 89036 73244
rect 88708 71052 88760 71058
rect 88708 70994 88760 71000
rect 87880 70984 87932 70990
rect 87880 70926 87932 70932
rect 87694 69048 87750 69057
rect 87694 68983 87750 68992
rect 87892 68746 87920 70926
rect 87880 68740 87932 68746
rect 87880 68682 87932 68688
rect 88248 68740 88300 68746
rect 88248 68682 88300 68688
rect 88260 68338 88288 68682
rect 88248 68332 88300 68338
rect 88248 68274 88300 68280
rect 86960 68128 87012 68134
rect 86960 68070 87012 68076
rect 86972 66570 87000 68070
rect 88432 67720 88484 67726
rect 88432 67662 88484 67668
rect 87052 67652 87104 67658
rect 87052 67594 87104 67600
rect 87064 67250 87092 67594
rect 87052 67244 87104 67250
rect 87052 67186 87104 67192
rect 88444 67046 88472 67662
rect 88720 67386 88748 70994
rect 88996 70922 89024 73238
rect 88984 70916 89036 70922
rect 88984 70858 89036 70864
rect 89180 69222 89208 76230
rect 89916 75954 89944 76774
rect 89904 75948 89956 75954
rect 89904 75890 89956 75896
rect 89916 75546 89944 75890
rect 90180 75744 90232 75750
rect 90180 75686 90232 75692
rect 90456 75744 90508 75750
rect 90456 75686 90508 75692
rect 89904 75540 89956 75546
rect 89904 75482 89956 75488
rect 90192 73166 90220 75686
rect 90364 75540 90416 75546
rect 90364 75482 90416 75488
rect 90272 73296 90324 73302
rect 90272 73238 90324 73244
rect 90180 73160 90232 73166
rect 90180 73102 90232 73108
rect 90284 70394 90312 73238
rect 90376 72010 90404 75482
rect 90468 75342 90496 75686
rect 90456 75336 90508 75342
rect 90456 75278 90508 75284
rect 90456 75200 90508 75206
rect 90456 75142 90508 75148
rect 90468 73166 90496 75142
rect 90456 73160 90508 73166
rect 90456 73102 90508 73108
rect 90364 72004 90416 72010
rect 90364 71946 90416 71952
rect 90192 70366 90312 70394
rect 88984 69216 89036 69222
rect 88984 69158 89036 69164
rect 89168 69216 89220 69222
rect 89168 69158 89220 69164
rect 88996 68950 89024 69158
rect 88984 68944 89036 68950
rect 88984 68886 89036 68892
rect 89812 68944 89864 68950
rect 89812 68886 89864 68892
rect 88996 68814 89024 68886
rect 89824 68814 89852 68886
rect 88984 68808 89036 68814
rect 88984 68750 89036 68756
rect 89812 68808 89864 68814
rect 89812 68750 89864 68756
rect 89812 67720 89864 67726
rect 89812 67662 89864 67668
rect 89352 67652 89404 67658
rect 89352 67594 89404 67600
rect 88708 67380 88760 67386
rect 88708 67322 88760 67328
rect 89168 67312 89220 67318
rect 89168 67254 89220 67260
rect 88708 67244 88760 67250
rect 88708 67186 88760 67192
rect 88432 67040 88484 67046
rect 88432 66982 88484 66988
rect 88156 66700 88208 66706
rect 88156 66642 88208 66648
rect 86960 66564 87012 66570
rect 86960 66506 87012 66512
rect 87604 66224 87656 66230
rect 86314 66192 86370 66201
rect 73526 66127 73582 66136
rect 85672 66156 85724 66162
rect 87604 66166 87656 66172
rect 86314 66127 86370 66136
rect 85672 66098 85724 66104
rect 87616 66094 87644 66166
rect 88168 66162 88196 66642
rect 88444 66298 88472 66982
rect 88720 66502 88748 67186
rect 88892 67040 88944 67046
rect 88892 66982 88944 66988
rect 88904 66570 88932 66982
rect 89180 66706 89208 67254
rect 89364 67250 89392 67594
rect 89720 67380 89772 67386
rect 89720 67322 89772 67328
rect 89352 67244 89404 67250
rect 89536 67244 89588 67250
rect 89352 67186 89404 67192
rect 89456 67204 89536 67232
rect 89260 67176 89312 67182
rect 89260 67118 89312 67124
rect 89272 66842 89300 67118
rect 89260 66836 89312 66842
rect 89260 66778 89312 66784
rect 89352 66768 89404 66774
rect 89352 66710 89404 66716
rect 89168 66700 89220 66706
rect 89168 66642 89220 66648
rect 89260 66632 89312 66638
rect 89260 66574 89312 66580
rect 88892 66564 88944 66570
rect 88892 66506 88944 66512
rect 88984 66564 89036 66570
rect 88984 66506 89036 66512
rect 88708 66496 88760 66502
rect 88708 66438 88760 66444
rect 88432 66292 88484 66298
rect 88432 66234 88484 66240
rect 88156 66156 88208 66162
rect 88156 66098 88208 66104
rect 87604 66088 87656 66094
rect 88064 66088 88116 66094
rect 87604 66030 87656 66036
rect 87892 66036 88064 66042
rect 87892 66030 88116 66036
rect 87892 66014 88104 66030
rect 87892 65958 87920 66014
rect 86224 65952 86276 65958
rect 86224 65894 86276 65900
rect 87880 65952 87932 65958
rect 87880 65894 87932 65900
rect 34934 65852 35242 65861
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65787 35242 65796
rect 65654 65852 65962 65861
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65787 65962 65796
rect 86236 65754 86264 65894
rect 86224 65748 86276 65754
rect 86224 65690 86276 65696
rect 88444 65686 88472 66234
rect 88996 66094 89024 66506
rect 88984 66088 89036 66094
rect 88984 66030 89036 66036
rect 89272 66026 89300 66574
rect 89364 66570 89392 66710
rect 89352 66564 89404 66570
rect 89352 66506 89404 66512
rect 89364 66201 89392 66506
rect 89456 66337 89484 67204
rect 89536 67186 89588 67192
rect 89732 66502 89760 67322
rect 89824 67046 89852 67662
rect 89996 67584 90048 67590
rect 89996 67526 90048 67532
rect 89904 67108 89956 67114
rect 89904 67050 89956 67056
rect 89812 67040 89864 67046
rect 89812 66982 89864 66988
rect 89720 66496 89772 66502
rect 89720 66438 89772 66444
rect 89442 66328 89498 66337
rect 89442 66263 89444 66272
rect 89496 66263 89498 66272
rect 89720 66292 89772 66298
rect 89444 66234 89496 66240
rect 89720 66234 89772 66240
rect 89350 66192 89406 66201
rect 89350 66127 89406 66136
rect 89364 66026 89392 66127
rect 89444 66088 89496 66094
rect 89444 66030 89496 66036
rect 89260 66020 89312 66026
rect 89260 65962 89312 65968
rect 89352 66020 89404 66026
rect 89352 65962 89404 65968
rect 89456 65906 89484 66030
rect 89732 65906 89760 66234
rect 89456 65878 89760 65906
rect 88432 65680 88484 65686
rect 88432 65622 88484 65628
rect 89824 65550 89852 66982
rect 89916 66706 89944 67050
rect 89904 66700 89956 66706
rect 89904 66642 89956 66648
rect 89916 66298 89944 66642
rect 90008 66638 90036 67526
rect 90192 67386 90220 70366
rect 90560 67930 90588 77143
rect 90652 73302 90680 79863
rect 90914 79520 90970 79529
rect 90914 79455 90970 79464
rect 90732 77920 90784 77926
rect 90732 77862 90784 77868
rect 90744 77654 90772 77862
rect 90732 77648 90784 77654
rect 90732 77590 90784 77596
rect 90732 75948 90784 75954
rect 90732 75890 90784 75896
rect 90744 75206 90772 75890
rect 90824 75268 90876 75274
rect 90824 75210 90876 75216
rect 90732 75200 90784 75206
rect 90732 75142 90784 75148
rect 90640 73296 90692 73302
rect 90640 73238 90692 73244
rect 90640 73160 90692 73166
rect 90640 73102 90692 73108
rect 90652 68814 90680 73102
rect 90744 71738 90772 75142
rect 90836 72078 90864 75210
rect 90824 72072 90876 72078
rect 90824 72014 90876 72020
rect 90732 71732 90784 71738
rect 90732 71674 90784 71680
rect 90640 68808 90692 68814
rect 90640 68750 90692 68756
rect 90732 68128 90784 68134
rect 90732 68070 90784 68076
rect 90548 67924 90600 67930
rect 90548 67866 90600 67872
rect 90548 67720 90600 67726
rect 90548 67662 90600 67668
rect 90180 67380 90232 67386
rect 90180 67322 90232 67328
rect 90272 67176 90324 67182
rect 90272 67118 90324 67124
rect 90284 66638 90312 67118
rect 89996 66632 90048 66638
rect 89996 66574 90048 66580
rect 90272 66632 90324 66638
rect 90272 66574 90324 66580
rect 90008 66502 90036 66574
rect 90560 66570 90588 67662
rect 90744 67318 90772 68070
rect 90732 67312 90784 67318
rect 90732 67254 90784 67260
rect 90640 66768 90692 66774
rect 90640 66710 90692 66716
rect 90652 66638 90680 66710
rect 90640 66632 90692 66638
rect 90640 66574 90692 66580
rect 90548 66564 90600 66570
rect 90548 66506 90600 66512
rect 89996 66496 90048 66502
rect 89996 66438 90048 66444
rect 90456 66496 90508 66502
rect 90456 66438 90508 66444
rect 90008 66298 90036 66438
rect 89904 66292 89956 66298
rect 89904 66234 89956 66240
rect 89996 66292 90048 66298
rect 89996 66234 90048 66240
rect 90468 66230 90496 66438
rect 90456 66224 90508 66230
rect 90456 66166 90508 66172
rect 90364 66156 90416 66162
rect 90364 66098 90416 66104
rect 90376 65754 90404 66098
rect 90560 65754 90588 66506
rect 90732 66292 90784 66298
rect 90732 66234 90784 66240
rect 90744 66094 90772 66234
rect 90928 66230 90956 79455
rect 101968 79354 101996 136206
rect 106658 136028 106966 136037
rect 106658 136026 106664 136028
rect 106720 136026 106744 136028
rect 106800 136026 106824 136028
rect 106880 136026 106904 136028
rect 106960 136026 106966 136028
rect 106720 135974 106722 136026
rect 106902 135974 106904 136026
rect 106658 135972 106664 135974
rect 106720 135972 106744 135974
rect 106800 135972 106824 135974
rect 106880 135972 106904 135974
rect 106960 135972 106966 135974
rect 106658 135963 106966 135972
rect 102140 135924 102192 135930
rect 102140 135866 102192 135872
rect 101956 79348 102008 79354
rect 101956 79290 102008 79296
rect 102152 78606 102180 135866
rect 103980 135856 104032 135862
rect 103980 135798 104032 135804
rect 102324 135788 102376 135794
rect 102324 135730 102376 135736
rect 102232 134020 102284 134026
rect 102232 133962 102284 133968
rect 96528 78600 96580 78606
rect 96526 78568 96528 78577
rect 102140 78600 102192 78606
rect 96580 78568 96582 78577
rect 91652 78532 91704 78538
rect 102140 78542 102192 78548
rect 96526 78503 96582 78512
rect 91652 78474 91704 78480
rect 91664 77450 91692 78474
rect 93124 78056 93176 78062
rect 93124 77998 93176 78004
rect 93136 77654 93164 77998
rect 94228 77988 94280 77994
rect 94228 77930 94280 77936
rect 93124 77648 93176 77654
rect 93124 77590 93176 77596
rect 94240 77450 94268 77930
rect 99656 77920 99708 77926
rect 99656 77862 99708 77868
rect 96374 77820 96682 77829
rect 96374 77818 96380 77820
rect 96436 77818 96460 77820
rect 96516 77818 96540 77820
rect 96596 77818 96620 77820
rect 96676 77818 96682 77820
rect 96436 77766 96438 77818
rect 96618 77766 96620 77818
rect 96374 77764 96380 77766
rect 96436 77764 96460 77766
rect 96516 77764 96540 77766
rect 96596 77764 96620 77766
rect 96676 77764 96682 77766
rect 96374 77755 96682 77764
rect 99668 77586 99696 77862
rect 99656 77580 99708 77586
rect 99656 77522 99708 77528
rect 91652 77444 91704 77450
rect 91652 77386 91704 77392
rect 92664 77444 92716 77450
rect 92664 77386 92716 77392
rect 94228 77444 94280 77450
rect 94228 77386 94280 77392
rect 95240 77444 95292 77450
rect 95240 77386 95292 77392
rect 92020 77376 92072 77382
rect 92020 77318 92072 77324
rect 92032 77178 92060 77318
rect 92020 77172 92072 77178
rect 92020 77114 92072 77120
rect 91468 77036 91520 77042
rect 91468 76978 91520 76984
rect 91480 76838 91508 76978
rect 91468 76832 91520 76838
rect 91468 76774 91520 76780
rect 91480 76294 91508 76774
rect 92676 76634 92704 77386
rect 95252 77110 95280 77386
rect 97034 77276 97342 77285
rect 97034 77274 97040 77276
rect 97096 77274 97120 77276
rect 97176 77274 97200 77276
rect 97256 77274 97280 77276
rect 97336 77274 97342 77276
rect 97096 77222 97098 77274
rect 97278 77222 97280 77274
rect 97034 77220 97040 77222
rect 97096 77220 97120 77222
rect 97176 77220 97200 77222
rect 97256 77220 97280 77222
rect 97336 77220 97342 77222
rect 97034 77211 97342 77220
rect 95240 77104 95292 77110
rect 95240 77046 95292 77052
rect 96374 76732 96682 76741
rect 96374 76730 96380 76732
rect 96436 76730 96460 76732
rect 96516 76730 96540 76732
rect 96596 76730 96620 76732
rect 96676 76730 96682 76732
rect 96436 76678 96438 76730
rect 96618 76678 96620 76730
rect 96374 76676 96380 76678
rect 96436 76676 96460 76678
rect 96516 76676 96540 76678
rect 96596 76676 96620 76678
rect 96676 76676 96682 76678
rect 96374 76667 96682 76676
rect 92664 76628 92716 76634
rect 92664 76570 92716 76576
rect 102244 76498 102272 133962
rect 102336 77625 102364 135730
rect 102416 135720 102468 135726
rect 102416 135662 102468 135668
rect 102428 78266 102456 135662
rect 103612 135652 103664 135658
rect 103612 135594 103664 135600
rect 102508 135516 102560 135522
rect 102508 135458 102560 135464
rect 102520 78305 102548 135458
rect 103520 134564 103572 134570
rect 103520 134506 103572 134512
rect 102600 133952 102652 133958
rect 102600 133894 102652 133900
rect 102506 78296 102562 78305
rect 102416 78260 102468 78266
rect 102506 78231 102562 78240
rect 102416 78202 102468 78208
rect 102612 78130 102640 133894
rect 102692 95328 102744 95334
rect 102692 95270 102744 95276
rect 102704 95033 102732 95270
rect 102690 95024 102746 95033
rect 102690 94959 102746 94968
rect 102600 78124 102652 78130
rect 102600 78066 102652 78072
rect 102322 77616 102378 77625
rect 102322 77551 102378 77560
rect 102232 76492 102284 76498
rect 102232 76434 102284 76440
rect 91468 76288 91520 76294
rect 91468 76230 91520 76236
rect 97034 76188 97342 76197
rect 97034 76186 97040 76188
rect 97096 76186 97120 76188
rect 97176 76186 97200 76188
rect 97256 76186 97280 76188
rect 97336 76186 97342 76188
rect 97096 76134 97098 76186
rect 97278 76134 97280 76186
rect 97034 76132 97040 76134
rect 97096 76132 97120 76134
rect 97176 76132 97200 76134
rect 97256 76132 97280 76134
rect 97336 76132 97342 76134
rect 97034 76123 97342 76132
rect 102704 75818 102732 94959
rect 103060 93900 103112 93906
rect 102888 93848 103060 93854
rect 102888 93842 103112 93848
rect 102888 93826 103100 93842
rect 102888 93401 102916 93826
rect 102874 93392 102930 93401
rect 102874 93327 102930 93336
rect 102692 75812 102744 75818
rect 102692 75754 102744 75760
rect 96374 75644 96682 75653
rect 96374 75642 96380 75644
rect 96436 75642 96460 75644
rect 96516 75642 96540 75644
rect 96596 75642 96620 75644
rect 96676 75642 96682 75644
rect 96436 75590 96438 75642
rect 96618 75590 96620 75642
rect 96374 75588 96380 75590
rect 96436 75588 96460 75590
rect 96516 75588 96540 75590
rect 96596 75588 96620 75590
rect 96676 75588 96682 75590
rect 96374 75579 96682 75588
rect 97034 75100 97342 75109
rect 97034 75098 97040 75100
rect 97096 75098 97120 75100
rect 97176 75098 97200 75100
rect 97256 75098 97280 75100
rect 97336 75098 97342 75100
rect 97096 75046 97098 75098
rect 97278 75046 97280 75098
rect 97034 75044 97040 75046
rect 97096 75044 97120 75046
rect 97176 75044 97200 75046
rect 97256 75044 97280 75046
rect 97336 75044 97342 75046
rect 97034 75035 97342 75044
rect 102140 74996 102192 75002
rect 102140 74938 102192 74944
rect 96374 74556 96682 74565
rect 96374 74554 96380 74556
rect 96436 74554 96460 74556
rect 96516 74554 96540 74556
rect 96596 74554 96620 74556
rect 96676 74554 96682 74556
rect 96436 74502 96438 74554
rect 96618 74502 96620 74554
rect 96374 74500 96380 74502
rect 96436 74500 96460 74502
rect 96516 74500 96540 74502
rect 96596 74500 96620 74502
rect 96676 74500 96682 74502
rect 96374 74491 96682 74500
rect 97034 74012 97342 74021
rect 97034 74010 97040 74012
rect 97096 74010 97120 74012
rect 97176 74010 97200 74012
rect 97256 74010 97280 74012
rect 97336 74010 97342 74012
rect 97096 73958 97098 74010
rect 97278 73958 97280 74010
rect 97034 73956 97040 73958
rect 97096 73956 97120 73958
rect 97176 73956 97200 73958
rect 97256 73956 97280 73958
rect 97336 73956 97342 73958
rect 97034 73947 97342 73956
rect 102152 73574 102180 74938
rect 102140 73568 102192 73574
rect 102140 73510 102192 73516
rect 96374 73468 96682 73477
rect 96374 73466 96380 73468
rect 96436 73466 96460 73468
rect 96516 73466 96540 73468
rect 96596 73466 96620 73468
rect 96676 73466 96682 73468
rect 96436 73414 96438 73466
rect 96618 73414 96620 73466
rect 96374 73412 96380 73414
rect 96436 73412 96460 73414
rect 96516 73412 96540 73414
rect 96596 73412 96620 73414
rect 96676 73412 96682 73414
rect 96374 73403 96682 73412
rect 97034 72924 97342 72933
rect 97034 72922 97040 72924
rect 97096 72922 97120 72924
rect 97176 72922 97200 72924
rect 97256 72922 97280 72924
rect 97336 72922 97342 72924
rect 97096 72870 97098 72922
rect 97278 72870 97280 72922
rect 97034 72868 97040 72870
rect 97096 72868 97120 72870
rect 97176 72868 97200 72870
rect 97256 72868 97280 72870
rect 97336 72868 97342 72870
rect 97034 72859 97342 72868
rect 95148 72480 95200 72486
rect 95148 72422 95200 72428
rect 95160 72282 95188 72422
rect 96374 72380 96682 72389
rect 96374 72378 96380 72380
rect 96436 72378 96460 72380
rect 96516 72378 96540 72380
rect 96596 72378 96620 72380
rect 96676 72378 96682 72380
rect 96436 72326 96438 72378
rect 96618 72326 96620 72378
rect 96374 72324 96380 72326
rect 96436 72324 96460 72326
rect 96516 72324 96540 72326
rect 96596 72324 96620 72326
rect 96676 72324 96682 72326
rect 96374 72315 96682 72324
rect 94320 72276 94372 72282
rect 94320 72218 94372 72224
rect 95148 72276 95200 72282
rect 95148 72218 95200 72224
rect 92388 72004 92440 72010
rect 92388 71946 92440 71952
rect 91836 71936 91888 71942
rect 91836 71878 91888 71884
rect 92112 71936 92164 71942
rect 92112 71878 92164 71884
rect 91848 71602 91876 71878
rect 91100 71596 91152 71602
rect 91100 71538 91152 71544
rect 91836 71596 91888 71602
rect 91836 71538 91888 71544
rect 91112 71194 91140 71538
rect 91100 71188 91152 71194
rect 91100 71130 91152 71136
rect 91100 68672 91152 68678
rect 91100 68614 91152 68620
rect 91112 67726 91140 68614
rect 92124 67794 92152 71878
rect 92400 68814 92428 71946
rect 92388 68808 92440 68814
rect 92388 68750 92440 68756
rect 91560 67788 91612 67794
rect 91560 67730 91612 67736
rect 92112 67788 92164 67794
rect 92112 67730 92164 67736
rect 91100 67720 91152 67726
rect 91100 67662 91152 67668
rect 91100 67584 91152 67590
rect 91100 67526 91152 67532
rect 91112 67386 91140 67526
rect 91100 67380 91152 67386
rect 91100 67322 91152 67328
rect 91572 67182 91600 67730
rect 92400 67726 92428 68750
rect 92388 67720 92440 67726
rect 92388 67662 92440 67668
rect 92400 67386 92428 67662
rect 92388 67380 92440 67386
rect 92388 67322 92440 67328
rect 91560 67176 91612 67182
rect 91560 67118 91612 67124
rect 91284 66632 91336 66638
rect 91284 66574 91336 66580
rect 91376 66632 91428 66638
rect 91376 66574 91428 66580
rect 91006 66328 91062 66337
rect 91006 66263 91008 66272
rect 91060 66263 91062 66272
rect 91008 66234 91060 66240
rect 90916 66224 90968 66230
rect 90916 66166 90968 66172
rect 91192 66156 91244 66162
rect 91192 66098 91244 66104
rect 90640 66088 90692 66094
rect 90640 66030 90692 66036
rect 90732 66088 90784 66094
rect 90732 66030 90784 66036
rect 90652 65958 90680 66030
rect 90640 65952 90692 65958
rect 90640 65894 90692 65900
rect 90364 65748 90416 65754
rect 90364 65690 90416 65696
rect 90548 65748 90600 65754
rect 90548 65690 90600 65696
rect 91204 65686 91232 66098
rect 91296 65958 91324 66574
rect 91388 66298 91416 66574
rect 91376 66292 91428 66298
rect 91376 66234 91428 66240
rect 91572 66230 91600 67118
rect 91928 66496 91980 66502
rect 91928 66438 91980 66444
rect 91940 66298 91968 66438
rect 91928 66292 91980 66298
rect 91928 66234 91980 66240
rect 94332 66230 94360 72218
rect 102888 72010 102916 93327
rect 102968 92608 103020 92614
rect 102968 92550 103020 92556
rect 102980 92313 103008 92550
rect 102966 92304 103022 92313
rect 102966 92239 103022 92248
rect 102876 72004 102928 72010
rect 102876 71946 102928 71952
rect 97034 71836 97342 71845
rect 97034 71834 97040 71836
rect 97096 71834 97120 71836
rect 97176 71834 97200 71836
rect 97256 71834 97280 71836
rect 97336 71834 97342 71836
rect 97096 71782 97098 71834
rect 97278 71782 97280 71834
rect 97034 71780 97040 71782
rect 97096 71780 97120 71782
rect 97176 71780 97200 71782
rect 97256 71780 97280 71782
rect 97336 71780 97342 71782
rect 97034 71771 97342 71780
rect 102232 71392 102284 71398
rect 102232 71334 102284 71340
rect 96374 71292 96682 71301
rect 96374 71290 96380 71292
rect 96436 71290 96460 71292
rect 96516 71290 96540 71292
rect 96596 71290 96620 71292
rect 96676 71290 96682 71292
rect 96436 71238 96438 71290
rect 96618 71238 96620 71290
rect 96374 71236 96380 71238
rect 96436 71236 96460 71238
rect 96516 71236 96540 71238
rect 96596 71236 96620 71238
rect 96676 71236 96682 71238
rect 96374 71227 96682 71236
rect 97034 70748 97342 70757
rect 97034 70746 97040 70748
rect 97096 70746 97120 70748
rect 97176 70746 97200 70748
rect 97256 70746 97280 70748
rect 97336 70746 97342 70748
rect 97096 70694 97098 70746
rect 97278 70694 97280 70746
rect 97034 70692 97040 70694
rect 97096 70692 97120 70694
rect 97176 70692 97200 70694
rect 97256 70692 97280 70694
rect 97336 70692 97342 70694
rect 97034 70683 97342 70692
rect 96374 70204 96682 70213
rect 96374 70202 96380 70204
rect 96436 70202 96460 70204
rect 96516 70202 96540 70204
rect 96596 70202 96620 70204
rect 96676 70202 96682 70204
rect 96436 70150 96438 70202
rect 96618 70150 96620 70202
rect 96374 70148 96380 70150
rect 96436 70148 96460 70150
rect 96516 70148 96540 70150
rect 96596 70148 96620 70150
rect 96676 70148 96682 70150
rect 96374 70139 96682 70148
rect 97034 69660 97342 69669
rect 97034 69658 97040 69660
rect 97096 69658 97120 69660
rect 97176 69658 97200 69660
rect 97256 69658 97280 69660
rect 97336 69658 97342 69660
rect 97096 69606 97098 69658
rect 97278 69606 97280 69658
rect 97034 69604 97040 69606
rect 97096 69604 97120 69606
rect 97176 69604 97200 69606
rect 97256 69604 97280 69606
rect 97336 69604 97342 69606
rect 97034 69595 97342 69604
rect 96374 69116 96682 69125
rect 96374 69114 96380 69116
rect 96436 69114 96460 69116
rect 96516 69114 96540 69116
rect 96596 69114 96620 69116
rect 96676 69114 96682 69116
rect 96436 69062 96438 69114
rect 96618 69062 96620 69114
rect 96374 69060 96380 69062
rect 96436 69060 96460 69062
rect 96516 69060 96540 69062
rect 96596 69060 96620 69062
rect 96676 69060 96682 69062
rect 96374 69051 96682 69060
rect 97034 68572 97342 68581
rect 97034 68570 97040 68572
rect 97096 68570 97120 68572
rect 97176 68570 97200 68572
rect 97256 68570 97280 68572
rect 97336 68570 97342 68572
rect 97096 68518 97098 68570
rect 97278 68518 97280 68570
rect 97034 68516 97040 68518
rect 97096 68516 97120 68518
rect 97176 68516 97200 68518
rect 97256 68516 97280 68518
rect 97336 68516 97342 68518
rect 97034 68507 97342 68516
rect 96374 68028 96682 68037
rect 96374 68026 96380 68028
rect 96436 68026 96460 68028
rect 96516 68026 96540 68028
rect 96596 68026 96620 68028
rect 96676 68026 96682 68028
rect 96436 67974 96438 68026
rect 96618 67974 96620 68026
rect 96374 67972 96380 67974
rect 96436 67972 96460 67974
rect 96516 67972 96540 67974
rect 96596 67972 96620 67974
rect 96676 67972 96682 67974
rect 96374 67963 96682 67972
rect 101956 67856 102008 67862
rect 101956 67798 102008 67804
rect 97034 67484 97342 67493
rect 97034 67482 97040 67484
rect 97096 67482 97120 67484
rect 97176 67482 97200 67484
rect 97256 67482 97280 67484
rect 97336 67482 97342 67484
rect 97096 67430 97098 67482
rect 97278 67430 97280 67482
rect 97034 67428 97040 67430
rect 97096 67428 97120 67430
rect 97176 67428 97200 67430
rect 97256 67428 97280 67430
rect 97336 67428 97342 67430
rect 97034 67419 97342 67428
rect 95884 67040 95936 67046
rect 95884 66982 95936 66988
rect 91560 66224 91612 66230
rect 94320 66224 94372 66230
rect 91560 66166 91612 66172
rect 91926 66192 91982 66201
rect 94320 66166 94372 66172
rect 91926 66127 91928 66136
rect 91980 66127 91982 66136
rect 91928 66098 91980 66104
rect 95896 65958 95924 66982
rect 96374 66940 96682 66949
rect 96374 66938 96380 66940
rect 96436 66938 96460 66940
rect 96516 66938 96540 66940
rect 96596 66938 96620 66940
rect 96676 66938 96682 66940
rect 96436 66886 96438 66938
rect 96618 66886 96620 66938
rect 96374 66884 96380 66886
rect 96436 66884 96460 66886
rect 96516 66884 96540 66886
rect 96596 66884 96620 66886
rect 96676 66884 96682 66886
rect 96374 66875 96682 66884
rect 97034 66396 97342 66405
rect 97034 66394 97040 66396
rect 97096 66394 97120 66396
rect 97176 66394 97200 66396
rect 97256 66394 97280 66396
rect 97336 66394 97342 66396
rect 97096 66342 97098 66394
rect 97278 66342 97280 66394
rect 97034 66340 97040 66342
rect 97096 66340 97120 66342
rect 97176 66340 97200 66342
rect 97256 66340 97280 66342
rect 97336 66340 97342 66342
rect 97034 66331 97342 66340
rect 91284 65952 91336 65958
rect 91284 65894 91336 65900
rect 91560 65952 91612 65958
rect 91560 65894 91612 65900
rect 92296 65952 92348 65958
rect 92296 65894 92348 65900
rect 95884 65952 95936 65958
rect 95884 65894 95936 65900
rect 91572 65754 91600 65894
rect 91560 65748 91612 65754
rect 91560 65690 91612 65696
rect 92308 65686 92336 65894
rect 91192 65680 91244 65686
rect 91192 65622 91244 65628
rect 92296 65680 92348 65686
rect 92296 65622 92348 65628
rect 89812 65544 89864 65550
rect 89812 65486 89864 65492
rect 95896 64161 95924 65894
rect 96374 65852 96682 65861
rect 96374 65850 96380 65852
rect 96436 65850 96460 65852
rect 96516 65850 96540 65852
rect 96596 65850 96620 65852
rect 96676 65850 96682 65852
rect 96436 65798 96438 65850
rect 96618 65798 96620 65850
rect 96374 65796 96380 65798
rect 96436 65796 96460 65798
rect 96516 65796 96540 65798
rect 96596 65796 96620 65798
rect 96676 65796 96682 65798
rect 96374 65787 96682 65796
rect 95882 64152 95938 64161
rect 95882 64087 95938 64096
rect 101968 23866 101996 67798
rect 102140 66292 102192 66298
rect 102140 66234 102192 66240
rect 101956 23860 102008 23866
rect 101956 23802 102008 23808
rect 101968 23374 101996 23802
rect 102046 23388 102102 23397
rect 101968 23346 102046 23374
rect 102046 23323 102102 23332
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 29564 9761 29592 9862
rect 23478 9752 23534 9761
rect 23478 9687 23534 9696
rect 25778 9752 25834 9761
rect 25778 9687 25834 9696
rect 28170 9752 28226 9761
rect 28170 9687 28226 9696
rect 29550 9752 29606 9761
rect 29550 9687 29606 9696
rect 30470 9752 30526 9761
rect 30470 9687 30526 9696
rect 90546 9752 90602 9761
rect 90546 9687 90602 9696
rect 90914 9752 90970 9761
rect 90914 9687 90970 9696
rect 9588 9648 9640 9654
rect 16120 9648 16172 9654
rect 9588 9590 9640 9596
rect 16026 9616 16082 9625
rect 16120 9590 16172 9596
rect 16026 9551 16028 9560
rect 16080 9551 16082 9560
rect 16028 9522 16080 9528
rect 16040 7546 16068 9522
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 1320 4865 1348 5170
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 1306 4856 1362 4865
rect 4214 4859 4522 4868
rect 1306 4791 1362 4800
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 16132 800 16160 9590
rect 23492 7546 23520 9687
rect 24674 9616 24730 9625
rect 24674 9551 24730 9560
rect 24688 8362 24716 9551
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24688 7546 24716 8298
rect 25792 7546 25820 9687
rect 26698 8936 26754 8945
rect 26698 8871 26754 8880
rect 26712 8838 26740 8871
rect 26700 8832 26752 8838
rect 26700 8774 26752 8780
rect 26712 7546 26740 8774
rect 28184 7546 28212 9687
rect 29564 7546 29592 9687
rect 30484 7750 30512 9687
rect 90560 9654 90588 9687
rect 90548 9648 90600 9654
rect 90548 9590 90600 9596
rect 90730 9616 90786 9625
rect 31666 8256 31722 8265
rect 31666 8191 31722 8200
rect 32954 8256 33010 8265
rect 32954 8191 33010 8200
rect 34242 8256 34298 8265
rect 34242 8191 34298 8200
rect 35438 8256 35494 8265
rect 35438 8191 35494 8200
rect 36358 8256 36414 8265
rect 36358 8191 36414 8200
rect 37462 8256 37518 8265
rect 37462 8191 37518 8200
rect 38750 8256 38806 8265
rect 38750 8191 38806 8200
rect 41326 8256 41382 8265
rect 41326 8191 41382 8200
rect 42154 8256 42210 8265
rect 42154 8191 42210 8200
rect 43442 8256 43498 8265
rect 43442 8191 43498 8200
rect 30472 7744 30524 7750
rect 30472 7686 30524 7692
rect 30484 7546 30512 7686
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 26700 7540 26752 7546
rect 26700 7482 26752 7488
rect 28172 7540 28224 7546
rect 28172 7482 28224 7488
rect 29552 7540 29604 7546
rect 29552 7482 29604 7488
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 23492 5030 23520 7482
rect 25792 6914 25820 7482
rect 28184 7274 28212 7482
rect 28172 7268 28224 7274
rect 28172 7210 28224 7216
rect 25792 6886 25912 6914
rect 25884 6118 25912 6886
rect 25872 6112 25924 6118
rect 25872 6054 25924 6060
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 31680 2650 31708 8191
rect 32968 2650 32996 8191
rect 34256 2650 34284 8191
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35452 2650 35480 8191
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 36372 2650 36400 8191
rect 37476 2650 37504 8191
rect 38764 2650 38792 8191
rect 39946 4584 40002 4593
rect 39946 4519 40002 4528
rect 39960 2650 39988 4519
rect 41340 2650 41368 8191
rect 42168 2650 42196 8191
rect 43456 2650 43484 8191
rect 66314 7644 66622 7653
rect 66314 7642 66320 7644
rect 66376 7642 66400 7644
rect 66456 7642 66480 7644
rect 66536 7642 66560 7644
rect 66616 7642 66622 7644
rect 66376 7590 66378 7642
rect 66558 7590 66560 7642
rect 66314 7588 66320 7590
rect 66376 7588 66400 7590
rect 66456 7588 66480 7590
rect 66536 7588 66560 7590
rect 66616 7588 66622 7590
rect 66314 7579 66622 7588
rect 90560 7546 90588 9590
rect 90928 9586 90956 9687
rect 90730 9551 90786 9560
rect 90916 9580 90968 9586
rect 90744 9518 90772 9551
rect 90916 9522 90968 9528
rect 90732 9512 90784 9518
rect 90732 9454 90784 9460
rect 90744 7546 90772 9454
rect 90928 7546 90956 9522
rect 102152 9518 102180 66234
rect 102244 25097 102272 71334
rect 102980 67658 103008 92239
rect 103532 90982 103560 134506
rect 103520 90976 103572 90982
rect 103520 90918 103572 90924
rect 103624 78033 103652 135594
rect 103704 135584 103756 135590
rect 103704 135526 103756 135532
rect 103716 78169 103744 135526
rect 103888 135448 103940 135454
rect 103888 135390 103940 135396
rect 103796 135380 103848 135386
rect 103796 135322 103848 135328
rect 103702 78160 103758 78169
rect 103702 78095 103758 78104
rect 103610 78024 103666 78033
rect 103610 77959 103666 77968
rect 103808 77722 103836 135322
rect 103900 78441 103928 135390
rect 103886 78432 103942 78441
rect 103886 78367 103942 78376
rect 103796 77716 103848 77722
rect 103796 77658 103848 77664
rect 103992 77489 104020 135798
rect 105922 135484 106230 135493
rect 105922 135482 105928 135484
rect 105984 135482 106008 135484
rect 106064 135482 106088 135484
rect 106144 135482 106168 135484
rect 106224 135482 106230 135484
rect 105984 135430 105986 135482
rect 106166 135430 106168 135482
rect 105922 135428 105928 135430
rect 105984 135428 106008 135430
rect 106064 135428 106088 135430
rect 106144 135428 106168 135430
rect 106224 135428 106230 135430
rect 105922 135419 106230 135428
rect 106658 134940 106966 134949
rect 106658 134938 106664 134940
rect 106720 134938 106744 134940
rect 106800 134938 106824 134940
rect 106880 134938 106904 134940
rect 106960 134938 106966 134940
rect 106720 134886 106722 134938
rect 106902 134886 106904 134938
rect 106658 134884 106664 134886
rect 106720 134884 106744 134886
rect 106800 134884 106824 134886
rect 106880 134884 106904 134886
rect 106960 134884 106966 134886
rect 106658 134875 106966 134884
rect 105922 134396 106230 134405
rect 105922 134394 105928 134396
rect 105984 134394 106008 134396
rect 106064 134394 106088 134396
rect 106144 134394 106168 134396
rect 106224 134394 106230 134396
rect 105984 134342 105986 134394
rect 106166 134342 106168 134394
rect 105922 134340 105928 134342
rect 105984 134340 106008 134342
rect 106064 134340 106088 134342
rect 106144 134340 106168 134342
rect 106224 134340 106230 134342
rect 105922 134331 106230 134340
rect 106658 133852 106966 133861
rect 106658 133850 106664 133852
rect 106720 133850 106744 133852
rect 106800 133850 106824 133852
rect 106880 133850 106904 133852
rect 106960 133850 106966 133852
rect 106720 133798 106722 133850
rect 106902 133798 106904 133850
rect 106658 133796 106664 133798
rect 106720 133796 106744 133798
rect 106800 133796 106824 133798
rect 106880 133796 106904 133798
rect 106960 133796 106966 133798
rect 106658 133787 106966 133796
rect 105922 133308 106230 133317
rect 105922 133306 105928 133308
rect 105984 133306 106008 133308
rect 106064 133306 106088 133308
rect 106144 133306 106168 133308
rect 106224 133306 106230 133308
rect 105984 133254 105986 133306
rect 106166 133254 106168 133306
rect 105922 133252 105928 133254
rect 105984 133252 106008 133254
rect 106064 133252 106088 133254
rect 106144 133252 106168 133254
rect 106224 133252 106230 133254
rect 105922 133243 106230 133252
rect 106658 132764 106966 132773
rect 106658 132762 106664 132764
rect 106720 132762 106744 132764
rect 106800 132762 106824 132764
rect 106880 132762 106904 132764
rect 106960 132762 106966 132764
rect 106720 132710 106722 132762
rect 106902 132710 106904 132762
rect 106658 132708 106664 132710
rect 106720 132708 106744 132710
rect 106800 132708 106824 132710
rect 106880 132708 106904 132710
rect 106960 132708 106966 132710
rect 106658 132699 106966 132708
rect 105922 132220 106230 132229
rect 105922 132218 105928 132220
rect 105984 132218 106008 132220
rect 106064 132218 106088 132220
rect 106144 132218 106168 132220
rect 106224 132218 106230 132220
rect 105984 132166 105986 132218
rect 106166 132166 106168 132218
rect 105922 132164 105928 132166
rect 105984 132164 106008 132166
rect 106064 132164 106088 132166
rect 106144 132164 106168 132166
rect 106224 132164 106230 132166
rect 105922 132155 106230 132164
rect 106658 131676 106966 131685
rect 106658 131674 106664 131676
rect 106720 131674 106744 131676
rect 106800 131674 106824 131676
rect 106880 131674 106904 131676
rect 106960 131674 106966 131676
rect 106720 131622 106722 131674
rect 106902 131622 106904 131674
rect 106658 131620 106664 131622
rect 106720 131620 106744 131622
rect 106800 131620 106824 131622
rect 106880 131620 106904 131622
rect 106960 131620 106966 131622
rect 106658 131611 106966 131620
rect 105922 131132 106230 131141
rect 105922 131130 105928 131132
rect 105984 131130 106008 131132
rect 106064 131130 106088 131132
rect 106144 131130 106168 131132
rect 106224 131130 106230 131132
rect 105984 131078 105986 131130
rect 106166 131078 106168 131130
rect 105922 131076 105928 131078
rect 105984 131076 106008 131078
rect 106064 131076 106088 131078
rect 106144 131076 106168 131078
rect 106224 131076 106230 131078
rect 105922 131067 106230 131076
rect 106658 130588 106966 130597
rect 106658 130586 106664 130588
rect 106720 130586 106744 130588
rect 106800 130586 106824 130588
rect 106880 130586 106904 130588
rect 106960 130586 106966 130588
rect 106720 130534 106722 130586
rect 106902 130534 106904 130586
rect 106658 130532 106664 130534
rect 106720 130532 106744 130534
rect 106800 130532 106824 130534
rect 106880 130532 106904 130534
rect 106960 130532 106966 130534
rect 106658 130523 106966 130532
rect 105922 130044 106230 130053
rect 105922 130042 105928 130044
rect 105984 130042 106008 130044
rect 106064 130042 106088 130044
rect 106144 130042 106168 130044
rect 106224 130042 106230 130044
rect 105984 129990 105986 130042
rect 106166 129990 106168 130042
rect 105922 129988 105928 129990
rect 105984 129988 106008 129990
rect 106064 129988 106088 129990
rect 106144 129988 106168 129990
rect 106224 129988 106230 129990
rect 105922 129979 106230 129988
rect 104348 129872 104400 129878
rect 104346 129840 104348 129849
rect 104400 129840 104402 129849
rect 104346 129775 104402 129784
rect 106658 129500 106966 129509
rect 106658 129498 106664 129500
rect 106720 129498 106744 129500
rect 106800 129498 106824 129500
rect 106880 129498 106904 129500
rect 106960 129498 106966 129500
rect 106720 129446 106722 129498
rect 106902 129446 106904 129498
rect 106658 129444 106664 129446
rect 106720 129444 106744 129446
rect 106800 129444 106824 129446
rect 106880 129444 106904 129446
rect 106960 129444 106966 129446
rect 106658 129435 106966 129444
rect 105922 128956 106230 128965
rect 105922 128954 105928 128956
rect 105984 128954 106008 128956
rect 106064 128954 106088 128956
rect 106144 128954 106168 128956
rect 106224 128954 106230 128956
rect 105984 128902 105986 128954
rect 106166 128902 106168 128954
rect 105922 128900 105928 128902
rect 105984 128900 106008 128902
rect 106064 128900 106088 128902
rect 106144 128900 106168 128902
rect 106224 128900 106230 128902
rect 105922 128891 106230 128900
rect 106658 128412 106966 128421
rect 106658 128410 106664 128412
rect 106720 128410 106744 128412
rect 106800 128410 106824 128412
rect 106880 128410 106904 128412
rect 106960 128410 106966 128412
rect 106720 128358 106722 128410
rect 106902 128358 106904 128410
rect 106658 128356 106664 128358
rect 106720 128356 106744 128358
rect 106800 128356 106824 128358
rect 106880 128356 106904 128358
rect 106960 128356 106966 128358
rect 106658 128347 106966 128356
rect 105922 127868 106230 127877
rect 105922 127866 105928 127868
rect 105984 127866 106008 127868
rect 106064 127866 106088 127868
rect 106144 127866 106168 127868
rect 106224 127866 106230 127868
rect 105984 127814 105986 127866
rect 106166 127814 106168 127866
rect 105922 127812 105928 127814
rect 105984 127812 106008 127814
rect 106064 127812 106088 127814
rect 106144 127812 106168 127814
rect 106224 127812 106230 127814
rect 105922 127803 106230 127812
rect 106658 127324 106966 127333
rect 106658 127322 106664 127324
rect 106720 127322 106744 127324
rect 106800 127322 106824 127324
rect 106880 127322 106904 127324
rect 106960 127322 106966 127324
rect 106720 127270 106722 127322
rect 106902 127270 106904 127322
rect 106658 127268 106664 127270
rect 106720 127268 106744 127270
rect 106800 127268 106824 127270
rect 106880 127268 106904 127270
rect 106960 127268 106966 127270
rect 106658 127259 106966 127268
rect 105922 126780 106230 126789
rect 105922 126778 105928 126780
rect 105984 126778 106008 126780
rect 106064 126778 106088 126780
rect 106144 126778 106168 126780
rect 106224 126778 106230 126780
rect 105984 126726 105986 126778
rect 106166 126726 106168 126778
rect 105922 126724 105928 126726
rect 105984 126724 106008 126726
rect 106064 126724 106088 126726
rect 106144 126724 106168 126726
rect 106224 126724 106230 126726
rect 105922 126715 106230 126724
rect 106658 126236 106966 126245
rect 106658 126234 106664 126236
rect 106720 126234 106744 126236
rect 106800 126234 106824 126236
rect 106880 126234 106904 126236
rect 106960 126234 106966 126236
rect 106720 126182 106722 126234
rect 106902 126182 106904 126234
rect 106658 126180 106664 126182
rect 106720 126180 106744 126182
rect 106800 126180 106824 126182
rect 106880 126180 106904 126182
rect 106960 126180 106966 126182
rect 106658 126171 106966 126180
rect 105922 125692 106230 125701
rect 105922 125690 105928 125692
rect 105984 125690 106008 125692
rect 106064 125690 106088 125692
rect 106144 125690 106168 125692
rect 106224 125690 106230 125692
rect 105984 125638 105986 125690
rect 106166 125638 106168 125690
rect 105922 125636 105928 125638
rect 105984 125636 106008 125638
rect 106064 125636 106088 125638
rect 106144 125636 106168 125638
rect 106224 125636 106230 125638
rect 105922 125627 106230 125636
rect 106658 125148 106966 125157
rect 106658 125146 106664 125148
rect 106720 125146 106744 125148
rect 106800 125146 106824 125148
rect 106880 125146 106904 125148
rect 106960 125146 106966 125148
rect 106720 125094 106722 125146
rect 106902 125094 106904 125146
rect 106658 125092 106664 125094
rect 106720 125092 106744 125094
rect 106800 125092 106824 125094
rect 106880 125092 106904 125094
rect 106960 125092 106966 125094
rect 106658 125083 106966 125092
rect 105922 124604 106230 124613
rect 105922 124602 105928 124604
rect 105984 124602 106008 124604
rect 106064 124602 106088 124604
rect 106144 124602 106168 124604
rect 106224 124602 106230 124604
rect 105984 124550 105986 124602
rect 106166 124550 106168 124602
rect 105922 124548 105928 124550
rect 105984 124548 106008 124550
rect 106064 124548 106088 124550
rect 106144 124548 106168 124550
rect 106224 124548 106230 124550
rect 105922 124539 106230 124548
rect 106658 124060 106966 124069
rect 106658 124058 106664 124060
rect 106720 124058 106744 124060
rect 106800 124058 106824 124060
rect 106880 124058 106904 124060
rect 106960 124058 106966 124060
rect 106720 124006 106722 124058
rect 106902 124006 106904 124058
rect 106658 124004 106664 124006
rect 106720 124004 106744 124006
rect 106800 124004 106824 124006
rect 106880 124004 106904 124006
rect 106960 124004 106966 124006
rect 106658 123995 106966 124004
rect 105922 123516 106230 123525
rect 105922 123514 105928 123516
rect 105984 123514 106008 123516
rect 106064 123514 106088 123516
rect 106144 123514 106168 123516
rect 106224 123514 106230 123516
rect 105984 123462 105986 123514
rect 106166 123462 106168 123514
rect 105922 123460 105928 123462
rect 105984 123460 106008 123462
rect 106064 123460 106088 123462
rect 106144 123460 106168 123462
rect 106224 123460 106230 123462
rect 105922 123451 106230 123460
rect 106658 122972 106966 122981
rect 106658 122970 106664 122972
rect 106720 122970 106744 122972
rect 106800 122970 106824 122972
rect 106880 122970 106904 122972
rect 106960 122970 106966 122972
rect 106720 122918 106722 122970
rect 106902 122918 106904 122970
rect 106658 122916 106664 122918
rect 106720 122916 106744 122918
rect 106800 122916 106824 122918
rect 106880 122916 106904 122918
rect 106960 122916 106966 122918
rect 106658 122907 106966 122916
rect 105922 122428 106230 122437
rect 105922 122426 105928 122428
rect 105984 122426 106008 122428
rect 106064 122426 106088 122428
rect 106144 122426 106168 122428
rect 106224 122426 106230 122428
rect 105984 122374 105986 122426
rect 106166 122374 106168 122426
rect 105922 122372 105928 122374
rect 105984 122372 106008 122374
rect 106064 122372 106088 122374
rect 106144 122372 106168 122374
rect 106224 122372 106230 122374
rect 105922 122363 106230 122372
rect 106658 121884 106966 121893
rect 106658 121882 106664 121884
rect 106720 121882 106744 121884
rect 106800 121882 106824 121884
rect 106880 121882 106904 121884
rect 106960 121882 106966 121884
rect 106720 121830 106722 121882
rect 106902 121830 106904 121882
rect 106658 121828 106664 121830
rect 106720 121828 106744 121830
rect 106800 121828 106824 121830
rect 106880 121828 106904 121830
rect 106960 121828 106966 121830
rect 106658 121819 106966 121828
rect 105922 121340 106230 121349
rect 105922 121338 105928 121340
rect 105984 121338 106008 121340
rect 106064 121338 106088 121340
rect 106144 121338 106168 121340
rect 106224 121338 106230 121340
rect 105984 121286 105986 121338
rect 106166 121286 106168 121338
rect 105922 121284 105928 121286
rect 105984 121284 106008 121286
rect 106064 121284 106088 121286
rect 106144 121284 106168 121286
rect 106224 121284 106230 121286
rect 105922 121275 106230 121284
rect 106658 120796 106966 120805
rect 106658 120794 106664 120796
rect 106720 120794 106744 120796
rect 106800 120794 106824 120796
rect 106880 120794 106904 120796
rect 106960 120794 106966 120796
rect 106720 120742 106722 120794
rect 106902 120742 106904 120794
rect 106658 120740 106664 120742
rect 106720 120740 106744 120742
rect 106800 120740 106824 120742
rect 106880 120740 106904 120742
rect 106960 120740 106966 120742
rect 106658 120731 106966 120740
rect 105922 120252 106230 120261
rect 105922 120250 105928 120252
rect 105984 120250 106008 120252
rect 106064 120250 106088 120252
rect 106144 120250 106168 120252
rect 106224 120250 106230 120252
rect 105984 120198 105986 120250
rect 106166 120198 106168 120250
rect 105922 120196 105928 120198
rect 105984 120196 106008 120198
rect 106064 120196 106088 120198
rect 106144 120196 106168 120198
rect 106224 120196 106230 120198
rect 105922 120187 106230 120196
rect 106658 119708 106966 119717
rect 106658 119706 106664 119708
rect 106720 119706 106744 119708
rect 106800 119706 106824 119708
rect 106880 119706 106904 119708
rect 106960 119706 106966 119708
rect 106720 119654 106722 119706
rect 106902 119654 106904 119706
rect 106658 119652 106664 119654
rect 106720 119652 106744 119654
rect 106800 119652 106824 119654
rect 106880 119652 106904 119654
rect 106960 119652 106966 119654
rect 106658 119643 106966 119652
rect 105922 119164 106230 119173
rect 105922 119162 105928 119164
rect 105984 119162 106008 119164
rect 106064 119162 106088 119164
rect 106144 119162 106168 119164
rect 106224 119162 106230 119164
rect 105984 119110 105986 119162
rect 106166 119110 106168 119162
rect 105922 119108 105928 119110
rect 105984 119108 106008 119110
rect 106064 119108 106088 119110
rect 106144 119108 106168 119110
rect 106224 119108 106230 119110
rect 105922 119099 106230 119108
rect 106658 118620 106966 118629
rect 106658 118618 106664 118620
rect 106720 118618 106744 118620
rect 106800 118618 106824 118620
rect 106880 118618 106904 118620
rect 106960 118618 106966 118620
rect 106720 118566 106722 118618
rect 106902 118566 106904 118618
rect 106658 118564 106664 118566
rect 106720 118564 106744 118566
rect 106800 118564 106824 118566
rect 106880 118564 106904 118566
rect 106960 118564 106966 118566
rect 106658 118555 106966 118564
rect 105922 118076 106230 118085
rect 105922 118074 105928 118076
rect 105984 118074 106008 118076
rect 106064 118074 106088 118076
rect 106144 118074 106168 118076
rect 106224 118074 106230 118076
rect 105984 118022 105986 118074
rect 106166 118022 106168 118074
rect 105922 118020 105928 118022
rect 105984 118020 106008 118022
rect 106064 118020 106088 118022
rect 106144 118020 106168 118022
rect 106224 118020 106230 118022
rect 105922 118011 106230 118020
rect 106658 117532 106966 117541
rect 106658 117530 106664 117532
rect 106720 117530 106744 117532
rect 106800 117530 106824 117532
rect 106880 117530 106904 117532
rect 106960 117530 106966 117532
rect 106720 117478 106722 117530
rect 106902 117478 106904 117530
rect 106658 117476 106664 117478
rect 106720 117476 106744 117478
rect 106800 117476 106824 117478
rect 106880 117476 106904 117478
rect 106960 117476 106966 117478
rect 106658 117467 106966 117476
rect 105922 116988 106230 116997
rect 105922 116986 105928 116988
rect 105984 116986 106008 116988
rect 106064 116986 106088 116988
rect 106144 116986 106168 116988
rect 106224 116986 106230 116988
rect 105984 116934 105986 116986
rect 106166 116934 106168 116986
rect 105922 116932 105928 116934
rect 105984 116932 106008 116934
rect 106064 116932 106088 116934
rect 106144 116932 106168 116934
rect 106224 116932 106230 116934
rect 105922 116923 106230 116932
rect 106658 116444 106966 116453
rect 106658 116442 106664 116444
rect 106720 116442 106744 116444
rect 106800 116442 106824 116444
rect 106880 116442 106904 116444
rect 106960 116442 106966 116444
rect 106720 116390 106722 116442
rect 106902 116390 106904 116442
rect 106658 116388 106664 116390
rect 106720 116388 106744 116390
rect 106800 116388 106824 116390
rect 106880 116388 106904 116390
rect 106960 116388 106966 116390
rect 106658 116379 106966 116388
rect 105922 115900 106230 115909
rect 105922 115898 105928 115900
rect 105984 115898 106008 115900
rect 106064 115898 106088 115900
rect 106144 115898 106168 115900
rect 106224 115898 106230 115900
rect 105984 115846 105986 115898
rect 106166 115846 106168 115898
rect 105922 115844 105928 115846
rect 105984 115844 106008 115846
rect 106064 115844 106088 115846
rect 106144 115844 106168 115846
rect 106224 115844 106230 115846
rect 105922 115835 106230 115844
rect 106658 115356 106966 115365
rect 106658 115354 106664 115356
rect 106720 115354 106744 115356
rect 106800 115354 106824 115356
rect 106880 115354 106904 115356
rect 106960 115354 106966 115356
rect 106720 115302 106722 115354
rect 106902 115302 106904 115354
rect 106658 115300 106664 115302
rect 106720 115300 106744 115302
rect 106800 115300 106824 115302
rect 106880 115300 106904 115302
rect 106960 115300 106966 115302
rect 106658 115291 106966 115300
rect 105922 114812 106230 114821
rect 105922 114810 105928 114812
rect 105984 114810 106008 114812
rect 106064 114810 106088 114812
rect 106144 114810 106168 114812
rect 106224 114810 106230 114812
rect 105984 114758 105986 114810
rect 106166 114758 106168 114810
rect 105922 114756 105928 114758
rect 105984 114756 106008 114758
rect 106064 114756 106088 114758
rect 106144 114756 106168 114758
rect 106224 114756 106230 114758
rect 105922 114747 106230 114756
rect 106658 114268 106966 114277
rect 106658 114266 106664 114268
rect 106720 114266 106744 114268
rect 106800 114266 106824 114268
rect 106880 114266 106904 114268
rect 106960 114266 106966 114268
rect 106720 114214 106722 114266
rect 106902 114214 106904 114266
rect 106658 114212 106664 114214
rect 106720 114212 106744 114214
rect 106800 114212 106824 114214
rect 106880 114212 106904 114214
rect 106960 114212 106966 114214
rect 106658 114203 106966 114212
rect 105922 113724 106230 113733
rect 105922 113722 105928 113724
rect 105984 113722 106008 113724
rect 106064 113722 106088 113724
rect 106144 113722 106168 113724
rect 106224 113722 106230 113724
rect 105984 113670 105986 113722
rect 106166 113670 106168 113722
rect 105922 113668 105928 113670
rect 105984 113668 106008 113670
rect 106064 113668 106088 113670
rect 106144 113668 106168 113670
rect 106224 113668 106230 113670
rect 105922 113659 106230 113668
rect 106658 113180 106966 113189
rect 106658 113178 106664 113180
rect 106720 113178 106744 113180
rect 106800 113178 106824 113180
rect 106880 113178 106904 113180
rect 106960 113178 106966 113180
rect 106720 113126 106722 113178
rect 106902 113126 106904 113178
rect 106658 113124 106664 113126
rect 106720 113124 106744 113126
rect 106800 113124 106824 113126
rect 106880 113124 106904 113126
rect 106960 113124 106966 113126
rect 106658 113115 106966 113124
rect 105922 112636 106230 112645
rect 105922 112634 105928 112636
rect 105984 112634 106008 112636
rect 106064 112634 106088 112636
rect 106144 112634 106168 112636
rect 106224 112634 106230 112636
rect 105984 112582 105986 112634
rect 106166 112582 106168 112634
rect 105922 112580 105928 112582
rect 105984 112580 106008 112582
rect 106064 112580 106088 112582
rect 106144 112580 106168 112582
rect 106224 112580 106230 112582
rect 105922 112571 106230 112580
rect 106658 112092 106966 112101
rect 106658 112090 106664 112092
rect 106720 112090 106744 112092
rect 106800 112090 106824 112092
rect 106880 112090 106904 112092
rect 106960 112090 106966 112092
rect 106720 112038 106722 112090
rect 106902 112038 106904 112090
rect 106658 112036 106664 112038
rect 106720 112036 106744 112038
rect 106800 112036 106824 112038
rect 106880 112036 106904 112038
rect 106960 112036 106966 112038
rect 106658 112027 106966 112036
rect 105922 111548 106230 111557
rect 105922 111546 105928 111548
rect 105984 111546 106008 111548
rect 106064 111546 106088 111548
rect 106144 111546 106168 111548
rect 106224 111546 106230 111548
rect 105984 111494 105986 111546
rect 106166 111494 106168 111546
rect 105922 111492 105928 111494
rect 105984 111492 106008 111494
rect 106064 111492 106088 111494
rect 106144 111492 106168 111494
rect 106224 111492 106230 111494
rect 105922 111483 106230 111492
rect 106658 111004 106966 111013
rect 106658 111002 106664 111004
rect 106720 111002 106744 111004
rect 106800 111002 106824 111004
rect 106880 111002 106904 111004
rect 106960 111002 106966 111004
rect 106720 110950 106722 111002
rect 106902 110950 106904 111002
rect 106658 110948 106664 110950
rect 106720 110948 106744 110950
rect 106800 110948 106824 110950
rect 106880 110948 106904 110950
rect 106960 110948 106966 110950
rect 106658 110939 106966 110948
rect 105922 110460 106230 110469
rect 105922 110458 105928 110460
rect 105984 110458 106008 110460
rect 106064 110458 106088 110460
rect 106144 110458 106168 110460
rect 106224 110458 106230 110460
rect 105984 110406 105986 110458
rect 106166 110406 106168 110458
rect 105922 110404 105928 110406
rect 105984 110404 106008 110406
rect 106064 110404 106088 110406
rect 106144 110404 106168 110406
rect 106224 110404 106230 110406
rect 105922 110395 106230 110404
rect 106658 109916 106966 109925
rect 106658 109914 106664 109916
rect 106720 109914 106744 109916
rect 106800 109914 106824 109916
rect 106880 109914 106904 109916
rect 106960 109914 106966 109916
rect 106720 109862 106722 109914
rect 106902 109862 106904 109914
rect 106658 109860 106664 109862
rect 106720 109860 106744 109862
rect 106800 109860 106824 109862
rect 106880 109860 106904 109862
rect 106960 109860 106966 109862
rect 106658 109851 106966 109860
rect 105922 109372 106230 109381
rect 105922 109370 105928 109372
rect 105984 109370 106008 109372
rect 106064 109370 106088 109372
rect 106144 109370 106168 109372
rect 106224 109370 106230 109372
rect 105984 109318 105986 109370
rect 106166 109318 106168 109370
rect 105922 109316 105928 109318
rect 105984 109316 106008 109318
rect 106064 109316 106088 109318
rect 106144 109316 106168 109318
rect 106224 109316 106230 109318
rect 105922 109307 106230 109316
rect 106658 108828 106966 108837
rect 106658 108826 106664 108828
rect 106720 108826 106744 108828
rect 106800 108826 106824 108828
rect 106880 108826 106904 108828
rect 106960 108826 106966 108828
rect 106720 108774 106722 108826
rect 106902 108774 106904 108826
rect 106658 108772 106664 108774
rect 106720 108772 106744 108774
rect 106800 108772 106824 108774
rect 106880 108772 106904 108774
rect 106960 108772 106966 108774
rect 106658 108763 106966 108772
rect 105922 108284 106230 108293
rect 105922 108282 105928 108284
rect 105984 108282 106008 108284
rect 106064 108282 106088 108284
rect 106144 108282 106168 108284
rect 106224 108282 106230 108284
rect 105984 108230 105986 108282
rect 106166 108230 106168 108282
rect 105922 108228 105928 108230
rect 105984 108228 106008 108230
rect 106064 108228 106088 108230
rect 106144 108228 106168 108230
rect 106224 108228 106230 108230
rect 105922 108219 106230 108228
rect 106658 107740 106966 107749
rect 106658 107738 106664 107740
rect 106720 107738 106744 107740
rect 106800 107738 106824 107740
rect 106880 107738 106904 107740
rect 106960 107738 106966 107740
rect 106720 107686 106722 107738
rect 106902 107686 106904 107738
rect 106658 107684 106664 107686
rect 106720 107684 106744 107686
rect 106800 107684 106824 107686
rect 106880 107684 106904 107686
rect 106960 107684 106966 107686
rect 106658 107675 106966 107684
rect 105922 107196 106230 107205
rect 105922 107194 105928 107196
rect 105984 107194 106008 107196
rect 106064 107194 106088 107196
rect 106144 107194 106168 107196
rect 106224 107194 106230 107196
rect 105984 107142 105986 107194
rect 106166 107142 106168 107194
rect 105922 107140 105928 107142
rect 105984 107140 106008 107142
rect 106064 107140 106088 107142
rect 106144 107140 106168 107142
rect 106224 107140 106230 107142
rect 105922 107131 106230 107140
rect 106658 106652 106966 106661
rect 106658 106650 106664 106652
rect 106720 106650 106744 106652
rect 106800 106650 106824 106652
rect 106880 106650 106904 106652
rect 106960 106650 106966 106652
rect 106720 106598 106722 106650
rect 106902 106598 106904 106650
rect 106658 106596 106664 106598
rect 106720 106596 106744 106598
rect 106800 106596 106824 106598
rect 106880 106596 106904 106598
rect 106960 106596 106966 106598
rect 106658 106587 106966 106596
rect 105922 106108 106230 106117
rect 105922 106106 105928 106108
rect 105984 106106 106008 106108
rect 106064 106106 106088 106108
rect 106144 106106 106168 106108
rect 106224 106106 106230 106108
rect 105984 106054 105986 106106
rect 106166 106054 106168 106106
rect 105922 106052 105928 106054
rect 105984 106052 106008 106054
rect 106064 106052 106088 106054
rect 106144 106052 106168 106054
rect 106224 106052 106230 106054
rect 105922 106043 106230 106052
rect 106658 105564 106966 105573
rect 106658 105562 106664 105564
rect 106720 105562 106744 105564
rect 106800 105562 106824 105564
rect 106880 105562 106904 105564
rect 106960 105562 106966 105564
rect 106720 105510 106722 105562
rect 106902 105510 106904 105562
rect 106658 105508 106664 105510
rect 106720 105508 106744 105510
rect 106800 105508 106824 105510
rect 106880 105508 106904 105510
rect 106960 105508 106966 105510
rect 106658 105499 106966 105508
rect 105922 105020 106230 105029
rect 105922 105018 105928 105020
rect 105984 105018 106008 105020
rect 106064 105018 106088 105020
rect 106144 105018 106168 105020
rect 106224 105018 106230 105020
rect 105984 104966 105986 105018
rect 106166 104966 106168 105018
rect 105922 104964 105928 104966
rect 105984 104964 106008 104966
rect 106064 104964 106088 104966
rect 106144 104964 106168 104966
rect 106224 104964 106230 104966
rect 105922 104955 106230 104964
rect 106658 104476 106966 104485
rect 106658 104474 106664 104476
rect 106720 104474 106744 104476
rect 106800 104474 106824 104476
rect 106880 104474 106904 104476
rect 106960 104474 106966 104476
rect 106720 104422 106722 104474
rect 106902 104422 106904 104474
rect 106658 104420 106664 104422
rect 106720 104420 106744 104422
rect 106800 104420 106824 104422
rect 106880 104420 106904 104422
rect 106960 104420 106966 104422
rect 106658 104411 106966 104420
rect 105922 103932 106230 103941
rect 105922 103930 105928 103932
rect 105984 103930 106008 103932
rect 106064 103930 106088 103932
rect 106144 103930 106168 103932
rect 106224 103930 106230 103932
rect 105984 103878 105986 103930
rect 106166 103878 106168 103930
rect 105922 103876 105928 103878
rect 105984 103876 106008 103878
rect 106064 103876 106088 103878
rect 106144 103876 106168 103878
rect 106224 103876 106230 103878
rect 105922 103867 106230 103876
rect 106658 103388 106966 103397
rect 106658 103386 106664 103388
rect 106720 103386 106744 103388
rect 106800 103386 106824 103388
rect 106880 103386 106904 103388
rect 106960 103386 106966 103388
rect 106720 103334 106722 103386
rect 106902 103334 106904 103386
rect 106658 103332 106664 103334
rect 106720 103332 106744 103334
rect 106800 103332 106824 103334
rect 106880 103332 106904 103334
rect 106960 103332 106966 103334
rect 106658 103323 106966 103332
rect 105922 102844 106230 102853
rect 105922 102842 105928 102844
rect 105984 102842 106008 102844
rect 106064 102842 106088 102844
rect 106144 102842 106168 102844
rect 106224 102842 106230 102844
rect 105984 102790 105986 102842
rect 106166 102790 106168 102842
rect 105922 102788 105928 102790
rect 105984 102788 106008 102790
rect 106064 102788 106088 102790
rect 106144 102788 106168 102790
rect 106224 102788 106230 102790
rect 105922 102779 106230 102788
rect 106658 102300 106966 102309
rect 106658 102298 106664 102300
rect 106720 102298 106744 102300
rect 106800 102298 106824 102300
rect 106880 102298 106904 102300
rect 106960 102298 106966 102300
rect 106720 102246 106722 102298
rect 106902 102246 106904 102298
rect 106658 102244 106664 102246
rect 106720 102244 106744 102246
rect 106800 102244 106824 102246
rect 106880 102244 106904 102246
rect 106960 102244 106966 102246
rect 106658 102235 106966 102244
rect 105922 101756 106230 101765
rect 105922 101754 105928 101756
rect 105984 101754 106008 101756
rect 106064 101754 106088 101756
rect 106144 101754 106168 101756
rect 106224 101754 106230 101756
rect 105984 101702 105986 101754
rect 106166 101702 106168 101754
rect 105922 101700 105928 101702
rect 105984 101700 106008 101702
rect 106064 101700 106088 101702
rect 106144 101700 106168 101702
rect 106224 101700 106230 101702
rect 105922 101691 106230 101700
rect 106658 101212 106966 101221
rect 106658 101210 106664 101212
rect 106720 101210 106744 101212
rect 106800 101210 106824 101212
rect 106880 101210 106904 101212
rect 106960 101210 106966 101212
rect 106720 101158 106722 101210
rect 106902 101158 106904 101210
rect 106658 101156 106664 101158
rect 106720 101156 106744 101158
rect 106800 101156 106824 101158
rect 106880 101156 106904 101158
rect 106960 101156 106966 101158
rect 106658 101147 106966 101156
rect 105922 100668 106230 100677
rect 105922 100666 105928 100668
rect 105984 100666 106008 100668
rect 106064 100666 106088 100668
rect 106144 100666 106168 100668
rect 106224 100666 106230 100668
rect 105984 100614 105986 100666
rect 106166 100614 106168 100666
rect 105922 100612 105928 100614
rect 105984 100612 106008 100614
rect 106064 100612 106088 100614
rect 106144 100612 106168 100614
rect 106224 100612 106230 100614
rect 105922 100603 106230 100612
rect 106658 100124 106966 100133
rect 106658 100122 106664 100124
rect 106720 100122 106744 100124
rect 106800 100122 106824 100124
rect 106880 100122 106904 100124
rect 106960 100122 106966 100124
rect 106720 100070 106722 100122
rect 106902 100070 106904 100122
rect 106658 100068 106664 100070
rect 106720 100068 106744 100070
rect 106800 100068 106824 100070
rect 106880 100068 106904 100070
rect 106960 100068 106966 100070
rect 106658 100059 106966 100068
rect 105922 99580 106230 99589
rect 105922 99578 105928 99580
rect 105984 99578 106008 99580
rect 106064 99578 106088 99580
rect 106144 99578 106168 99580
rect 106224 99578 106230 99580
rect 105984 99526 105986 99578
rect 106166 99526 106168 99578
rect 105922 99524 105928 99526
rect 105984 99524 106008 99526
rect 106064 99524 106088 99526
rect 106144 99524 106168 99526
rect 106224 99524 106230 99526
rect 105922 99515 106230 99524
rect 106658 99036 106966 99045
rect 106658 99034 106664 99036
rect 106720 99034 106744 99036
rect 106800 99034 106824 99036
rect 106880 99034 106904 99036
rect 106960 99034 106966 99036
rect 106720 98982 106722 99034
rect 106902 98982 106904 99034
rect 106658 98980 106664 98982
rect 106720 98980 106744 98982
rect 106800 98980 106824 98982
rect 106880 98980 106904 98982
rect 106960 98980 106966 98982
rect 106658 98971 106966 98980
rect 105922 98492 106230 98501
rect 105922 98490 105928 98492
rect 105984 98490 106008 98492
rect 106064 98490 106088 98492
rect 106144 98490 106168 98492
rect 106224 98490 106230 98492
rect 105984 98438 105986 98490
rect 106166 98438 106168 98490
rect 105922 98436 105928 98438
rect 105984 98436 106008 98438
rect 106064 98436 106088 98438
rect 106144 98436 106168 98438
rect 106224 98436 106230 98438
rect 105922 98427 106230 98436
rect 106658 97948 106966 97957
rect 106658 97946 106664 97948
rect 106720 97946 106744 97948
rect 106800 97946 106824 97948
rect 106880 97946 106904 97948
rect 106960 97946 106966 97948
rect 106720 97894 106722 97946
rect 106902 97894 106904 97946
rect 106658 97892 106664 97894
rect 106720 97892 106744 97894
rect 106800 97892 106824 97894
rect 106880 97892 106904 97894
rect 106960 97892 106966 97894
rect 106658 97883 106966 97892
rect 105922 97404 106230 97413
rect 105922 97402 105928 97404
rect 105984 97402 106008 97404
rect 106064 97402 106088 97404
rect 106144 97402 106168 97404
rect 106224 97402 106230 97404
rect 105984 97350 105986 97402
rect 106166 97350 106168 97402
rect 105922 97348 105928 97350
rect 105984 97348 106008 97350
rect 106064 97348 106088 97350
rect 106144 97348 106168 97350
rect 106224 97348 106230 97350
rect 105922 97339 106230 97348
rect 106658 96860 106966 96869
rect 106658 96858 106664 96860
rect 106720 96858 106744 96860
rect 106800 96858 106824 96860
rect 106880 96858 106904 96860
rect 106960 96858 106966 96860
rect 106720 96806 106722 96858
rect 106902 96806 106904 96858
rect 106658 96804 106664 96806
rect 106720 96804 106744 96806
rect 106800 96804 106824 96806
rect 106880 96804 106904 96806
rect 106960 96804 106966 96806
rect 106658 96795 106966 96804
rect 105922 96316 106230 96325
rect 105922 96314 105928 96316
rect 105984 96314 106008 96316
rect 106064 96314 106088 96316
rect 106144 96314 106168 96316
rect 106224 96314 106230 96316
rect 105984 96262 105986 96314
rect 106166 96262 106168 96314
rect 105922 96260 105928 96262
rect 105984 96260 106008 96262
rect 106064 96260 106088 96262
rect 106144 96260 106168 96262
rect 106224 96260 106230 96262
rect 105922 96251 106230 96260
rect 106658 95772 106966 95781
rect 106658 95770 106664 95772
rect 106720 95770 106744 95772
rect 106800 95770 106824 95772
rect 106880 95770 106904 95772
rect 106960 95770 106966 95772
rect 106720 95718 106722 95770
rect 106902 95718 106904 95770
rect 106658 95716 106664 95718
rect 106720 95716 106744 95718
rect 106800 95716 106824 95718
rect 106880 95716 106904 95718
rect 106960 95716 106966 95718
rect 106658 95707 106966 95716
rect 105922 95228 106230 95237
rect 105922 95226 105928 95228
rect 105984 95226 106008 95228
rect 106064 95226 106088 95228
rect 106144 95226 106168 95228
rect 106224 95226 106230 95228
rect 105984 95174 105986 95226
rect 106166 95174 106168 95226
rect 105922 95172 105928 95174
rect 105984 95172 106008 95174
rect 106064 95172 106088 95174
rect 106144 95172 106168 95174
rect 106224 95172 106230 95174
rect 105922 95163 106230 95172
rect 106658 94684 106966 94693
rect 106658 94682 106664 94684
rect 106720 94682 106744 94684
rect 106800 94682 106824 94684
rect 106880 94682 106904 94684
rect 106960 94682 106966 94684
rect 106720 94630 106722 94682
rect 106902 94630 106904 94682
rect 106658 94628 106664 94630
rect 106720 94628 106744 94630
rect 106800 94628 106824 94630
rect 106880 94628 106904 94630
rect 106960 94628 106966 94630
rect 106658 94619 106966 94628
rect 105922 94140 106230 94149
rect 105922 94138 105928 94140
rect 105984 94138 106008 94140
rect 106064 94138 106088 94140
rect 106144 94138 106168 94140
rect 106224 94138 106230 94140
rect 105984 94086 105986 94138
rect 106166 94086 106168 94138
rect 105922 94084 105928 94086
rect 105984 94084 106008 94086
rect 106064 94084 106088 94086
rect 106144 94084 106168 94086
rect 106224 94084 106230 94086
rect 105922 94075 106230 94084
rect 106658 93596 106966 93605
rect 106658 93594 106664 93596
rect 106720 93594 106744 93596
rect 106800 93594 106824 93596
rect 106880 93594 106904 93596
rect 106960 93594 106966 93596
rect 106720 93542 106722 93594
rect 106902 93542 106904 93594
rect 106658 93540 106664 93542
rect 106720 93540 106744 93542
rect 106800 93540 106824 93542
rect 106880 93540 106904 93542
rect 106960 93540 106966 93542
rect 106658 93531 106966 93540
rect 105922 93052 106230 93061
rect 105922 93050 105928 93052
rect 105984 93050 106008 93052
rect 106064 93050 106088 93052
rect 106144 93050 106168 93052
rect 106224 93050 106230 93052
rect 105984 92998 105986 93050
rect 106166 92998 106168 93050
rect 105922 92996 105928 92998
rect 105984 92996 106008 92998
rect 106064 92996 106088 92998
rect 106144 92996 106168 92998
rect 106224 92996 106230 92998
rect 105922 92987 106230 92996
rect 106658 92508 106966 92517
rect 106658 92506 106664 92508
rect 106720 92506 106744 92508
rect 106800 92506 106824 92508
rect 106880 92506 106904 92508
rect 106960 92506 106966 92508
rect 106720 92454 106722 92506
rect 106902 92454 106904 92506
rect 106658 92452 106664 92454
rect 106720 92452 106744 92454
rect 106800 92452 106824 92454
rect 106880 92452 106904 92454
rect 106960 92452 106966 92454
rect 106658 92443 106966 92452
rect 105922 91964 106230 91973
rect 105922 91962 105928 91964
rect 105984 91962 106008 91964
rect 106064 91962 106088 91964
rect 106144 91962 106168 91964
rect 106224 91962 106230 91964
rect 105984 91910 105986 91962
rect 106166 91910 106168 91962
rect 105922 91908 105928 91910
rect 105984 91908 106008 91910
rect 106064 91908 106088 91910
rect 106144 91908 106168 91910
rect 106224 91908 106230 91910
rect 105922 91899 106230 91908
rect 106658 91420 106966 91429
rect 106658 91418 106664 91420
rect 106720 91418 106744 91420
rect 106800 91418 106824 91420
rect 106880 91418 106904 91420
rect 106960 91418 106966 91420
rect 106720 91366 106722 91418
rect 106902 91366 106904 91418
rect 106658 91364 106664 91366
rect 106720 91364 106744 91366
rect 106800 91364 106824 91366
rect 106880 91364 106904 91366
rect 106960 91364 106966 91366
rect 106658 91355 106966 91364
rect 104348 91180 104400 91186
rect 104348 91122 104400 91128
rect 104164 90976 104216 90982
rect 104164 90918 104216 90924
rect 103978 77480 104034 77489
rect 103978 77415 104034 77424
rect 104176 77382 104204 90918
rect 104360 90438 104388 91122
rect 105922 90876 106230 90885
rect 105922 90874 105928 90876
rect 105984 90874 106008 90876
rect 106064 90874 106088 90876
rect 106144 90874 106168 90876
rect 106224 90874 106230 90876
rect 105984 90822 105986 90874
rect 106166 90822 106168 90874
rect 105922 90820 105928 90822
rect 105984 90820 106008 90822
rect 106064 90820 106088 90822
rect 106144 90820 106168 90822
rect 106224 90820 106230 90822
rect 105922 90811 106230 90820
rect 104348 90432 104400 90438
rect 104348 90374 104400 90380
rect 104164 77376 104216 77382
rect 104164 77318 104216 77324
rect 104360 72486 104388 90374
rect 106658 90332 106966 90341
rect 106658 90330 106664 90332
rect 106720 90330 106744 90332
rect 106800 90330 106824 90332
rect 106880 90330 106904 90332
rect 106960 90330 106966 90332
rect 106720 90278 106722 90330
rect 106902 90278 106904 90330
rect 106658 90276 106664 90278
rect 106720 90276 106744 90278
rect 106800 90276 106824 90278
rect 106880 90276 106904 90278
rect 106960 90276 106966 90278
rect 106658 90267 106966 90276
rect 105922 89788 106230 89797
rect 105922 89786 105928 89788
rect 105984 89786 106008 89788
rect 106064 89786 106088 89788
rect 106144 89786 106168 89788
rect 106224 89786 106230 89788
rect 105984 89734 105986 89786
rect 106166 89734 106168 89786
rect 105922 89732 105928 89734
rect 105984 89732 106008 89734
rect 106064 89732 106088 89734
rect 106144 89732 106168 89734
rect 106224 89732 106230 89734
rect 105922 89723 106230 89732
rect 106658 89244 106966 89253
rect 106658 89242 106664 89244
rect 106720 89242 106744 89244
rect 106800 89242 106824 89244
rect 106880 89242 106904 89244
rect 106960 89242 106966 89244
rect 106720 89190 106722 89242
rect 106902 89190 106904 89242
rect 106658 89188 106664 89190
rect 106720 89188 106744 89190
rect 106800 89188 106824 89190
rect 106880 89188 106904 89190
rect 106960 89188 106966 89190
rect 106658 89179 106966 89188
rect 105922 88700 106230 88709
rect 105922 88698 105928 88700
rect 105984 88698 106008 88700
rect 106064 88698 106088 88700
rect 106144 88698 106168 88700
rect 106224 88698 106230 88700
rect 105984 88646 105986 88698
rect 106166 88646 106168 88698
rect 105922 88644 105928 88646
rect 105984 88644 106008 88646
rect 106064 88644 106088 88646
rect 106144 88644 106168 88646
rect 106224 88644 106230 88646
rect 105922 88635 106230 88644
rect 106658 88156 106966 88165
rect 106658 88154 106664 88156
rect 106720 88154 106744 88156
rect 106800 88154 106824 88156
rect 106880 88154 106904 88156
rect 106960 88154 106966 88156
rect 106720 88102 106722 88154
rect 106902 88102 106904 88154
rect 106658 88100 106664 88102
rect 106720 88100 106744 88102
rect 106800 88100 106824 88102
rect 106880 88100 106904 88102
rect 106960 88100 106966 88102
rect 106658 88091 106966 88100
rect 105922 87612 106230 87621
rect 105922 87610 105928 87612
rect 105984 87610 106008 87612
rect 106064 87610 106088 87612
rect 106144 87610 106168 87612
rect 106224 87610 106230 87612
rect 105984 87558 105986 87610
rect 106166 87558 106168 87610
rect 105922 87556 105928 87558
rect 105984 87556 106008 87558
rect 106064 87556 106088 87558
rect 106144 87556 106168 87558
rect 106224 87556 106230 87558
rect 105922 87547 106230 87556
rect 106658 87068 106966 87077
rect 106658 87066 106664 87068
rect 106720 87066 106744 87068
rect 106800 87066 106824 87068
rect 106880 87066 106904 87068
rect 106960 87066 106966 87068
rect 106720 87014 106722 87066
rect 106902 87014 106904 87066
rect 106658 87012 106664 87014
rect 106720 87012 106744 87014
rect 106800 87012 106824 87014
rect 106880 87012 106904 87014
rect 106960 87012 106966 87014
rect 106658 87003 106966 87012
rect 105922 86524 106230 86533
rect 105922 86522 105928 86524
rect 105984 86522 106008 86524
rect 106064 86522 106088 86524
rect 106144 86522 106168 86524
rect 106224 86522 106230 86524
rect 105984 86470 105986 86522
rect 106166 86470 106168 86522
rect 105922 86468 105928 86470
rect 105984 86468 106008 86470
rect 106064 86468 106088 86470
rect 106144 86468 106168 86470
rect 106224 86468 106230 86470
rect 105922 86459 106230 86468
rect 106658 85980 106966 85989
rect 106658 85978 106664 85980
rect 106720 85978 106744 85980
rect 106800 85978 106824 85980
rect 106880 85978 106904 85980
rect 106960 85978 106966 85980
rect 106720 85926 106722 85978
rect 106902 85926 106904 85978
rect 106658 85924 106664 85926
rect 106720 85924 106744 85926
rect 106800 85924 106824 85926
rect 106880 85924 106904 85926
rect 106960 85924 106966 85926
rect 106658 85915 106966 85924
rect 105922 85436 106230 85445
rect 105922 85434 105928 85436
rect 105984 85434 106008 85436
rect 106064 85434 106088 85436
rect 106144 85434 106168 85436
rect 106224 85434 106230 85436
rect 105984 85382 105986 85434
rect 106166 85382 106168 85434
rect 105922 85380 105928 85382
rect 105984 85380 106008 85382
rect 106064 85380 106088 85382
rect 106144 85380 106168 85382
rect 106224 85380 106230 85382
rect 105922 85371 106230 85380
rect 106658 84892 106966 84901
rect 106658 84890 106664 84892
rect 106720 84890 106744 84892
rect 106800 84890 106824 84892
rect 106880 84890 106904 84892
rect 106960 84890 106966 84892
rect 106720 84838 106722 84890
rect 106902 84838 106904 84890
rect 106658 84836 106664 84838
rect 106720 84836 106744 84838
rect 106800 84836 106824 84838
rect 106880 84836 106904 84838
rect 106960 84836 106966 84838
rect 106658 84827 106966 84836
rect 105922 84348 106230 84357
rect 105922 84346 105928 84348
rect 105984 84346 106008 84348
rect 106064 84346 106088 84348
rect 106144 84346 106168 84348
rect 106224 84346 106230 84348
rect 105984 84294 105986 84346
rect 106166 84294 106168 84346
rect 105922 84292 105928 84294
rect 105984 84292 106008 84294
rect 106064 84292 106088 84294
rect 106144 84292 106168 84294
rect 106224 84292 106230 84294
rect 105922 84283 106230 84292
rect 106658 83804 106966 83813
rect 106658 83802 106664 83804
rect 106720 83802 106744 83804
rect 106800 83802 106824 83804
rect 106880 83802 106904 83804
rect 106960 83802 106966 83804
rect 106720 83750 106722 83802
rect 106902 83750 106904 83802
rect 106658 83748 106664 83750
rect 106720 83748 106744 83750
rect 106800 83748 106824 83750
rect 106880 83748 106904 83750
rect 106960 83748 106966 83750
rect 106658 83739 106966 83748
rect 105922 83260 106230 83269
rect 105922 83258 105928 83260
rect 105984 83258 106008 83260
rect 106064 83258 106088 83260
rect 106144 83258 106168 83260
rect 106224 83258 106230 83260
rect 105984 83206 105986 83258
rect 106166 83206 106168 83258
rect 105922 83204 105928 83206
rect 105984 83204 106008 83206
rect 106064 83204 106088 83206
rect 106144 83204 106168 83206
rect 106224 83204 106230 83206
rect 105922 83195 106230 83204
rect 106658 82716 106966 82725
rect 106658 82714 106664 82716
rect 106720 82714 106744 82716
rect 106800 82714 106824 82716
rect 106880 82714 106904 82716
rect 106960 82714 106966 82716
rect 106720 82662 106722 82714
rect 106902 82662 106904 82714
rect 106658 82660 106664 82662
rect 106720 82660 106744 82662
rect 106800 82660 106824 82662
rect 106880 82660 106904 82662
rect 106960 82660 106966 82662
rect 106658 82651 106966 82660
rect 105922 82172 106230 82181
rect 105922 82170 105928 82172
rect 105984 82170 106008 82172
rect 106064 82170 106088 82172
rect 106144 82170 106168 82172
rect 106224 82170 106230 82172
rect 105984 82118 105986 82170
rect 106166 82118 106168 82170
rect 105922 82116 105928 82118
rect 105984 82116 106008 82118
rect 106064 82116 106088 82118
rect 106144 82116 106168 82118
rect 106224 82116 106230 82118
rect 105922 82107 106230 82116
rect 106658 81628 106966 81637
rect 106658 81626 106664 81628
rect 106720 81626 106744 81628
rect 106800 81626 106824 81628
rect 106880 81626 106904 81628
rect 106960 81626 106966 81628
rect 106720 81574 106722 81626
rect 106902 81574 106904 81626
rect 106658 81572 106664 81574
rect 106720 81572 106744 81574
rect 106800 81572 106824 81574
rect 106880 81572 106904 81574
rect 106960 81572 106966 81574
rect 106658 81563 106966 81572
rect 105922 81084 106230 81093
rect 105922 81082 105928 81084
rect 105984 81082 106008 81084
rect 106064 81082 106088 81084
rect 106144 81082 106168 81084
rect 106224 81082 106230 81084
rect 105984 81030 105986 81082
rect 106166 81030 106168 81082
rect 105922 81028 105928 81030
rect 105984 81028 106008 81030
rect 106064 81028 106088 81030
rect 106144 81028 106168 81030
rect 106224 81028 106230 81030
rect 105922 81019 106230 81028
rect 106658 80540 106966 80549
rect 106658 80538 106664 80540
rect 106720 80538 106744 80540
rect 106800 80538 106824 80540
rect 106880 80538 106904 80540
rect 106960 80538 106966 80540
rect 106720 80486 106722 80538
rect 106902 80486 106904 80538
rect 106658 80484 106664 80486
rect 106720 80484 106744 80486
rect 106800 80484 106824 80486
rect 106880 80484 106904 80486
rect 106960 80484 106966 80486
rect 106658 80475 106966 80484
rect 105922 79996 106230 80005
rect 105922 79994 105928 79996
rect 105984 79994 106008 79996
rect 106064 79994 106088 79996
rect 106144 79994 106168 79996
rect 106224 79994 106230 79996
rect 105984 79942 105986 79994
rect 106166 79942 106168 79994
rect 105922 79940 105928 79942
rect 105984 79940 106008 79942
rect 106064 79940 106088 79942
rect 106144 79940 106168 79942
rect 106224 79940 106230 79942
rect 105922 79931 106230 79940
rect 106658 79452 106966 79461
rect 106658 79450 106664 79452
rect 106720 79450 106744 79452
rect 106800 79450 106824 79452
rect 106880 79450 106904 79452
rect 106960 79450 106966 79452
rect 106720 79398 106722 79450
rect 106902 79398 106904 79450
rect 106658 79396 106664 79398
rect 106720 79396 106744 79398
rect 106800 79396 106824 79398
rect 106880 79396 106904 79398
rect 106960 79396 106966 79398
rect 106658 79387 106966 79396
rect 108488 79008 108540 79014
rect 108486 78976 108488 78985
rect 108540 78976 108542 78985
rect 105922 78908 106230 78917
rect 108486 78911 108542 78920
rect 105922 78906 105928 78908
rect 105984 78906 106008 78908
rect 106064 78906 106088 78908
rect 106144 78906 106168 78908
rect 106224 78906 106230 78908
rect 105984 78854 105986 78906
rect 106166 78854 106168 78906
rect 105922 78852 105928 78854
rect 105984 78852 106008 78854
rect 106064 78852 106088 78854
rect 106144 78852 106168 78854
rect 106224 78852 106230 78854
rect 105922 78843 106230 78852
rect 108120 78464 108172 78470
rect 108120 78406 108172 78412
rect 108488 78464 108540 78470
rect 108488 78406 108540 78412
rect 106658 78364 106966 78373
rect 106658 78362 106664 78364
rect 106720 78362 106744 78364
rect 106800 78362 106824 78364
rect 106880 78362 106904 78364
rect 106960 78362 106966 78364
rect 106720 78310 106722 78362
rect 106902 78310 106904 78362
rect 106658 78308 106664 78310
rect 106720 78308 106744 78310
rect 106800 78308 106824 78310
rect 106880 78308 106904 78310
rect 106960 78308 106966 78310
rect 106658 78299 106966 78308
rect 107660 78056 107712 78062
rect 107660 77998 107712 78004
rect 105820 77920 105872 77926
rect 105820 77862 105872 77868
rect 105832 76906 105860 77862
rect 105922 77820 106230 77829
rect 105922 77818 105928 77820
rect 105984 77818 106008 77820
rect 106064 77818 106088 77820
rect 106144 77818 106168 77820
rect 106224 77818 106230 77820
rect 105984 77766 105986 77818
rect 106166 77766 106168 77818
rect 105922 77764 105928 77766
rect 105984 77764 106008 77766
rect 106064 77764 106088 77766
rect 106144 77764 106168 77766
rect 106224 77764 106230 77766
rect 105922 77755 106230 77764
rect 106280 77444 106332 77450
rect 106280 77386 106332 77392
rect 106292 77042 106320 77386
rect 106658 77276 106966 77285
rect 106658 77274 106664 77276
rect 106720 77274 106744 77276
rect 106800 77274 106824 77276
rect 106880 77274 106904 77276
rect 106960 77274 106966 77276
rect 106720 77222 106722 77274
rect 106902 77222 106904 77274
rect 106658 77220 106664 77222
rect 106720 77220 106744 77222
rect 106800 77220 106824 77222
rect 106880 77220 106904 77222
rect 106960 77220 106966 77222
rect 106658 77211 106966 77220
rect 106280 77036 106332 77042
rect 106280 76978 106332 76984
rect 105820 76900 105872 76906
rect 105820 76842 105872 76848
rect 107672 76430 107700 77998
rect 108132 77586 108160 78406
rect 108500 78305 108528 78406
rect 108486 78296 108542 78305
rect 108486 78231 108542 78240
rect 108488 77920 108540 77926
rect 108488 77862 108540 77868
rect 108500 77625 108528 77862
rect 108486 77616 108542 77625
rect 108120 77580 108172 77586
rect 108486 77551 108542 77560
rect 108120 77522 108172 77528
rect 108486 76936 108542 76945
rect 108486 76871 108488 76880
rect 108540 76871 108542 76880
rect 108488 76842 108540 76848
rect 107660 76424 107712 76430
rect 107660 76366 107712 76372
rect 108120 76356 108172 76362
rect 108120 76298 108172 76304
rect 108132 76090 108160 76298
rect 108488 76288 108540 76294
rect 108486 76256 108488 76265
rect 108540 76256 108542 76265
rect 108486 76191 108542 76200
rect 108120 76084 108172 76090
rect 108120 76026 108172 76032
rect 108488 76084 108540 76090
rect 108488 76026 108540 76032
rect 108120 75744 108172 75750
rect 108120 75686 108172 75692
rect 108132 73370 108160 75686
rect 108500 75585 108528 76026
rect 108486 75576 108542 75585
rect 108486 75511 108542 75520
rect 108488 75200 108540 75206
rect 108488 75142 108540 75148
rect 108500 74905 108528 75142
rect 108486 74896 108542 74905
rect 108486 74831 108542 74840
rect 108486 74216 108542 74225
rect 108486 74151 108542 74160
rect 108500 74118 108528 74151
rect 108488 74112 108540 74118
rect 108488 74054 108540 74060
rect 108488 73568 108540 73574
rect 108486 73536 108488 73545
rect 108540 73536 108542 73545
rect 108486 73471 108542 73480
rect 108120 73364 108172 73370
rect 108120 73306 108172 73312
rect 108132 73166 108160 73306
rect 108120 73160 108172 73166
rect 108120 73102 108172 73108
rect 108488 73024 108540 73030
rect 108488 72966 108540 72972
rect 108500 72865 108528 72966
rect 108486 72856 108542 72865
rect 108486 72791 108542 72800
rect 104348 72480 104400 72486
rect 104348 72422 104400 72428
rect 107936 68672 107988 68678
rect 107936 68614 107988 68620
rect 107948 67930 107976 68614
rect 107936 67924 107988 67930
rect 107936 67866 107988 67872
rect 108488 67720 108540 67726
rect 108488 67662 108540 67668
rect 102968 67652 103020 67658
rect 102968 67594 103020 67600
rect 108500 67425 108528 67662
rect 108486 67416 108542 67425
rect 108486 67351 108542 67360
rect 102324 66632 102376 66638
rect 102324 66574 102376 66580
rect 102230 25088 102286 25097
rect 102230 25023 102286 25032
rect 102336 22778 102364 66574
rect 106658 66396 106966 66405
rect 106658 66394 106664 66396
rect 106720 66394 106744 66396
rect 106800 66394 106824 66396
rect 106880 66394 106904 66396
rect 106960 66394 106966 66396
rect 106720 66342 106722 66394
rect 106902 66342 106904 66394
rect 106658 66340 106664 66342
rect 106720 66340 106744 66342
rect 106800 66340 106824 66342
rect 106880 66340 106904 66342
rect 106960 66340 106966 66342
rect 106658 66331 106966 66340
rect 105922 65852 106230 65861
rect 105922 65850 105928 65852
rect 105984 65850 106008 65852
rect 106064 65850 106088 65852
rect 106144 65850 106168 65852
rect 106224 65850 106230 65852
rect 105984 65798 105986 65850
rect 106166 65798 106168 65850
rect 105922 65796 105928 65798
rect 105984 65796 106008 65798
rect 106064 65796 106088 65798
rect 106144 65796 106168 65798
rect 106224 65796 106230 65798
rect 105922 65787 106230 65796
rect 103520 65680 103572 65686
rect 103520 65622 103572 65628
rect 102600 25152 102652 25158
rect 102598 25120 102600 25129
rect 102652 25120 102654 25129
rect 102598 25055 102654 25064
rect 102324 22772 102376 22778
rect 102324 22714 102376 22720
rect 102336 22269 102364 22714
rect 102322 22260 102378 22269
rect 102322 22195 102378 22204
rect 103532 9586 103560 65622
rect 103612 65544 103664 65550
rect 103612 65486 103664 65492
rect 103624 9654 103652 65486
rect 106658 65308 106966 65317
rect 106658 65306 106664 65308
rect 106720 65306 106744 65308
rect 106800 65306 106824 65308
rect 106880 65306 106904 65308
rect 106960 65306 106966 65308
rect 106720 65254 106722 65306
rect 106902 65254 106904 65306
rect 106658 65252 106664 65254
rect 106720 65252 106744 65254
rect 106800 65252 106824 65254
rect 106880 65252 106904 65254
rect 106960 65252 106966 65254
rect 106658 65243 106966 65252
rect 105922 64764 106230 64773
rect 105922 64762 105928 64764
rect 105984 64762 106008 64764
rect 106064 64762 106088 64764
rect 106144 64762 106168 64764
rect 106224 64762 106230 64764
rect 105984 64710 105986 64762
rect 106166 64710 106168 64762
rect 105922 64708 105928 64710
rect 105984 64708 106008 64710
rect 106064 64708 106088 64710
rect 106144 64708 106168 64710
rect 106224 64708 106230 64710
rect 105922 64699 106230 64708
rect 106658 64220 106966 64229
rect 106658 64218 106664 64220
rect 106720 64218 106744 64220
rect 106800 64218 106824 64220
rect 106880 64218 106904 64220
rect 106960 64218 106966 64220
rect 106720 64166 106722 64218
rect 106902 64166 106904 64218
rect 106658 64164 106664 64166
rect 106720 64164 106744 64166
rect 106800 64164 106824 64166
rect 106880 64164 106904 64166
rect 106960 64164 106966 64166
rect 106658 64155 106966 64164
rect 105922 63676 106230 63685
rect 105922 63674 105928 63676
rect 105984 63674 106008 63676
rect 106064 63674 106088 63676
rect 106144 63674 106168 63676
rect 106224 63674 106230 63676
rect 105984 63622 105986 63674
rect 106166 63622 106168 63674
rect 105922 63620 105928 63622
rect 105984 63620 106008 63622
rect 106064 63620 106088 63622
rect 106144 63620 106168 63622
rect 106224 63620 106230 63622
rect 105922 63611 106230 63620
rect 106658 63132 106966 63141
rect 106658 63130 106664 63132
rect 106720 63130 106744 63132
rect 106800 63130 106824 63132
rect 106880 63130 106904 63132
rect 106960 63130 106966 63132
rect 106720 63078 106722 63130
rect 106902 63078 106904 63130
rect 106658 63076 106664 63078
rect 106720 63076 106744 63078
rect 106800 63076 106824 63078
rect 106880 63076 106904 63078
rect 106960 63076 106966 63078
rect 106658 63067 106966 63076
rect 105922 62588 106230 62597
rect 105922 62586 105928 62588
rect 105984 62586 106008 62588
rect 106064 62586 106088 62588
rect 106144 62586 106168 62588
rect 106224 62586 106230 62588
rect 105984 62534 105986 62586
rect 106166 62534 106168 62586
rect 105922 62532 105928 62534
rect 105984 62532 106008 62534
rect 106064 62532 106088 62534
rect 106144 62532 106168 62534
rect 106224 62532 106230 62534
rect 105922 62523 106230 62532
rect 106658 62044 106966 62053
rect 106658 62042 106664 62044
rect 106720 62042 106744 62044
rect 106800 62042 106824 62044
rect 106880 62042 106904 62044
rect 106960 62042 106966 62044
rect 106720 61990 106722 62042
rect 106902 61990 106904 62042
rect 106658 61988 106664 61990
rect 106720 61988 106744 61990
rect 106800 61988 106824 61990
rect 106880 61988 106904 61990
rect 106960 61988 106966 61990
rect 106658 61979 106966 61988
rect 105922 61500 106230 61509
rect 105922 61498 105928 61500
rect 105984 61498 106008 61500
rect 106064 61498 106088 61500
rect 106144 61498 106168 61500
rect 106224 61498 106230 61500
rect 105984 61446 105986 61498
rect 106166 61446 106168 61498
rect 105922 61444 105928 61446
rect 105984 61444 106008 61446
rect 106064 61444 106088 61446
rect 106144 61444 106168 61446
rect 106224 61444 106230 61446
rect 105922 61435 106230 61444
rect 106658 60956 106966 60965
rect 106658 60954 106664 60956
rect 106720 60954 106744 60956
rect 106800 60954 106824 60956
rect 106880 60954 106904 60956
rect 106960 60954 106966 60956
rect 106720 60902 106722 60954
rect 106902 60902 106904 60954
rect 106658 60900 106664 60902
rect 106720 60900 106744 60902
rect 106800 60900 106824 60902
rect 106880 60900 106904 60902
rect 106960 60900 106966 60902
rect 106658 60891 106966 60900
rect 105922 60412 106230 60421
rect 105922 60410 105928 60412
rect 105984 60410 106008 60412
rect 106064 60410 106088 60412
rect 106144 60410 106168 60412
rect 106224 60410 106230 60412
rect 105984 60358 105986 60410
rect 106166 60358 106168 60410
rect 105922 60356 105928 60358
rect 105984 60356 106008 60358
rect 106064 60356 106088 60358
rect 106144 60356 106168 60358
rect 106224 60356 106230 60358
rect 105922 60347 106230 60356
rect 104348 60104 104400 60110
rect 104348 60046 104400 60052
rect 104360 59809 104388 60046
rect 106658 59868 106966 59877
rect 106658 59866 106664 59868
rect 106720 59866 106744 59868
rect 106800 59866 106824 59868
rect 106880 59866 106904 59868
rect 106960 59866 106966 59868
rect 106720 59814 106722 59866
rect 106902 59814 106904 59866
rect 106658 59812 106664 59814
rect 106720 59812 106744 59814
rect 106800 59812 106824 59814
rect 106880 59812 106904 59814
rect 106960 59812 106966 59814
rect 104346 59800 104402 59809
rect 106658 59803 106966 59812
rect 104346 59735 104402 59744
rect 105922 59324 106230 59333
rect 105922 59322 105928 59324
rect 105984 59322 106008 59324
rect 106064 59322 106088 59324
rect 106144 59322 106168 59324
rect 106224 59322 106230 59324
rect 105984 59270 105986 59322
rect 106166 59270 106168 59322
rect 105922 59268 105928 59270
rect 105984 59268 106008 59270
rect 106064 59268 106088 59270
rect 106144 59268 106168 59270
rect 106224 59268 106230 59270
rect 105922 59259 106230 59268
rect 106658 58780 106966 58789
rect 106658 58778 106664 58780
rect 106720 58778 106744 58780
rect 106800 58778 106824 58780
rect 106880 58778 106904 58780
rect 106960 58778 106966 58780
rect 106720 58726 106722 58778
rect 106902 58726 106904 58778
rect 106658 58724 106664 58726
rect 106720 58724 106744 58726
rect 106800 58724 106824 58726
rect 106880 58724 106904 58726
rect 106960 58724 106966 58726
rect 106658 58715 106966 58724
rect 105922 58236 106230 58245
rect 105922 58234 105928 58236
rect 105984 58234 106008 58236
rect 106064 58234 106088 58236
rect 106144 58234 106168 58236
rect 106224 58234 106230 58236
rect 105984 58182 105986 58234
rect 106166 58182 106168 58234
rect 105922 58180 105928 58182
rect 105984 58180 106008 58182
rect 106064 58180 106088 58182
rect 106144 58180 106168 58182
rect 106224 58180 106230 58182
rect 105922 58171 106230 58180
rect 106658 57692 106966 57701
rect 106658 57690 106664 57692
rect 106720 57690 106744 57692
rect 106800 57690 106824 57692
rect 106880 57690 106904 57692
rect 106960 57690 106966 57692
rect 106720 57638 106722 57690
rect 106902 57638 106904 57690
rect 106658 57636 106664 57638
rect 106720 57636 106744 57638
rect 106800 57636 106824 57638
rect 106880 57636 106904 57638
rect 106960 57636 106966 57638
rect 106658 57627 106966 57636
rect 105922 57148 106230 57157
rect 105922 57146 105928 57148
rect 105984 57146 106008 57148
rect 106064 57146 106088 57148
rect 106144 57146 106168 57148
rect 106224 57146 106230 57148
rect 105984 57094 105986 57146
rect 106166 57094 106168 57146
rect 105922 57092 105928 57094
rect 105984 57092 106008 57094
rect 106064 57092 106088 57094
rect 106144 57092 106168 57094
rect 106224 57092 106230 57094
rect 105922 57083 106230 57092
rect 106658 56604 106966 56613
rect 106658 56602 106664 56604
rect 106720 56602 106744 56604
rect 106800 56602 106824 56604
rect 106880 56602 106904 56604
rect 106960 56602 106966 56604
rect 106720 56550 106722 56602
rect 106902 56550 106904 56602
rect 106658 56548 106664 56550
rect 106720 56548 106744 56550
rect 106800 56548 106824 56550
rect 106880 56548 106904 56550
rect 106960 56548 106966 56550
rect 106658 56539 106966 56548
rect 105922 56060 106230 56069
rect 105922 56058 105928 56060
rect 105984 56058 106008 56060
rect 106064 56058 106088 56060
rect 106144 56058 106168 56060
rect 106224 56058 106230 56060
rect 105984 56006 105986 56058
rect 106166 56006 106168 56058
rect 105922 56004 105928 56006
rect 105984 56004 106008 56006
rect 106064 56004 106088 56006
rect 106144 56004 106168 56006
rect 106224 56004 106230 56006
rect 105922 55995 106230 56004
rect 106658 55516 106966 55525
rect 106658 55514 106664 55516
rect 106720 55514 106744 55516
rect 106800 55514 106824 55516
rect 106880 55514 106904 55516
rect 106960 55514 106966 55516
rect 106720 55462 106722 55514
rect 106902 55462 106904 55514
rect 106658 55460 106664 55462
rect 106720 55460 106744 55462
rect 106800 55460 106824 55462
rect 106880 55460 106904 55462
rect 106960 55460 106966 55462
rect 106658 55451 106966 55460
rect 105922 54972 106230 54981
rect 105922 54970 105928 54972
rect 105984 54970 106008 54972
rect 106064 54970 106088 54972
rect 106144 54970 106168 54972
rect 106224 54970 106230 54972
rect 105984 54918 105986 54970
rect 106166 54918 106168 54970
rect 105922 54916 105928 54918
rect 105984 54916 106008 54918
rect 106064 54916 106088 54918
rect 106144 54916 106168 54918
rect 106224 54916 106230 54918
rect 105922 54907 106230 54916
rect 106658 54428 106966 54437
rect 106658 54426 106664 54428
rect 106720 54426 106744 54428
rect 106800 54426 106824 54428
rect 106880 54426 106904 54428
rect 106960 54426 106966 54428
rect 106720 54374 106722 54426
rect 106902 54374 106904 54426
rect 106658 54372 106664 54374
rect 106720 54372 106744 54374
rect 106800 54372 106824 54374
rect 106880 54372 106904 54374
rect 106960 54372 106966 54374
rect 106658 54363 106966 54372
rect 105922 53884 106230 53893
rect 105922 53882 105928 53884
rect 105984 53882 106008 53884
rect 106064 53882 106088 53884
rect 106144 53882 106168 53884
rect 106224 53882 106230 53884
rect 105984 53830 105986 53882
rect 106166 53830 106168 53882
rect 105922 53828 105928 53830
rect 105984 53828 106008 53830
rect 106064 53828 106088 53830
rect 106144 53828 106168 53830
rect 106224 53828 106230 53830
rect 105922 53819 106230 53828
rect 106658 53340 106966 53349
rect 106658 53338 106664 53340
rect 106720 53338 106744 53340
rect 106800 53338 106824 53340
rect 106880 53338 106904 53340
rect 106960 53338 106966 53340
rect 106720 53286 106722 53338
rect 106902 53286 106904 53338
rect 106658 53284 106664 53286
rect 106720 53284 106744 53286
rect 106800 53284 106824 53286
rect 106880 53284 106904 53286
rect 106960 53284 106966 53286
rect 106658 53275 106966 53284
rect 105922 52796 106230 52805
rect 105922 52794 105928 52796
rect 105984 52794 106008 52796
rect 106064 52794 106088 52796
rect 106144 52794 106168 52796
rect 106224 52794 106230 52796
rect 105984 52742 105986 52794
rect 106166 52742 106168 52794
rect 105922 52740 105928 52742
rect 105984 52740 106008 52742
rect 106064 52740 106088 52742
rect 106144 52740 106168 52742
rect 106224 52740 106230 52742
rect 105922 52731 106230 52740
rect 106658 52252 106966 52261
rect 106658 52250 106664 52252
rect 106720 52250 106744 52252
rect 106800 52250 106824 52252
rect 106880 52250 106904 52252
rect 106960 52250 106966 52252
rect 106720 52198 106722 52250
rect 106902 52198 106904 52250
rect 106658 52196 106664 52198
rect 106720 52196 106744 52198
rect 106800 52196 106824 52198
rect 106880 52196 106904 52198
rect 106960 52196 106966 52198
rect 106658 52187 106966 52196
rect 105922 51708 106230 51717
rect 105922 51706 105928 51708
rect 105984 51706 106008 51708
rect 106064 51706 106088 51708
rect 106144 51706 106168 51708
rect 106224 51706 106230 51708
rect 105984 51654 105986 51706
rect 106166 51654 106168 51706
rect 105922 51652 105928 51654
rect 105984 51652 106008 51654
rect 106064 51652 106088 51654
rect 106144 51652 106168 51654
rect 106224 51652 106230 51654
rect 105922 51643 106230 51652
rect 106658 51164 106966 51173
rect 106658 51162 106664 51164
rect 106720 51162 106744 51164
rect 106800 51162 106824 51164
rect 106880 51162 106904 51164
rect 106960 51162 106966 51164
rect 106720 51110 106722 51162
rect 106902 51110 106904 51162
rect 106658 51108 106664 51110
rect 106720 51108 106744 51110
rect 106800 51108 106824 51110
rect 106880 51108 106904 51110
rect 106960 51108 106966 51110
rect 106658 51099 106966 51108
rect 105922 50620 106230 50629
rect 105922 50618 105928 50620
rect 105984 50618 106008 50620
rect 106064 50618 106088 50620
rect 106144 50618 106168 50620
rect 106224 50618 106230 50620
rect 105984 50566 105986 50618
rect 106166 50566 106168 50618
rect 105922 50564 105928 50566
rect 105984 50564 106008 50566
rect 106064 50564 106088 50566
rect 106144 50564 106168 50566
rect 106224 50564 106230 50566
rect 105922 50555 106230 50564
rect 106658 50076 106966 50085
rect 106658 50074 106664 50076
rect 106720 50074 106744 50076
rect 106800 50074 106824 50076
rect 106880 50074 106904 50076
rect 106960 50074 106966 50076
rect 106720 50022 106722 50074
rect 106902 50022 106904 50074
rect 106658 50020 106664 50022
rect 106720 50020 106744 50022
rect 106800 50020 106824 50022
rect 106880 50020 106904 50022
rect 106960 50020 106966 50022
rect 106658 50011 106966 50020
rect 105922 49532 106230 49541
rect 105922 49530 105928 49532
rect 105984 49530 106008 49532
rect 106064 49530 106088 49532
rect 106144 49530 106168 49532
rect 106224 49530 106230 49532
rect 105984 49478 105986 49530
rect 106166 49478 106168 49530
rect 105922 49476 105928 49478
rect 105984 49476 106008 49478
rect 106064 49476 106088 49478
rect 106144 49476 106168 49478
rect 106224 49476 106230 49478
rect 105922 49467 106230 49476
rect 106658 48988 106966 48997
rect 106658 48986 106664 48988
rect 106720 48986 106744 48988
rect 106800 48986 106824 48988
rect 106880 48986 106904 48988
rect 106960 48986 106966 48988
rect 106720 48934 106722 48986
rect 106902 48934 106904 48986
rect 106658 48932 106664 48934
rect 106720 48932 106744 48934
rect 106800 48932 106824 48934
rect 106880 48932 106904 48934
rect 106960 48932 106966 48934
rect 106658 48923 106966 48932
rect 105922 48444 106230 48453
rect 105922 48442 105928 48444
rect 105984 48442 106008 48444
rect 106064 48442 106088 48444
rect 106144 48442 106168 48444
rect 106224 48442 106230 48444
rect 105984 48390 105986 48442
rect 106166 48390 106168 48442
rect 105922 48388 105928 48390
rect 105984 48388 106008 48390
rect 106064 48388 106088 48390
rect 106144 48388 106168 48390
rect 106224 48388 106230 48390
rect 105922 48379 106230 48388
rect 106658 47900 106966 47909
rect 106658 47898 106664 47900
rect 106720 47898 106744 47900
rect 106800 47898 106824 47900
rect 106880 47898 106904 47900
rect 106960 47898 106966 47900
rect 106720 47846 106722 47898
rect 106902 47846 106904 47898
rect 106658 47844 106664 47846
rect 106720 47844 106744 47846
rect 106800 47844 106824 47846
rect 106880 47844 106904 47846
rect 106960 47844 106966 47846
rect 106658 47835 106966 47844
rect 105922 47356 106230 47365
rect 105922 47354 105928 47356
rect 105984 47354 106008 47356
rect 106064 47354 106088 47356
rect 106144 47354 106168 47356
rect 106224 47354 106230 47356
rect 105984 47302 105986 47354
rect 106166 47302 106168 47354
rect 105922 47300 105928 47302
rect 105984 47300 106008 47302
rect 106064 47300 106088 47302
rect 106144 47300 106168 47302
rect 106224 47300 106230 47302
rect 105922 47291 106230 47300
rect 106658 46812 106966 46821
rect 106658 46810 106664 46812
rect 106720 46810 106744 46812
rect 106800 46810 106824 46812
rect 106880 46810 106904 46812
rect 106960 46810 106966 46812
rect 106720 46758 106722 46810
rect 106902 46758 106904 46810
rect 106658 46756 106664 46758
rect 106720 46756 106744 46758
rect 106800 46756 106824 46758
rect 106880 46756 106904 46758
rect 106960 46756 106966 46758
rect 106658 46747 106966 46756
rect 105922 46268 106230 46277
rect 105922 46266 105928 46268
rect 105984 46266 106008 46268
rect 106064 46266 106088 46268
rect 106144 46266 106168 46268
rect 106224 46266 106230 46268
rect 105984 46214 105986 46266
rect 106166 46214 106168 46266
rect 105922 46212 105928 46214
rect 105984 46212 106008 46214
rect 106064 46212 106088 46214
rect 106144 46212 106168 46214
rect 106224 46212 106230 46214
rect 105922 46203 106230 46212
rect 106658 45724 106966 45733
rect 106658 45722 106664 45724
rect 106720 45722 106744 45724
rect 106800 45722 106824 45724
rect 106880 45722 106904 45724
rect 106960 45722 106966 45724
rect 106720 45670 106722 45722
rect 106902 45670 106904 45722
rect 106658 45668 106664 45670
rect 106720 45668 106744 45670
rect 106800 45668 106824 45670
rect 106880 45668 106904 45670
rect 106960 45668 106966 45670
rect 106658 45659 106966 45668
rect 105922 45180 106230 45189
rect 105922 45178 105928 45180
rect 105984 45178 106008 45180
rect 106064 45178 106088 45180
rect 106144 45178 106168 45180
rect 106224 45178 106230 45180
rect 105984 45126 105986 45178
rect 106166 45126 106168 45178
rect 105922 45124 105928 45126
rect 105984 45124 106008 45126
rect 106064 45124 106088 45126
rect 106144 45124 106168 45126
rect 106224 45124 106230 45126
rect 105922 45115 106230 45124
rect 106658 44636 106966 44645
rect 106658 44634 106664 44636
rect 106720 44634 106744 44636
rect 106800 44634 106824 44636
rect 106880 44634 106904 44636
rect 106960 44634 106966 44636
rect 106720 44582 106722 44634
rect 106902 44582 106904 44634
rect 106658 44580 106664 44582
rect 106720 44580 106744 44582
rect 106800 44580 106824 44582
rect 106880 44580 106904 44582
rect 106960 44580 106966 44582
rect 106658 44571 106966 44580
rect 105922 44092 106230 44101
rect 105922 44090 105928 44092
rect 105984 44090 106008 44092
rect 106064 44090 106088 44092
rect 106144 44090 106168 44092
rect 106224 44090 106230 44092
rect 105984 44038 105986 44090
rect 106166 44038 106168 44090
rect 105922 44036 105928 44038
rect 105984 44036 106008 44038
rect 106064 44036 106088 44038
rect 106144 44036 106168 44038
rect 106224 44036 106230 44038
rect 105922 44027 106230 44036
rect 106658 43548 106966 43557
rect 106658 43546 106664 43548
rect 106720 43546 106744 43548
rect 106800 43546 106824 43548
rect 106880 43546 106904 43548
rect 106960 43546 106966 43548
rect 106720 43494 106722 43546
rect 106902 43494 106904 43546
rect 106658 43492 106664 43494
rect 106720 43492 106744 43494
rect 106800 43492 106824 43494
rect 106880 43492 106904 43494
rect 106960 43492 106966 43494
rect 106658 43483 106966 43492
rect 105922 43004 106230 43013
rect 105922 43002 105928 43004
rect 105984 43002 106008 43004
rect 106064 43002 106088 43004
rect 106144 43002 106168 43004
rect 106224 43002 106230 43004
rect 105984 42950 105986 43002
rect 106166 42950 106168 43002
rect 105922 42948 105928 42950
rect 105984 42948 106008 42950
rect 106064 42948 106088 42950
rect 106144 42948 106168 42950
rect 106224 42948 106230 42950
rect 105922 42939 106230 42948
rect 106658 42460 106966 42469
rect 106658 42458 106664 42460
rect 106720 42458 106744 42460
rect 106800 42458 106824 42460
rect 106880 42458 106904 42460
rect 106960 42458 106966 42460
rect 106720 42406 106722 42458
rect 106902 42406 106904 42458
rect 106658 42404 106664 42406
rect 106720 42404 106744 42406
rect 106800 42404 106824 42406
rect 106880 42404 106904 42406
rect 106960 42404 106966 42406
rect 106658 42395 106966 42404
rect 105922 41916 106230 41925
rect 105922 41914 105928 41916
rect 105984 41914 106008 41916
rect 106064 41914 106088 41916
rect 106144 41914 106168 41916
rect 106224 41914 106230 41916
rect 105984 41862 105986 41914
rect 106166 41862 106168 41914
rect 105922 41860 105928 41862
rect 105984 41860 106008 41862
rect 106064 41860 106088 41862
rect 106144 41860 106168 41862
rect 106224 41860 106230 41862
rect 105922 41851 106230 41860
rect 106658 41372 106966 41381
rect 106658 41370 106664 41372
rect 106720 41370 106744 41372
rect 106800 41370 106824 41372
rect 106880 41370 106904 41372
rect 106960 41370 106966 41372
rect 106720 41318 106722 41370
rect 106902 41318 106904 41370
rect 106658 41316 106664 41318
rect 106720 41316 106744 41318
rect 106800 41316 106824 41318
rect 106880 41316 106904 41318
rect 106960 41316 106966 41318
rect 106658 41307 106966 41316
rect 105922 40828 106230 40837
rect 105922 40826 105928 40828
rect 105984 40826 106008 40828
rect 106064 40826 106088 40828
rect 106144 40826 106168 40828
rect 106224 40826 106230 40828
rect 105984 40774 105986 40826
rect 106166 40774 106168 40826
rect 105922 40772 105928 40774
rect 105984 40772 106008 40774
rect 106064 40772 106088 40774
rect 106144 40772 106168 40774
rect 106224 40772 106230 40774
rect 105922 40763 106230 40772
rect 106658 40284 106966 40293
rect 106658 40282 106664 40284
rect 106720 40282 106744 40284
rect 106800 40282 106824 40284
rect 106880 40282 106904 40284
rect 106960 40282 106966 40284
rect 106720 40230 106722 40282
rect 106902 40230 106904 40282
rect 106658 40228 106664 40230
rect 106720 40228 106744 40230
rect 106800 40228 106824 40230
rect 106880 40228 106904 40230
rect 106960 40228 106966 40230
rect 106658 40219 106966 40228
rect 105922 39740 106230 39749
rect 105922 39738 105928 39740
rect 105984 39738 106008 39740
rect 106064 39738 106088 39740
rect 106144 39738 106168 39740
rect 106224 39738 106230 39740
rect 105984 39686 105986 39738
rect 106166 39686 106168 39738
rect 105922 39684 105928 39686
rect 105984 39684 106008 39686
rect 106064 39684 106088 39686
rect 106144 39684 106168 39686
rect 106224 39684 106230 39686
rect 105922 39675 106230 39684
rect 106658 39196 106966 39205
rect 106658 39194 106664 39196
rect 106720 39194 106744 39196
rect 106800 39194 106824 39196
rect 106880 39194 106904 39196
rect 106960 39194 106966 39196
rect 106720 39142 106722 39194
rect 106902 39142 106904 39194
rect 106658 39140 106664 39142
rect 106720 39140 106744 39142
rect 106800 39140 106824 39142
rect 106880 39140 106904 39142
rect 106960 39140 106966 39142
rect 106658 39131 106966 39140
rect 105922 38652 106230 38661
rect 105922 38650 105928 38652
rect 105984 38650 106008 38652
rect 106064 38650 106088 38652
rect 106144 38650 106168 38652
rect 106224 38650 106230 38652
rect 105984 38598 105986 38650
rect 106166 38598 106168 38650
rect 105922 38596 105928 38598
rect 105984 38596 106008 38598
rect 106064 38596 106088 38598
rect 106144 38596 106168 38598
rect 106224 38596 106230 38598
rect 105922 38587 106230 38596
rect 106658 38108 106966 38117
rect 106658 38106 106664 38108
rect 106720 38106 106744 38108
rect 106800 38106 106824 38108
rect 106880 38106 106904 38108
rect 106960 38106 106966 38108
rect 106720 38054 106722 38106
rect 106902 38054 106904 38106
rect 106658 38052 106664 38054
rect 106720 38052 106744 38054
rect 106800 38052 106824 38054
rect 106880 38052 106904 38054
rect 106960 38052 106966 38054
rect 106658 38043 106966 38052
rect 105922 37564 106230 37573
rect 105922 37562 105928 37564
rect 105984 37562 106008 37564
rect 106064 37562 106088 37564
rect 106144 37562 106168 37564
rect 106224 37562 106230 37564
rect 105984 37510 105986 37562
rect 106166 37510 106168 37562
rect 105922 37508 105928 37510
rect 105984 37508 106008 37510
rect 106064 37508 106088 37510
rect 106144 37508 106168 37510
rect 106224 37508 106230 37510
rect 105922 37499 106230 37508
rect 106658 37020 106966 37029
rect 106658 37018 106664 37020
rect 106720 37018 106744 37020
rect 106800 37018 106824 37020
rect 106880 37018 106904 37020
rect 106960 37018 106966 37020
rect 106720 36966 106722 37018
rect 106902 36966 106904 37018
rect 106658 36964 106664 36966
rect 106720 36964 106744 36966
rect 106800 36964 106824 36966
rect 106880 36964 106904 36966
rect 106960 36964 106966 36966
rect 106658 36955 106966 36964
rect 105922 36476 106230 36485
rect 105922 36474 105928 36476
rect 105984 36474 106008 36476
rect 106064 36474 106088 36476
rect 106144 36474 106168 36476
rect 106224 36474 106230 36476
rect 105984 36422 105986 36474
rect 106166 36422 106168 36474
rect 105922 36420 105928 36422
rect 105984 36420 106008 36422
rect 106064 36420 106088 36422
rect 106144 36420 106168 36422
rect 106224 36420 106230 36422
rect 105922 36411 106230 36420
rect 106658 35932 106966 35941
rect 106658 35930 106664 35932
rect 106720 35930 106744 35932
rect 106800 35930 106824 35932
rect 106880 35930 106904 35932
rect 106960 35930 106966 35932
rect 106720 35878 106722 35930
rect 106902 35878 106904 35930
rect 106658 35876 106664 35878
rect 106720 35876 106744 35878
rect 106800 35876 106824 35878
rect 106880 35876 106904 35878
rect 106960 35876 106966 35878
rect 106658 35867 106966 35876
rect 105922 35388 106230 35397
rect 105922 35386 105928 35388
rect 105984 35386 106008 35388
rect 106064 35386 106088 35388
rect 106144 35386 106168 35388
rect 106224 35386 106230 35388
rect 105984 35334 105986 35386
rect 106166 35334 106168 35386
rect 105922 35332 105928 35334
rect 105984 35332 106008 35334
rect 106064 35332 106088 35334
rect 106144 35332 106168 35334
rect 106224 35332 106230 35334
rect 105922 35323 106230 35332
rect 106658 34844 106966 34853
rect 106658 34842 106664 34844
rect 106720 34842 106744 34844
rect 106800 34842 106824 34844
rect 106880 34842 106904 34844
rect 106960 34842 106966 34844
rect 106720 34790 106722 34842
rect 106902 34790 106904 34842
rect 106658 34788 106664 34790
rect 106720 34788 106744 34790
rect 106800 34788 106824 34790
rect 106880 34788 106904 34790
rect 106960 34788 106966 34790
rect 106658 34779 106966 34788
rect 105922 34300 106230 34309
rect 105922 34298 105928 34300
rect 105984 34298 106008 34300
rect 106064 34298 106088 34300
rect 106144 34298 106168 34300
rect 106224 34298 106230 34300
rect 105984 34246 105986 34298
rect 106166 34246 106168 34298
rect 105922 34244 105928 34246
rect 105984 34244 106008 34246
rect 106064 34244 106088 34246
rect 106144 34244 106168 34246
rect 106224 34244 106230 34246
rect 105922 34235 106230 34244
rect 106658 33756 106966 33765
rect 106658 33754 106664 33756
rect 106720 33754 106744 33756
rect 106800 33754 106824 33756
rect 106880 33754 106904 33756
rect 106960 33754 106966 33756
rect 106720 33702 106722 33754
rect 106902 33702 106904 33754
rect 106658 33700 106664 33702
rect 106720 33700 106744 33702
rect 106800 33700 106824 33702
rect 106880 33700 106904 33702
rect 106960 33700 106966 33702
rect 106658 33691 106966 33700
rect 105922 33212 106230 33221
rect 105922 33210 105928 33212
rect 105984 33210 106008 33212
rect 106064 33210 106088 33212
rect 106144 33210 106168 33212
rect 106224 33210 106230 33212
rect 105984 33158 105986 33210
rect 106166 33158 106168 33210
rect 105922 33156 105928 33158
rect 105984 33156 106008 33158
rect 106064 33156 106088 33158
rect 106144 33156 106168 33158
rect 106224 33156 106230 33158
rect 105922 33147 106230 33156
rect 106658 32668 106966 32677
rect 106658 32666 106664 32668
rect 106720 32666 106744 32668
rect 106800 32666 106824 32668
rect 106880 32666 106904 32668
rect 106960 32666 106966 32668
rect 106720 32614 106722 32666
rect 106902 32614 106904 32666
rect 106658 32612 106664 32614
rect 106720 32612 106744 32614
rect 106800 32612 106824 32614
rect 106880 32612 106904 32614
rect 106960 32612 106966 32614
rect 106658 32603 106966 32612
rect 105922 32124 106230 32133
rect 105922 32122 105928 32124
rect 105984 32122 106008 32124
rect 106064 32122 106088 32124
rect 106144 32122 106168 32124
rect 106224 32122 106230 32124
rect 105984 32070 105986 32122
rect 106166 32070 106168 32122
rect 105922 32068 105928 32070
rect 105984 32068 106008 32070
rect 106064 32068 106088 32070
rect 106144 32068 106168 32070
rect 106224 32068 106230 32070
rect 105922 32059 106230 32068
rect 106658 31580 106966 31589
rect 106658 31578 106664 31580
rect 106720 31578 106744 31580
rect 106800 31578 106824 31580
rect 106880 31578 106904 31580
rect 106960 31578 106966 31580
rect 106720 31526 106722 31578
rect 106902 31526 106904 31578
rect 106658 31524 106664 31526
rect 106720 31524 106744 31526
rect 106800 31524 106824 31526
rect 106880 31524 106904 31526
rect 106960 31524 106966 31526
rect 106658 31515 106966 31524
rect 105922 31036 106230 31045
rect 105922 31034 105928 31036
rect 105984 31034 106008 31036
rect 106064 31034 106088 31036
rect 106144 31034 106168 31036
rect 106224 31034 106230 31036
rect 105984 30982 105986 31034
rect 106166 30982 106168 31034
rect 105922 30980 105928 30982
rect 105984 30980 106008 30982
rect 106064 30980 106088 30982
rect 106144 30980 106168 30982
rect 106224 30980 106230 30982
rect 105922 30971 106230 30980
rect 106658 30492 106966 30501
rect 106658 30490 106664 30492
rect 106720 30490 106744 30492
rect 106800 30490 106824 30492
rect 106880 30490 106904 30492
rect 106960 30490 106966 30492
rect 106720 30438 106722 30490
rect 106902 30438 106904 30490
rect 106658 30436 106664 30438
rect 106720 30436 106744 30438
rect 106800 30436 106824 30438
rect 106880 30436 106904 30438
rect 106960 30436 106966 30438
rect 106658 30427 106966 30436
rect 105922 29948 106230 29957
rect 105922 29946 105928 29948
rect 105984 29946 106008 29948
rect 106064 29946 106088 29948
rect 106144 29946 106168 29948
rect 106224 29946 106230 29948
rect 105984 29894 105986 29946
rect 106166 29894 106168 29946
rect 105922 29892 105928 29894
rect 105984 29892 106008 29894
rect 106064 29892 106088 29894
rect 106144 29892 106168 29894
rect 106224 29892 106230 29894
rect 105922 29883 106230 29892
rect 106658 29404 106966 29413
rect 106658 29402 106664 29404
rect 106720 29402 106744 29404
rect 106800 29402 106824 29404
rect 106880 29402 106904 29404
rect 106960 29402 106966 29404
rect 106720 29350 106722 29402
rect 106902 29350 106904 29402
rect 106658 29348 106664 29350
rect 106720 29348 106744 29350
rect 106800 29348 106824 29350
rect 106880 29348 106904 29350
rect 106960 29348 106966 29350
rect 106658 29339 106966 29348
rect 105922 28860 106230 28869
rect 105922 28858 105928 28860
rect 105984 28858 106008 28860
rect 106064 28858 106088 28860
rect 106144 28858 106168 28860
rect 106224 28858 106230 28860
rect 105984 28806 105986 28858
rect 106166 28806 106168 28858
rect 105922 28804 105928 28806
rect 105984 28804 106008 28806
rect 106064 28804 106088 28806
rect 106144 28804 106168 28806
rect 106224 28804 106230 28806
rect 105922 28795 106230 28804
rect 106658 28316 106966 28325
rect 106658 28314 106664 28316
rect 106720 28314 106744 28316
rect 106800 28314 106824 28316
rect 106880 28314 106904 28316
rect 106960 28314 106966 28316
rect 106720 28262 106722 28314
rect 106902 28262 106904 28314
rect 106658 28260 106664 28262
rect 106720 28260 106744 28262
rect 106800 28260 106824 28262
rect 106880 28260 106904 28262
rect 106960 28260 106966 28262
rect 106658 28251 106966 28260
rect 105922 27772 106230 27781
rect 105922 27770 105928 27772
rect 105984 27770 106008 27772
rect 106064 27770 106088 27772
rect 106144 27770 106168 27772
rect 106224 27770 106230 27772
rect 105984 27718 105986 27770
rect 106166 27718 106168 27770
rect 105922 27716 105928 27718
rect 105984 27716 106008 27718
rect 106064 27716 106088 27718
rect 106144 27716 106168 27718
rect 106224 27716 106230 27718
rect 105922 27707 106230 27716
rect 106658 27228 106966 27237
rect 106658 27226 106664 27228
rect 106720 27226 106744 27228
rect 106800 27226 106824 27228
rect 106880 27226 106904 27228
rect 106960 27226 106966 27228
rect 106720 27174 106722 27226
rect 106902 27174 106904 27226
rect 106658 27172 106664 27174
rect 106720 27172 106744 27174
rect 106800 27172 106824 27174
rect 106880 27172 106904 27174
rect 106960 27172 106966 27174
rect 106658 27163 106966 27172
rect 105922 26684 106230 26693
rect 105922 26682 105928 26684
rect 105984 26682 106008 26684
rect 106064 26682 106088 26684
rect 106144 26682 106168 26684
rect 106224 26682 106230 26684
rect 105984 26630 105986 26682
rect 106166 26630 106168 26682
rect 105922 26628 105928 26630
rect 105984 26628 106008 26630
rect 106064 26628 106088 26630
rect 106144 26628 106168 26630
rect 106224 26628 106230 26630
rect 105922 26619 106230 26628
rect 106658 26140 106966 26149
rect 106658 26138 106664 26140
rect 106720 26138 106744 26140
rect 106800 26138 106824 26140
rect 106880 26138 106904 26140
rect 106960 26138 106966 26140
rect 106720 26086 106722 26138
rect 106902 26086 106904 26138
rect 106658 26084 106664 26086
rect 106720 26084 106744 26086
rect 106800 26084 106824 26086
rect 106880 26084 106904 26086
rect 106960 26084 106966 26086
rect 106658 26075 106966 26084
rect 105922 25596 106230 25605
rect 105922 25594 105928 25596
rect 105984 25594 106008 25596
rect 106064 25594 106088 25596
rect 106144 25594 106168 25596
rect 106224 25594 106230 25596
rect 105984 25542 105986 25594
rect 106166 25542 106168 25594
rect 105922 25540 105928 25542
rect 105984 25540 106008 25542
rect 106064 25540 106088 25542
rect 106144 25540 106168 25542
rect 106224 25540 106230 25542
rect 105922 25531 106230 25540
rect 106658 25052 106966 25061
rect 106658 25050 106664 25052
rect 106720 25050 106744 25052
rect 106800 25050 106824 25052
rect 106880 25050 106904 25052
rect 106960 25050 106966 25052
rect 106720 24998 106722 25050
rect 106902 24998 106904 25050
rect 106658 24996 106664 24998
rect 106720 24996 106744 24998
rect 106800 24996 106824 24998
rect 106880 24996 106904 24998
rect 106960 24996 106966 24998
rect 106658 24987 106966 24996
rect 105922 24508 106230 24517
rect 105922 24506 105928 24508
rect 105984 24506 106008 24508
rect 106064 24506 106088 24508
rect 106144 24506 106168 24508
rect 106224 24506 106230 24508
rect 105984 24454 105986 24506
rect 106166 24454 106168 24506
rect 105922 24452 105928 24454
rect 105984 24452 106008 24454
rect 106064 24452 106088 24454
rect 106144 24452 106168 24454
rect 106224 24452 106230 24454
rect 105922 24443 106230 24452
rect 106658 23964 106966 23973
rect 106658 23962 106664 23964
rect 106720 23962 106744 23964
rect 106800 23962 106824 23964
rect 106880 23962 106904 23964
rect 106960 23962 106966 23964
rect 106720 23910 106722 23962
rect 106902 23910 106904 23962
rect 106658 23908 106664 23910
rect 106720 23908 106744 23910
rect 106800 23908 106824 23910
rect 106880 23908 106904 23910
rect 106960 23908 106966 23910
rect 106658 23899 106966 23908
rect 105922 23420 106230 23429
rect 105922 23418 105928 23420
rect 105984 23418 106008 23420
rect 106064 23418 106088 23420
rect 106144 23418 106168 23420
rect 106224 23418 106230 23420
rect 105984 23366 105986 23418
rect 106166 23366 106168 23418
rect 105922 23364 105928 23366
rect 105984 23364 106008 23366
rect 106064 23364 106088 23366
rect 106144 23364 106168 23366
rect 106224 23364 106230 23366
rect 105922 23355 106230 23364
rect 106658 22876 106966 22885
rect 106658 22874 106664 22876
rect 106720 22874 106744 22876
rect 106800 22874 106824 22876
rect 106880 22874 106904 22876
rect 106960 22874 106966 22876
rect 106720 22822 106722 22874
rect 106902 22822 106904 22874
rect 106658 22820 106664 22822
rect 106720 22820 106744 22822
rect 106800 22820 106824 22822
rect 106880 22820 106904 22822
rect 106960 22820 106966 22822
rect 106658 22811 106966 22820
rect 105922 22332 106230 22341
rect 105922 22330 105928 22332
rect 105984 22330 106008 22332
rect 106064 22330 106088 22332
rect 106144 22330 106168 22332
rect 106224 22330 106230 22332
rect 105984 22278 105986 22330
rect 106166 22278 106168 22330
rect 105922 22276 105928 22278
rect 105984 22276 106008 22278
rect 106064 22276 106088 22278
rect 106144 22276 106168 22278
rect 106224 22276 106230 22278
rect 105922 22267 106230 22276
rect 106658 21788 106966 21797
rect 106658 21786 106664 21788
rect 106720 21786 106744 21788
rect 106800 21786 106824 21788
rect 106880 21786 106904 21788
rect 106960 21786 106966 21788
rect 106720 21734 106722 21786
rect 106902 21734 106904 21786
rect 106658 21732 106664 21734
rect 106720 21732 106744 21734
rect 106800 21732 106824 21734
rect 106880 21732 106904 21734
rect 106960 21732 106966 21734
rect 106658 21723 106966 21732
rect 105922 21244 106230 21253
rect 105922 21242 105928 21244
rect 105984 21242 106008 21244
rect 106064 21242 106088 21244
rect 106144 21242 106168 21244
rect 106224 21242 106230 21244
rect 105984 21190 105986 21242
rect 106166 21190 106168 21242
rect 105922 21188 105928 21190
rect 105984 21188 106008 21190
rect 106064 21188 106088 21190
rect 106144 21188 106168 21190
rect 106224 21188 106230 21190
rect 105922 21179 106230 21188
rect 106658 20700 106966 20709
rect 106658 20698 106664 20700
rect 106720 20698 106744 20700
rect 106800 20698 106824 20700
rect 106880 20698 106904 20700
rect 106960 20698 106966 20700
rect 106720 20646 106722 20698
rect 106902 20646 106904 20698
rect 106658 20644 106664 20646
rect 106720 20644 106744 20646
rect 106800 20644 106824 20646
rect 106880 20644 106904 20646
rect 106960 20644 106966 20646
rect 106658 20635 106966 20644
rect 105922 20156 106230 20165
rect 105922 20154 105928 20156
rect 105984 20154 106008 20156
rect 106064 20154 106088 20156
rect 106144 20154 106168 20156
rect 106224 20154 106230 20156
rect 105984 20102 105986 20154
rect 106166 20102 106168 20154
rect 105922 20100 105928 20102
rect 105984 20100 106008 20102
rect 106064 20100 106088 20102
rect 106144 20100 106168 20102
rect 106224 20100 106230 20102
rect 105922 20091 106230 20100
rect 106658 19612 106966 19621
rect 106658 19610 106664 19612
rect 106720 19610 106744 19612
rect 106800 19610 106824 19612
rect 106880 19610 106904 19612
rect 106960 19610 106966 19612
rect 106720 19558 106722 19610
rect 106902 19558 106904 19610
rect 106658 19556 106664 19558
rect 106720 19556 106744 19558
rect 106800 19556 106824 19558
rect 106880 19556 106904 19558
rect 106960 19556 106966 19558
rect 106658 19547 106966 19556
rect 105922 19068 106230 19077
rect 105922 19066 105928 19068
rect 105984 19066 106008 19068
rect 106064 19066 106088 19068
rect 106144 19066 106168 19068
rect 106224 19066 106230 19068
rect 105984 19014 105986 19066
rect 106166 19014 106168 19066
rect 105922 19012 105928 19014
rect 105984 19012 106008 19014
rect 106064 19012 106088 19014
rect 106144 19012 106168 19014
rect 106224 19012 106230 19014
rect 105922 19003 106230 19012
rect 106658 18524 106966 18533
rect 106658 18522 106664 18524
rect 106720 18522 106744 18524
rect 106800 18522 106824 18524
rect 106880 18522 106904 18524
rect 106960 18522 106966 18524
rect 106720 18470 106722 18522
rect 106902 18470 106904 18522
rect 106658 18468 106664 18470
rect 106720 18468 106744 18470
rect 106800 18468 106824 18470
rect 106880 18468 106904 18470
rect 106960 18468 106966 18470
rect 106658 18459 106966 18468
rect 105922 17980 106230 17989
rect 105922 17978 105928 17980
rect 105984 17978 106008 17980
rect 106064 17978 106088 17980
rect 106144 17978 106168 17980
rect 106224 17978 106230 17980
rect 105984 17926 105986 17978
rect 106166 17926 106168 17978
rect 105922 17924 105928 17926
rect 105984 17924 106008 17926
rect 106064 17924 106088 17926
rect 106144 17924 106168 17926
rect 106224 17924 106230 17926
rect 105922 17915 106230 17924
rect 106658 17436 106966 17445
rect 106658 17434 106664 17436
rect 106720 17434 106744 17436
rect 106800 17434 106824 17436
rect 106880 17434 106904 17436
rect 106960 17434 106966 17436
rect 106720 17382 106722 17434
rect 106902 17382 106904 17434
rect 106658 17380 106664 17382
rect 106720 17380 106744 17382
rect 106800 17380 106824 17382
rect 106880 17380 106904 17382
rect 106960 17380 106966 17382
rect 106658 17371 106966 17380
rect 105922 16892 106230 16901
rect 105922 16890 105928 16892
rect 105984 16890 106008 16892
rect 106064 16890 106088 16892
rect 106144 16890 106168 16892
rect 106224 16890 106230 16892
rect 105984 16838 105986 16890
rect 106166 16838 106168 16890
rect 105922 16836 105928 16838
rect 105984 16836 106008 16838
rect 106064 16836 106088 16838
rect 106144 16836 106168 16838
rect 106224 16836 106230 16838
rect 105922 16827 106230 16836
rect 106658 16348 106966 16357
rect 106658 16346 106664 16348
rect 106720 16346 106744 16348
rect 106800 16346 106824 16348
rect 106880 16346 106904 16348
rect 106960 16346 106966 16348
rect 106720 16294 106722 16346
rect 106902 16294 106904 16346
rect 106658 16292 106664 16294
rect 106720 16292 106744 16294
rect 106800 16292 106824 16294
rect 106880 16292 106904 16294
rect 106960 16292 106966 16294
rect 106658 16283 106966 16292
rect 105922 15804 106230 15813
rect 105922 15802 105928 15804
rect 105984 15802 106008 15804
rect 106064 15802 106088 15804
rect 106144 15802 106168 15804
rect 106224 15802 106230 15804
rect 105984 15750 105986 15802
rect 106166 15750 106168 15802
rect 105922 15748 105928 15750
rect 105984 15748 106008 15750
rect 106064 15748 106088 15750
rect 106144 15748 106168 15750
rect 106224 15748 106230 15750
rect 105922 15739 106230 15748
rect 106658 15260 106966 15269
rect 106658 15258 106664 15260
rect 106720 15258 106744 15260
rect 106800 15258 106824 15260
rect 106880 15258 106904 15260
rect 106960 15258 106966 15260
rect 106720 15206 106722 15258
rect 106902 15206 106904 15258
rect 106658 15204 106664 15206
rect 106720 15204 106744 15206
rect 106800 15204 106824 15206
rect 106880 15204 106904 15206
rect 106960 15204 106966 15206
rect 106658 15195 106966 15204
rect 105922 14716 106230 14725
rect 105922 14714 105928 14716
rect 105984 14714 106008 14716
rect 106064 14714 106088 14716
rect 106144 14714 106168 14716
rect 106224 14714 106230 14716
rect 105984 14662 105986 14714
rect 106166 14662 106168 14714
rect 105922 14660 105928 14662
rect 105984 14660 106008 14662
rect 106064 14660 106088 14662
rect 106144 14660 106168 14662
rect 106224 14660 106230 14662
rect 105922 14651 106230 14660
rect 106658 14172 106966 14181
rect 106658 14170 106664 14172
rect 106720 14170 106744 14172
rect 106800 14170 106824 14172
rect 106880 14170 106904 14172
rect 106960 14170 106966 14172
rect 106720 14118 106722 14170
rect 106902 14118 106904 14170
rect 106658 14116 106664 14118
rect 106720 14116 106744 14118
rect 106800 14116 106824 14118
rect 106880 14116 106904 14118
rect 106960 14116 106966 14118
rect 106658 14107 106966 14116
rect 105922 13628 106230 13637
rect 105922 13626 105928 13628
rect 105984 13626 106008 13628
rect 106064 13626 106088 13628
rect 106144 13626 106168 13628
rect 106224 13626 106230 13628
rect 105984 13574 105986 13626
rect 106166 13574 106168 13626
rect 105922 13572 105928 13574
rect 105984 13572 106008 13574
rect 106064 13572 106088 13574
rect 106144 13572 106168 13574
rect 106224 13572 106230 13574
rect 105922 13563 106230 13572
rect 106658 13084 106966 13093
rect 106658 13082 106664 13084
rect 106720 13082 106744 13084
rect 106800 13082 106824 13084
rect 106880 13082 106904 13084
rect 106960 13082 106966 13084
rect 106720 13030 106722 13082
rect 106902 13030 106904 13082
rect 106658 13028 106664 13030
rect 106720 13028 106744 13030
rect 106800 13028 106824 13030
rect 106880 13028 106904 13030
rect 106960 13028 106966 13030
rect 106658 13019 106966 13028
rect 105922 12540 106230 12549
rect 105922 12538 105928 12540
rect 105984 12538 106008 12540
rect 106064 12538 106088 12540
rect 106144 12538 106168 12540
rect 106224 12538 106230 12540
rect 105984 12486 105986 12538
rect 106166 12486 106168 12538
rect 105922 12484 105928 12486
rect 105984 12484 106008 12486
rect 106064 12484 106088 12486
rect 106144 12484 106168 12486
rect 106224 12484 106230 12486
rect 105922 12475 106230 12484
rect 106658 11996 106966 12005
rect 106658 11994 106664 11996
rect 106720 11994 106744 11996
rect 106800 11994 106824 11996
rect 106880 11994 106904 11996
rect 106960 11994 106966 11996
rect 106720 11942 106722 11994
rect 106902 11942 106904 11994
rect 106658 11940 106664 11942
rect 106720 11940 106744 11942
rect 106800 11940 106824 11942
rect 106880 11940 106904 11942
rect 106960 11940 106966 11942
rect 106658 11931 106966 11940
rect 105922 11452 106230 11461
rect 105922 11450 105928 11452
rect 105984 11450 106008 11452
rect 106064 11450 106088 11452
rect 106144 11450 106168 11452
rect 106224 11450 106230 11452
rect 105984 11398 105986 11450
rect 106166 11398 106168 11450
rect 105922 11396 105928 11398
rect 105984 11396 106008 11398
rect 106064 11396 106088 11398
rect 106144 11396 106168 11398
rect 106224 11396 106230 11398
rect 105922 11387 106230 11396
rect 106658 10908 106966 10917
rect 106658 10906 106664 10908
rect 106720 10906 106744 10908
rect 106800 10906 106824 10908
rect 106880 10906 106904 10908
rect 106960 10906 106966 10908
rect 106720 10854 106722 10906
rect 106902 10854 106904 10906
rect 106658 10852 106664 10854
rect 106720 10852 106744 10854
rect 106800 10852 106824 10854
rect 106880 10852 106904 10854
rect 106960 10852 106966 10854
rect 106658 10843 106966 10852
rect 105922 10364 106230 10373
rect 105922 10362 105928 10364
rect 105984 10362 106008 10364
rect 106064 10362 106088 10364
rect 106144 10362 106168 10364
rect 106224 10362 106230 10364
rect 105984 10310 105986 10362
rect 106166 10310 106168 10362
rect 105922 10308 105928 10310
rect 105984 10308 106008 10310
rect 106064 10308 106088 10310
rect 106144 10308 106168 10310
rect 106224 10308 106230 10310
rect 105922 10299 106230 10308
rect 106658 9820 106966 9829
rect 106658 9818 106664 9820
rect 106720 9818 106744 9820
rect 106800 9818 106824 9820
rect 106880 9818 106904 9820
rect 106960 9818 106966 9820
rect 106720 9766 106722 9818
rect 106902 9766 106904 9818
rect 106658 9764 106664 9766
rect 106720 9764 106744 9766
rect 106800 9764 106824 9766
rect 106880 9764 106904 9766
rect 106960 9764 106966 9766
rect 106658 9755 106966 9764
rect 103612 9648 103664 9654
rect 103612 9590 103664 9596
rect 103520 9580 103572 9586
rect 103520 9522 103572 9528
rect 102140 9512 102192 9518
rect 102140 9454 102192 9460
rect 105922 9276 106230 9285
rect 105922 9274 105928 9276
rect 105984 9274 106008 9276
rect 106064 9274 106088 9276
rect 106144 9274 106168 9276
rect 106224 9274 106230 9276
rect 105984 9222 105986 9274
rect 106166 9222 106168 9274
rect 105922 9220 105928 9222
rect 105984 9220 106008 9222
rect 106064 9220 106088 9222
rect 106144 9220 106168 9222
rect 106224 9220 106230 9222
rect 105922 9211 106230 9220
rect 106658 8732 106966 8741
rect 106658 8730 106664 8732
rect 106720 8730 106744 8732
rect 106800 8730 106824 8732
rect 106880 8730 106904 8732
rect 106960 8730 106966 8732
rect 106720 8678 106722 8730
rect 106902 8678 106904 8730
rect 106658 8676 106664 8678
rect 106720 8676 106744 8678
rect 106800 8676 106824 8678
rect 106880 8676 106904 8678
rect 106960 8676 106966 8678
rect 106658 8667 106966 8676
rect 105922 8188 106230 8197
rect 105922 8186 105928 8188
rect 105984 8186 106008 8188
rect 106064 8186 106088 8188
rect 106144 8186 106168 8188
rect 106224 8186 106230 8188
rect 105984 8134 105986 8186
rect 106166 8134 106168 8186
rect 105922 8132 105928 8134
rect 105984 8132 106008 8134
rect 106064 8132 106088 8134
rect 106144 8132 106168 8134
rect 106224 8132 106230 8134
rect 105922 8123 106230 8132
rect 97034 7644 97342 7653
rect 97034 7642 97040 7644
rect 97096 7642 97120 7644
rect 97176 7642 97200 7644
rect 97256 7642 97280 7644
rect 97336 7642 97342 7644
rect 97096 7590 97098 7642
rect 97278 7590 97280 7642
rect 97034 7588 97040 7590
rect 97096 7588 97120 7590
rect 97176 7588 97200 7590
rect 97256 7588 97280 7590
rect 97336 7588 97342 7590
rect 97034 7579 97342 7588
rect 106658 7644 106966 7653
rect 106658 7642 106664 7644
rect 106720 7642 106744 7644
rect 106800 7642 106824 7644
rect 106880 7642 106904 7644
rect 106960 7642 106966 7644
rect 106720 7590 106722 7642
rect 106902 7590 106904 7642
rect 106658 7588 106664 7590
rect 106720 7588 106744 7590
rect 106800 7588 106824 7590
rect 106880 7588 106904 7590
rect 106960 7588 106966 7590
rect 106658 7579 106966 7588
rect 90548 7540 90600 7546
rect 90548 7482 90600 7488
rect 90732 7540 90784 7546
rect 90732 7482 90784 7488
rect 90916 7540 90968 7546
rect 90916 7482 90968 7488
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 96374 7100 96682 7109
rect 96374 7098 96380 7100
rect 96436 7098 96460 7100
rect 96516 7098 96540 7100
rect 96596 7098 96620 7100
rect 96676 7098 96682 7100
rect 96436 7046 96438 7098
rect 96618 7046 96620 7098
rect 96374 7044 96380 7046
rect 96436 7044 96460 7046
rect 96516 7044 96540 7046
rect 96596 7044 96620 7046
rect 96676 7044 96682 7046
rect 96374 7035 96682 7044
rect 105922 7100 106230 7109
rect 105922 7098 105928 7100
rect 105984 7098 106008 7100
rect 106064 7098 106088 7100
rect 106144 7098 106168 7100
rect 106224 7098 106230 7100
rect 105984 7046 105986 7098
rect 106166 7046 106168 7098
rect 105922 7044 105928 7046
rect 105984 7044 106008 7046
rect 106064 7044 106088 7046
rect 106144 7044 106168 7046
rect 106224 7044 106230 7046
rect 105922 7035 106230 7044
rect 66314 6556 66622 6565
rect 66314 6554 66320 6556
rect 66376 6554 66400 6556
rect 66456 6554 66480 6556
rect 66536 6554 66560 6556
rect 66616 6554 66622 6556
rect 66376 6502 66378 6554
rect 66558 6502 66560 6554
rect 66314 6500 66320 6502
rect 66376 6500 66400 6502
rect 66456 6500 66480 6502
rect 66536 6500 66560 6502
rect 66616 6500 66622 6502
rect 66314 6491 66622 6500
rect 97034 6556 97342 6565
rect 97034 6554 97040 6556
rect 97096 6554 97120 6556
rect 97176 6554 97200 6556
rect 97256 6554 97280 6556
rect 97336 6554 97342 6556
rect 97096 6502 97098 6554
rect 97278 6502 97280 6554
rect 97034 6500 97040 6502
rect 97096 6500 97120 6502
rect 97176 6500 97200 6502
rect 97256 6500 97280 6502
rect 97336 6500 97342 6502
rect 97034 6491 97342 6500
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 96374 6012 96682 6021
rect 96374 6010 96380 6012
rect 96436 6010 96460 6012
rect 96516 6010 96540 6012
rect 96596 6010 96620 6012
rect 96676 6010 96682 6012
rect 96436 5958 96438 6010
rect 96618 5958 96620 6010
rect 96374 5956 96380 5958
rect 96436 5956 96460 5958
rect 96516 5956 96540 5958
rect 96596 5956 96620 5958
rect 96676 5956 96682 5958
rect 96374 5947 96682 5956
rect 66314 5468 66622 5477
rect 66314 5466 66320 5468
rect 66376 5466 66400 5468
rect 66456 5466 66480 5468
rect 66536 5466 66560 5468
rect 66616 5466 66622 5468
rect 66376 5414 66378 5466
rect 66558 5414 66560 5466
rect 66314 5412 66320 5414
rect 66376 5412 66400 5414
rect 66456 5412 66480 5414
rect 66536 5412 66560 5414
rect 66616 5412 66622 5414
rect 66314 5403 66622 5412
rect 97034 5468 97342 5477
rect 97034 5466 97040 5468
rect 97096 5466 97120 5468
rect 97176 5466 97200 5468
rect 97256 5466 97280 5468
rect 97336 5466 97342 5468
rect 97096 5414 97098 5466
rect 97278 5414 97280 5466
rect 97034 5412 97040 5414
rect 97096 5412 97120 5414
rect 97176 5412 97200 5414
rect 97256 5412 97280 5414
rect 97336 5412 97342 5414
rect 97034 5403 97342 5412
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 96374 4924 96682 4933
rect 96374 4922 96380 4924
rect 96436 4922 96460 4924
rect 96516 4922 96540 4924
rect 96596 4922 96620 4924
rect 96676 4922 96682 4924
rect 96436 4870 96438 4922
rect 96618 4870 96620 4922
rect 96374 4868 96380 4870
rect 96436 4868 96460 4870
rect 96516 4868 96540 4870
rect 96596 4868 96620 4870
rect 96676 4868 96682 4870
rect 96374 4859 96682 4868
rect 66314 4380 66622 4389
rect 66314 4378 66320 4380
rect 66376 4378 66400 4380
rect 66456 4378 66480 4380
rect 66536 4378 66560 4380
rect 66616 4378 66622 4380
rect 66376 4326 66378 4378
rect 66558 4326 66560 4378
rect 66314 4324 66320 4326
rect 66376 4324 66400 4326
rect 66456 4324 66480 4326
rect 66536 4324 66560 4326
rect 66616 4324 66622 4326
rect 66314 4315 66622 4324
rect 97034 4380 97342 4389
rect 97034 4378 97040 4380
rect 97096 4378 97120 4380
rect 97176 4378 97200 4380
rect 97256 4378 97280 4380
rect 97336 4378 97342 4380
rect 97096 4326 97098 4378
rect 97278 4326 97280 4378
rect 97034 4324 97040 4326
rect 97096 4324 97120 4326
rect 97176 4324 97200 4326
rect 97256 4324 97280 4326
rect 97336 4324 97342 4326
rect 97034 4315 97342 4324
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 96374 3836 96682 3845
rect 96374 3834 96380 3836
rect 96436 3834 96460 3836
rect 96516 3834 96540 3836
rect 96596 3834 96620 3836
rect 96676 3834 96682 3836
rect 96436 3782 96438 3834
rect 96618 3782 96620 3834
rect 96374 3780 96380 3782
rect 96436 3780 96460 3782
rect 96516 3780 96540 3782
rect 96596 3780 96620 3782
rect 96676 3780 96682 3782
rect 96374 3771 96682 3780
rect 66314 3292 66622 3301
rect 66314 3290 66320 3292
rect 66376 3290 66400 3292
rect 66456 3290 66480 3292
rect 66536 3290 66560 3292
rect 66616 3290 66622 3292
rect 66376 3238 66378 3290
rect 66558 3238 66560 3290
rect 66314 3236 66320 3238
rect 66376 3236 66400 3238
rect 66456 3236 66480 3238
rect 66536 3236 66560 3238
rect 66616 3236 66622 3238
rect 66314 3227 66622 3236
rect 97034 3292 97342 3301
rect 97034 3290 97040 3292
rect 97096 3290 97120 3292
rect 97176 3290 97200 3292
rect 97256 3290 97280 3292
rect 97336 3290 97342 3292
rect 97096 3238 97098 3290
rect 97278 3238 97280 3290
rect 97034 3236 97040 3238
rect 97096 3236 97120 3238
rect 97176 3236 97200 3238
rect 97256 3236 97280 3238
rect 97336 3236 97342 3238
rect 97034 3227 97342 3236
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 96374 2748 96682 2757
rect 96374 2746 96380 2748
rect 96436 2746 96460 2748
rect 96516 2746 96540 2748
rect 96596 2746 96620 2748
rect 96676 2746 96682 2748
rect 96436 2694 96438 2746
rect 96618 2694 96620 2746
rect 96374 2692 96380 2694
rect 96436 2692 96460 2694
rect 96516 2692 96540 2694
rect 96596 2692 96620 2694
rect 96676 2692 96682 2694
rect 96374 2683 96682 2692
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 32956 2644 33008 2650
rect 32956 2586 33008 2592
rect 34244 2644 34296 2650
rect 34244 2586 34296 2592
rect 35440 2644 35492 2650
rect 35440 2586 35492 2592
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 38752 2644 38804 2650
rect 38752 2586 38804 2592
rect 39948 2644 40000 2650
rect 39948 2586 40000 2592
rect 41328 2644 41380 2650
rect 41328 2586 41380 2592
rect 42156 2644 42208 2650
rect 42156 2586 42208 2592
rect 43444 2644 43496 2650
rect 43444 2586 43496 2592
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 39948 2304 40000 2310
rect 39948 2246 40000 2252
rect 41236 2304 41288 2310
rect 41236 2246 41288 2252
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 43168 2304 43220 2310
rect 43168 2246 43220 2252
rect 31588 800 31616 2246
rect 32876 800 32904 2246
rect 34164 800 34192 2246
rect 35452 800 35480 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 36096 800 36124 2246
rect 37384 800 37412 2246
rect 38672 800 38700 2246
rect 39960 800 39988 2246
rect 41248 800 41276 2246
rect 41892 800 41920 2246
rect 43180 800 43208 2246
rect 66314 2204 66622 2213
rect 66314 2202 66320 2204
rect 66376 2202 66400 2204
rect 66456 2202 66480 2204
rect 66536 2202 66560 2204
rect 66616 2202 66622 2204
rect 66376 2150 66378 2202
rect 66558 2150 66560 2202
rect 66314 2148 66320 2150
rect 66376 2148 66400 2150
rect 66456 2148 66480 2150
rect 66536 2148 66560 2150
rect 66616 2148 66622 2150
rect 66314 2139 66622 2148
rect 97034 2204 97342 2213
rect 97034 2202 97040 2204
rect 97096 2202 97120 2204
rect 97176 2202 97200 2204
rect 97256 2202 97280 2204
rect 97336 2202 97342 2204
rect 97096 2150 97098 2202
rect 97278 2150 97280 2202
rect 97034 2148 97040 2150
rect 97096 2148 97120 2150
rect 97176 2148 97200 2150
rect 97256 2148 97280 2150
rect 97336 2148 97342 2150
rect 97034 2139 97342 2148
rect 16118 0 16174 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 43166 0 43222 800
<< via2 >>
rect 4220 147450 4276 147452
rect 4300 147450 4356 147452
rect 4380 147450 4436 147452
rect 4460 147450 4516 147452
rect 4220 147398 4266 147450
rect 4266 147398 4276 147450
rect 4300 147398 4330 147450
rect 4330 147398 4342 147450
rect 4342 147398 4356 147450
rect 4380 147398 4394 147450
rect 4394 147398 4406 147450
rect 4406 147398 4436 147450
rect 4460 147398 4470 147450
rect 4470 147398 4516 147450
rect 4220 147396 4276 147398
rect 4300 147396 4356 147398
rect 4380 147396 4436 147398
rect 4460 147396 4516 147398
rect 34940 147450 34996 147452
rect 35020 147450 35076 147452
rect 35100 147450 35156 147452
rect 35180 147450 35236 147452
rect 34940 147398 34986 147450
rect 34986 147398 34996 147450
rect 35020 147398 35050 147450
rect 35050 147398 35062 147450
rect 35062 147398 35076 147450
rect 35100 147398 35114 147450
rect 35114 147398 35126 147450
rect 35126 147398 35156 147450
rect 35180 147398 35190 147450
rect 35190 147398 35236 147450
rect 34940 147396 34996 147398
rect 35020 147396 35076 147398
rect 35100 147396 35156 147398
rect 35180 147396 35236 147398
rect 65660 147450 65716 147452
rect 65740 147450 65796 147452
rect 65820 147450 65876 147452
rect 65900 147450 65956 147452
rect 65660 147398 65706 147450
rect 65706 147398 65716 147450
rect 65740 147398 65770 147450
rect 65770 147398 65782 147450
rect 65782 147398 65796 147450
rect 65820 147398 65834 147450
rect 65834 147398 65846 147450
rect 65846 147398 65876 147450
rect 65900 147398 65910 147450
rect 65910 147398 65956 147450
rect 65660 147396 65716 147398
rect 65740 147396 65796 147398
rect 65820 147396 65876 147398
rect 65900 147396 65956 147398
rect 96380 147450 96436 147452
rect 96460 147450 96516 147452
rect 96540 147450 96596 147452
rect 96620 147450 96676 147452
rect 96380 147398 96426 147450
rect 96426 147398 96436 147450
rect 96460 147398 96490 147450
rect 96490 147398 96502 147450
rect 96502 147398 96516 147450
rect 96540 147398 96554 147450
rect 96554 147398 96566 147450
rect 96566 147398 96596 147450
rect 96620 147398 96630 147450
rect 96630 147398 96676 147450
rect 96380 147396 96436 147398
rect 96460 147396 96516 147398
rect 96540 147396 96596 147398
rect 96620 147396 96676 147398
rect 4880 146906 4936 146908
rect 4960 146906 5016 146908
rect 5040 146906 5096 146908
rect 5120 146906 5176 146908
rect 4880 146854 4926 146906
rect 4926 146854 4936 146906
rect 4960 146854 4990 146906
rect 4990 146854 5002 146906
rect 5002 146854 5016 146906
rect 5040 146854 5054 146906
rect 5054 146854 5066 146906
rect 5066 146854 5096 146906
rect 5120 146854 5130 146906
rect 5130 146854 5176 146906
rect 4880 146852 4936 146854
rect 4960 146852 5016 146854
rect 5040 146852 5096 146854
rect 5120 146852 5176 146854
rect 35600 146906 35656 146908
rect 35680 146906 35736 146908
rect 35760 146906 35816 146908
rect 35840 146906 35896 146908
rect 35600 146854 35646 146906
rect 35646 146854 35656 146906
rect 35680 146854 35710 146906
rect 35710 146854 35722 146906
rect 35722 146854 35736 146906
rect 35760 146854 35774 146906
rect 35774 146854 35786 146906
rect 35786 146854 35816 146906
rect 35840 146854 35850 146906
rect 35850 146854 35896 146906
rect 35600 146852 35656 146854
rect 35680 146852 35736 146854
rect 35760 146852 35816 146854
rect 35840 146852 35896 146854
rect 66320 146906 66376 146908
rect 66400 146906 66456 146908
rect 66480 146906 66536 146908
rect 66560 146906 66616 146908
rect 66320 146854 66366 146906
rect 66366 146854 66376 146906
rect 66400 146854 66430 146906
rect 66430 146854 66442 146906
rect 66442 146854 66456 146906
rect 66480 146854 66494 146906
rect 66494 146854 66506 146906
rect 66506 146854 66536 146906
rect 66560 146854 66570 146906
rect 66570 146854 66616 146906
rect 66320 146852 66376 146854
rect 66400 146852 66456 146854
rect 66480 146852 66536 146854
rect 66560 146852 66616 146854
rect 97040 146906 97096 146908
rect 97120 146906 97176 146908
rect 97200 146906 97256 146908
rect 97280 146906 97336 146908
rect 97040 146854 97086 146906
rect 97086 146854 97096 146906
rect 97120 146854 97150 146906
rect 97150 146854 97162 146906
rect 97162 146854 97176 146906
rect 97200 146854 97214 146906
rect 97214 146854 97226 146906
rect 97226 146854 97256 146906
rect 97280 146854 97290 146906
rect 97290 146854 97336 146906
rect 97040 146852 97096 146854
rect 97120 146852 97176 146854
rect 97200 146852 97256 146854
rect 97280 146852 97336 146854
rect 4220 146362 4276 146364
rect 4300 146362 4356 146364
rect 4380 146362 4436 146364
rect 4460 146362 4516 146364
rect 4220 146310 4266 146362
rect 4266 146310 4276 146362
rect 4300 146310 4330 146362
rect 4330 146310 4342 146362
rect 4342 146310 4356 146362
rect 4380 146310 4394 146362
rect 4394 146310 4406 146362
rect 4406 146310 4436 146362
rect 4460 146310 4470 146362
rect 4470 146310 4516 146362
rect 4220 146308 4276 146310
rect 4300 146308 4356 146310
rect 4380 146308 4436 146310
rect 4460 146308 4516 146310
rect 34940 146362 34996 146364
rect 35020 146362 35076 146364
rect 35100 146362 35156 146364
rect 35180 146362 35236 146364
rect 34940 146310 34986 146362
rect 34986 146310 34996 146362
rect 35020 146310 35050 146362
rect 35050 146310 35062 146362
rect 35062 146310 35076 146362
rect 35100 146310 35114 146362
rect 35114 146310 35126 146362
rect 35126 146310 35156 146362
rect 35180 146310 35190 146362
rect 35190 146310 35236 146362
rect 34940 146308 34996 146310
rect 35020 146308 35076 146310
rect 35100 146308 35156 146310
rect 35180 146308 35236 146310
rect 65660 146362 65716 146364
rect 65740 146362 65796 146364
rect 65820 146362 65876 146364
rect 65900 146362 65956 146364
rect 65660 146310 65706 146362
rect 65706 146310 65716 146362
rect 65740 146310 65770 146362
rect 65770 146310 65782 146362
rect 65782 146310 65796 146362
rect 65820 146310 65834 146362
rect 65834 146310 65846 146362
rect 65846 146310 65876 146362
rect 65900 146310 65910 146362
rect 65910 146310 65956 146362
rect 65660 146308 65716 146310
rect 65740 146308 65796 146310
rect 65820 146308 65876 146310
rect 65900 146308 65956 146310
rect 96380 146362 96436 146364
rect 96460 146362 96516 146364
rect 96540 146362 96596 146364
rect 96620 146362 96676 146364
rect 96380 146310 96426 146362
rect 96426 146310 96436 146362
rect 96460 146310 96490 146362
rect 96490 146310 96502 146362
rect 96502 146310 96516 146362
rect 96540 146310 96554 146362
rect 96554 146310 96566 146362
rect 96566 146310 96596 146362
rect 96620 146310 96630 146362
rect 96630 146310 96676 146362
rect 96380 146308 96436 146310
rect 96460 146308 96516 146310
rect 96540 146308 96596 146310
rect 96620 146308 96676 146310
rect 4880 145818 4936 145820
rect 4960 145818 5016 145820
rect 5040 145818 5096 145820
rect 5120 145818 5176 145820
rect 4880 145766 4926 145818
rect 4926 145766 4936 145818
rect 4960 145766 4990 145818
rect 4990 145766 5002 145818
rect 5002 145766 5016 145818
rect 5040 145766 5054 145818
rect 5054 145766 5066 145818
rect 5066 145766 5096 145818
rect 5120 145766 5130 145818
rect 5130 145766 5176 145818
rect 4880 145764 4936 145766
rect 4960 145764 5016 145766
rect 5040 145764 5096 145766
rect 5120 145764 5176 145766
rect 35600 145818 35656 145820
rect 35680 145818 35736 145820
rect 35760 145818 35816 145820
rect 35840 145818 35896 145820
rect 35600 145766 35646 145818
rect 35646 145766 35656 145818
rect 35680 145766 35710 145818
rect 35710 145766 35722 145818
rect 35722 145766 35736 145818
rect 35760 145766 35774 145818
rect 35774 145766 35786 145818
rect 35786 145766 35816 145818
rect 35840 145766 35850 145818
rect 35850 145766 35896 145818
rect 35600 145764 35656 145766
rect 35680 145764 35736 145766
rect 35760 145764 35816 145766
rect 35840 145764 35896 145766
rect 66320 145818 66376 145820
rect 66400 145818 66456 145820
rect 66480 145818 66536 145820
rect 66560 145818 66616 145820
rect 66320 145766 66366 145818
rect 66366 145766 66376 145818
rect 66400 145766 66430 145818
rect 66430 145766 66442 145818
rect 66442 145766 66456 145818
rect 66480 145766 66494 145818
rect 66494 145766 66506 145818
rect 66506 145766 66536 145818
rect 66560 145766 66570 145818
rect 66570 145766 66616 145818
rect 66320 145764 66376 145766
rect 66400 145764 66456 145766
rect 66480 145764 66536 145766
rect 66560 145764 66616 145766
rect 97040 145818 97096 145820
rect 97120 145818 97176 145820
rect 97200 145818 97256 145820
rect 97280 145818 97336 145820
rect 97040 145766 97086 145818
rect 97086 145766 97096 145818
rect 97120 145766 97150 145818
rect 97150 145766 97162 145818
rect 97162 145766 97176 145818
rect 97200 145766 97214 145818
rect 97214 145766 97226 145818
rect 97226 145766 97256 145818
rect 97280 145766 97290 145818
rect 97290 145766 97336 145818
rect 97040 145764 97096 145766
rect 97120 145764 97176 145766
rect 97200 145764 97256 145766
rect 97280 145764 97336 145766
rect 4220 145274 4276 145276
rect 4300 145274 4356 145276
rect 4380 145274 4436 145276
rect 4460 145274 4516 145276
rect 4220 145222 4266 145274
rect 4266 145222 4276 145274
rect 4300 145222 4330 145274
rect 4330 145222 4342 145274
rect 4342 145222 4356 145274
rect 4380 145222 4394 145274
rect 4394 145222 4406 145274
rect 4406 145222 4436 145274
rect 4460 145222 4470 145274
rect 4470 145222 4516 145274
rect 4220 145220 4276 145222
rect 4300 145220 4356 145222
rect 4380 145220 4436 145222
rect 4460 145220 4516 145222
rect 34940 145274 34996 145276
rect 35020 145274 35076 145276
rect 35100 145274 35156 145276
rect 35180 145274 35236 145276
rect 34940 145222 34986 145274
rect 34986 145222 34996 145274
rect 35020 145222 35050 145274
rect 35050 145222 35062 145274
rect 35062 145222 35076 145274
rect 35100 145222 35114 145274
rect 35114 145222 35126 145274
rect 35126 145222 35156 145274
rect 35180 145222 35190 145274
rect 35190 145222 35236 145274
rect 34940 145220 34996 145222
rect 35020 145220 35076 145222
rect 35100 145220 35156 145222
rect 35180 145220 35236 145222
rect 65660 145274 65716 145276
rect 65740 145274 65796 145276
rect 65820 145274 65876 145276
rect 65900 145274 65956 145276
rect 65660 145222 65706 145274
rect 65706 145222 65716 145274
rect 65740 145222 65770 145274
rect 65770 145222 65782 145274
rect 65782 145222 65796 145274
rect 65820 145222 65834 145274
rect 65834 145222 65846 145274
rect 65846 145222 65876 145274
rect 65900 145222 65910 145274
rect 65910 145222 65956 145274
rect 65660 145220 65716 145222
rect 65740 145220 65796 145222
rect 65820 145220 65876 145222
rect 65900 145220 65956 145222
rect 96380 145274 96436 145276
rect 96460 145274 96516 145276
rect 96540 145274 96596 145276
rect 96620 145274 96676 145276
rect 96380 145222 96426 145274
rect 96426 145222 96436 145274
rect 96460 145222 96490 145274
rect 96490 145222 96502 145274
rect 96502 145222 96516 145274
rect 96540 145222 96554 145274
rect 96554 145222 96566 145274
rect 96566 145222 96596 145274
rect 96620 145222 96630 145274
rect 96630 145222 96676 145274
rect 96380 145220 96436 145222
rect 96460 145220 96516 145222
rect 96540 145220 96596 145222
rect 96620 145220 96676 145222
rect 4880 144730 4936 144732
rect 4960 144730 5016 144732
rect 5040 144730 5096 144732
rect 5120 144730 5176 144732
rect 4880 144678 4926 144730
rect 4926 144678 4936 144730
rect 4960 144678 4990 144730
rect 4990 144678 5002 144730
rect 5002 144678 5016 144730
rect 5040 144678 5054 144730
rect 5054 144678 5066 144730
rect 5066 144678 5096 144730
rect 5120 144678 5130 144730
rect 5130 144678 5176 144730
rect 4880 144676 4936 144678
rect 4960 144676 5016 144678
rect 5040 144676 5096 144678
rect 5120 144676 5176 144678
rect 35600 144730 35656 144732
rect 35680 144730 35736 144732
rect 35760 144730 35816 144732
rect 35840 144730 35896 144732
rect 35600 144678 35646 144730
rect 35646 144678 35656 144730
rect 35680 144678 35710 144730
rect 35710 144678 35722 144730
rect 35722 144678 35736 144730
rect 35760 144678 35774 144730
rect 35774 144678 35786 144730
rect 35786 144678 35816 144730
rect 35840 144678 35850 144730
rect 35850 144678 35896 144730
rect 35600 144676 35656 144678
rect 35680 144676 35736 144678
rect 35760 144676 35816 144678
rect 35840 144676 35896 144678
rect 66320 144730 66376 144732
rect 66400 144730 66456 144732
rect 66480 144730 66536 144732
rect 66560 144730 66616 144732
rect 66320 144678 66366 144730
rect 66366 144678 66376 144730
rect 66400 144678 66430 144730
rect 66430 144678 66442 144730
rect 66442 144678 66456 144730
rect 66480 144678 66494 144730
rect 66494 144678 66506 144730
rect 66506 144678 66536 144730
rect 66560 144678 66570 144730
rect 66570 144678 66616 144730
rect 66320 144676 66376 144678
rect 66400 144676 66456 144678
rect 66480 144676 66536 144678
rect 66560 144676 66616 144678
rect 97040 144730 97096 144732
rect 97120 144730 97176 144732
rect 97200 144730 97256 144732
rect 97280 144730 97336 144732
rect 97040 144678 97086 144730
rect 97086 144678 97096 144730
rect 97120 144678 97150 144730
rect 97150 144678 97162 144730
rect 97162 144678 97176 144730
rect 97200 144678 97214 144730
rect 97214 144678 97226 144730
rect 97226 144678 97256 144730
rect 97280 144678 97290 144730
rect 97290 144678 97336 144730
rect 97040 144676 97096 144678
rect 97120 144676 97176 144678
rect 97200 144676 97256 144678
rect 97280 144676 97336 144678
rect 4220 144186 4276 144188
rect 4300 144186 4356 144188
rect 4380 144186 4436 144188
rect 4460 144186 4516 144188
rect 4220 144134 4266 144186
rect 4266 144134 4276 144186
rect 4300 144134 4330 144186
rect 4330 144134 4342 144186
rect 4342 144134 4356 144186
rect 4380 144134 4394 144186
rect 4394 144134 4406 144186
rect 4406 144134 4436 144186
rect 4460 144134 4470 144186
rect 4470 144134 4516 144186
rect 4220 144132 4276 144134
rect 4300 144132 4356 144134
rect 4380 144132 4436 144134
rect 4460 144132 4516 144134
rect 34940 144186 34996 144188
rect 35020 144186 35076 144188
rect 35100 144186 35156 144188
rect 35180 144186 35236 144188
rect 34940 144134 34986 144186
rect 34986 144134 34996 144186
rect 35020 144134 35050 144186
rect 35050 144134 35062 144186
rect 35062 144134 35076 144186
rect 35100 144134 35114 144186
rect 35114 144134 35126 144186
rect 35126 144134 35156 144186
rect 35180 144134 35190 144186
rect 35190 144134 35236 144186
rect 34940 144132 34996 144134
rect 35020 144132 35076 144134
rect 35100 144132 35156 144134
rect 35180 144132 35236 144134
rect 65660 144186 65716 144188
rect 65740 144186 65796 144188
rect 65820 144186 65876 144188
rect 65900 144186 65956 144188
rect 65660 144134 65706 144186
rect 65706 144134 65716 144186
rect 65740 144134 65770 144186
rect 65770 144134 65782 144186
rect 65782 144134 65796 144186
rect 65820 144134 65834 144186
rect 65834 144134 65846 144186
rect 65846 144134 65876 144186
rect 65900 144134 65910 144186
rect 65910 144134 65956 144186
rect 65660 144132 65716 144134
rect 65740 144132 65796 144134
rect 65820 144132 65876 144134
rect 65900 144132 65956 144134
rect 96380 144186 96436 144188
rect 96460 144186 96516 144188
rect 96540 144186 96596 144188
rect 96620 144186 96676 144188
rect 96380 144134 96426 144186
rect 96426 144134 96436 144186
rect 96460 144134 96490 144186
rect 96490 144134 96502 144186
rect 96502 144134 96516 144186
rect 96540 144134 96554 144186
rect 96554 144134 96566 144186
rect 96566 144134 96596 144186
rect 96620 144134 96630 144186
rect 96630 144134 96676 144186
rect 96380 144132 96436 144134
rect 96460 144132 96516 144134
rect 96540 144132 96596 144134
rect 96620 144132 96676 144134
rect 4880 143642 4936 143644
rect 4960 143642 5016 143644
rect 5040 143642 5096 143644
rect 5120 143642 5176 143644
rect 4880 143590 4926 143642
rect 4926 143590 4936 143642
rect 4960 143590 4990 143642
rect 4990 143590 5002 143642
rect 5002 143590 5016 143642
rect 5040 143590 5054 143642
rect 5054 143590 5066 143642
rect 5066 143590 5096 143642
rect 5120 143590 5130 143642
rect 5130 143590 5176 143642
rect 4880 143588 4936 143590
rect 4960 143588 5016 143590
rect 5040 143588 5096 143590
rect 5120 143588 5176 143590
rect 35600 143642 35656 143644
rect 35680 143642 35736 143644
rect 35760 143642 35816 143644
rect 35840 143642 35896 143644
rect 35600 143590 35646 143642
rect 35646 143590 35656 143642
rect 35680 143590 35710 143642
rect 35710 143590 35722 143642
rect 35722 143590 35736 143642
rect 35760 143590 35774 143642
rect 35774 143590 35786 143642
rect 35786 143590 35816 143642
rect 35840 143590 35850 143642
rect 35850 143590 35896 143642
rect 35600 143588 35656 143590
rect 35680 143588 35736 143590
rect 35760 143588 35816 143590
rect 35840 143588 35896 143590
rect 66320 143642 66376 143644
rect 66400 143642 66456 143644
rect 66480 143642 66536 143644
rect 66560 143642 66616 143644
rect 66320 143590 66366 143642
rect 66366 143590 66376 143642
rect 66400 143590 66430 143642
rect 66430 143590 66442 143642
rect 66442 143590 66456 143642
rect 66480 143590 66494 143642
rect 66494 143590 66506 143642
rect 66506 143590 66536 143642
rect 66560 143590 66570 143642
rect 66570 143590 66616 143642
rect 66320 143588 66376 143590
rect 66400 143588 66456 143590
rect 66480 143588 66536 143590
rect 66560 143588 66616 143590
rect 97040 143642 97096 143644
rect 97120 143642 97176 143644
rect 97200 143642 97256 143644
rect 97280 143642 97336 143644
rect 97040 143590 97086 143642
rect 97086 143590 97096 143642
rect 97120 143590 97150 143642
rect 97150 143590 97162 143642
rect 97162 143590 97176 143642
rect 97200 143590 97214 143642
rect 97214 143590 97226 143642
rect 97226 143590 97256 143642
rect 97280 143590 97290 143642
rect 97290 143590 97336 143642
rect 97040 143588 97096 143590
rect 97120 143588 97176 143590
rect 97200 143588 97256 143590
rect 97280 143588 97336 143590
rect 4220 143098 4276 143100
rect 4300 143098 4356 143100
rect 4380 143098 4436 143100
rect 4460 143098 4516 143100
rect 4220 143046 4266 143098
rect 4266 143046 4276 143098
rect 4300 143046 4330 143098
rect 4330 143046 4342 143098
rect 4342 143046 4356 143098
rect 4380 143046 4394 143098
rect 4394 143046 4406 143098
rect 4406 143046 4436 143098
rect 4460 143046 4470 143098
rect 4470 143046 4516 143098
rect 4220 143044 4276 143046
rect 4300 143044 4356 143046
rect 4380 143044 4436 143046
rect 4460 143044 4516 143046
rect 34940 143098 34996 143100
rect 35020 143098 35076 143100
rect 35100 143098 35156 143100
rect 35180 143098 35236 143100
rect 34940 143046 34986 143098
rect 34986 143046 34996 143098
rect 35020 143046 35050 143098
rect 35050 143046 35062 143098
rect 35062 143046 35076 143098
rect 35100 143046 35114 143098
rect 35114 143046 35126 143098
rect 35126 143046 35156 143098
rect 35180 143046 35190 143098
rect 35190 143046 35236 143098
rect 34940 143044 34996 143046
rect 35020 143044 35076 143046
rect 35100 143044 35156 143046
rect 35180 143044 35236 143046
rect 65660 143098 65716 143100
rect 65740 143098 65796 143100
rect 65820 143098 65876 143100
rect 65900 143098 65956 143100
rect 65660 143046 65706 143098
rect 65706 143046 65716 143098
rect 65740 143046 65770 143098
rect 65770 143046 65782 143098
rect 65782 143046 65796 143098
rect 65820 143046 65834 143098
rect 65834 143046 65846 143098
rect 65846 143046 65876 143098
rect 65900 143046 65910 143098
rect 65910 143046 65956 143098
rect 65660 143044 65716 143046
rect 65740 143044 65796 143046
rect 65820 143044 65876 143046
rect 65900 143044 65956 143046
rect 96380 143098 96436 143100
rect 96460 143098 96516 143100
rect 96540 143098 96596 143100
rect 96620 143098 96676 143100
rect 96380 143046 96426 143098
rect 96426 143046 96436 143098
rect 96460 143046 96490 143098
rect 96490 143046 96502 143098
rect 96502 143046 96516 143098
rect 96540 143046 96554 143098
rect 96554 143046 96566 143098
rect 96566 143046 96596 143098
rect 96620 143046 96630 143098
rect 96630 143046 96676 143098
rect 96380 143044 96436 143046
rect 96460 143044 96516 143046
rect 96540 143044 96596 143046
rect 96620 143044 96676 143046
rect 4880 142554 4936 142556
rect 4960 142554 5016 142556
rect 5040 142554 5096 142556
rect 5120 142554 5176 142556
rect 4880 142502 4926 142554
rect 4926 142502 4936 142554
rect 4960 142502 4990 142554
rect 4990 142502 5002 142554
rect 5002 142502 5016 142554
rect 5040 142502 5054 142554
rect 5054 142502 5066 142554
rect 5066 142502 5096 142554
rect 5120 142502 5130 142554
rect 5130 142502 5176 142554
rect 4880 142500 4936 142502
rect 4960 142500 5016 142502
rect 5040 142500 5096 142502
rect 5120 142500 5176 142502
rect 35600 142554 35656 142556
rect 35680 142554 35736 142556
rect 35760 142554 35816 142556
rect 35840 142554 35896 142556
rect 35600 142502 35646 142554
rect 35646 142502 35656 142554
rect 35680 142502 35710 142554
rect 35710 142502 35722 142554
rect 35722 142502 35736 142554
rect 35760 142502 35774 142554
rect 35774 142502 35786 142554
rect 35786 142502 35816 142554
rect 35840 142502 35850 142554
rect 35850 142502 35896 142554
rect 35600 142500 35656 142502
rect 35680 142500 35736 142502
rect 35760 142500 35816 142502
rect 35840 142500 35896 142502
rect 66320 142554 66376 142556
rect 66400 142554 66456 142556
rect 66480 142554 66536 142556
rect 66560 142554 66616 142556
rect 66320 142502 66366 142554
rect 66366 142502 66376 142554
rect 66400 142502 66430 142554
rect 66430 142502 66442 142554
rect 66442 142502 66456 142554
rect 66480 142502 66494 142554
rect 66494 142502 66506 142554
rect 66506 142502 66536 142554
rect 66560 142502 66570 142554
rect 66570 142502 66616 142554
rect 66320 142500 66376 142502
rect 66400 142500 66456 142502
rect 66480 142500 66536 142502
rect 66560 142500 66616 142502
rect 97040 142554 97096 142556
rect 97120 142554 97176 142556
rect 97200 142554 97256 142556
rect 97280 142554 97336 142556
rect 97040 142502 97086 142554
rect 97086 142502 97096 142554
rect 97120 142502 97150 142554
rect 97150 142502 97162 142554
rect 97162 142502 97176 142554
rect 97200 142502 97214 142554
rect 97214 142502 97226 142554
rect 97226 142502 97256 142554
rect 97280 142502 97290 142554
rect 97290 142502 97336 142554
rect 97040 142500 97096 142502
rect 97120 142500 97176 142502
rect 97200 142500 97256 142502
rect 97280 142500 97336 142502
rect 4220 142010 4276 142012
rect 4300 142010 4356 142012
rect 4380 142010 4436 142012
rect 4460 142010 4516 142012
rect 4220 141958 4266 142010
rect 4266 141958 4276 142010
rect 4300 141958 4330 142010
rect 4330 141958 4342 142010
rect 4342 141958 4356 142010
rect 4380 141958 4394 142010
rect 4394 141958 4406 142010
rect 4406 141958 4436 142010
rect 4460 141958 4470 142010
rect 4470 141958 4516 142010
rect 4220 141956 4276 141958
rect 4300 141956 4356 141958
rect 4380 141956 4436 141958
rect 4460 141956 4516 141958
rect 34940 142010 34996 142012
rect 35020 142010 35076 142012
rect 35100 142010 35156 142012
rect 35180 142010 35236 142012
rect 34940 141958 34986 142010
rect 34986 141958 34996 142010
rect 35020 141958 35050 142010
rect 35050 141958 35062 142010
rect 35062 141958 35076 142010
rect 35100 141958 35114 142010
rect 35114 141958 35126 142010
rect 35126 141958 35156 142010
rect 35180 141958 35190 142010
rect 35190 141958 35236 142010
rect 34940 141956 34996 141958
rect 35020 141956 35076 141958
rect 35100 141956 35156 141958
rect 35180 141956 35236 141958
rect 65660 142010 65716 142012
rect 65740 142010 65796 142012
rect 65820 142010 65876 142012
rect 65900 142010 65956 142012
rect 65660 141958 65706 142010
rect 65706 141958 65716 142010
rect 65740 141958 65770 142010
rect 65770 141958 65782 142010
rect 65782 141958 65796 142010
rect 65820 141958 65834 142010
rect 65834 141958 65846 142010
rect 65846 141958 65876 142010
rect 65900 141958 65910 142010
rect 65910 141958 65956 142010
rect 65660 141956 65716 141958
rect 65740 141956 65796 141958
rect 65820 141956 65876 141958
rect 65900 141956 65956 141958
rect 96380 142010 96436 142012
rect 96460 142010 96516 142012
rect 96540 142010 96596 142012
rect 96620 142010 96676 142012
rect 96380 141958 96426 142010
rect 96426 141958 96436 142010
rect 96460 141958 96490 142010
rect 96490 141958 96502 142010
rect 96502 141958 96516 142010
rect 96540 141958 96554 142010
rect 96554 141958 96566 142010
rect 96566 141958 96596 142010
rect 96620 141958 96630 142010
rect 96630 141958 96676 142010
rect 96380 141956 96436 141958
rect 96460 141956 96516 141958
rect 96540 141956 96596 141958
rect 96620 141956 96676 141958
rect 4880 141466 4936 141468
rect 4960 141466 5016 141468
rect 5040 141466 5096 141468
rect 5120 141466 5176 141468
rect 4880 141414 4926 141466
rect 4926 141414 4936 141466
rect 4960 141414 4990 141466
rect 4990 141414 5002 141466
rect 5002 141414 5016 141466
rect 5040 141414 5054 141466
rect 5054 141414 5066 141466
rect 5066 141414 5096 141466
rect 5120 141414 5130 141466
rect 5130 141414 5176 141466
rect 4880 141412 4936 141414
rect 4960 141412 5016 141414
rect 5040 141412 5096 141414
rect 5120 141412 5176 141414
rect 35600 141466 35656 141468
rect 35680 141466 35736 141468
rect 35760 141466 35816 141468
rect 35840 141466 35896 141468
rect 35600 141414 35646 141466
rect 35646 141414 35656 141466
rect 35680 141414 35710 141466
rect 35710 141414 35722 141466
rect 35722 141414 35736 141466
rect 35760 141414 35774 141466
rect 35774 141414 35786 141466
rect 35786 141414 35816 141466
rect 35840 141414 35850 141466
rect 35850 141414 35896 141466
rect 35600 141412 35656 141414
rect 35680 141412 35736 141414
rect 35760 141412 35816 141414
rect 35840 141412 35896 141414
rect 66320 141466 66376 141468
rect 66400 141466 66456 141468
rect 66480 141466 66536 141468
rect 66560 141466 66616 141468
rect 66320 141414 66366 141466
rect 66366 141414 66376 141466
rect 66400 141414 66430 141466
rect 66430 141414 66442 141466
rect 66442 141414 66456 141466
rect 66480 141414 66494 141466
rect 66494 141414 66506 141466
rect 66506 141414 66536 141466
rect 66560 141414 66570 141466
rect 66570 141414 66616 141466
rect 66320 141412 66376 141414
rect 66400 141412 66456 141414
rect 66480 141412 66536 141414
rect 66560 141412 66616 141414
rect 97040 141466 97096 141468
rect 97120 141466 97176 141468
rect 97200 141466 97256 141468
rect 97280 141466 97336 141468
rect 97040 141414 97086 141466
rect 97086 141414 97096 141466
rect 97120 141414 97150 141466
rect 97150 141414 97162 141466
rect 97162 141414 97176 141466
rect 97200 141414 97214 141466
rect 97214 141414 97226 141466
rect 97226 141414 97256 141466
rect 97280 141414 97290 141466
rect 97290 141414 97336 141466
rect 97040 141412 97096 141414
rect 97120 141412 97176 141414
rect 97200 141412 97256 141414
rect 97280 141412 97336 141414
rect 4220 140922 4276 140924
rect 4300 140922 4356 140924
rect 4380 140922 4436 140924
rect 4460 140922 4516 140924
rect 4220 140870 4266 140922
rect 4266 140870 4276 140922
rect 4300 140870 4330 140922
rect 4330 140870 4342 140922
rect 4342 140870 4356 140922
rect 4380 140870 4394 140922
rect 4394 140870 4406 140922
rect 4406 140870 4436 140922
rect 4460 140870 4470 140922
rect 4470 140870 4516 140922
rect 4220 140868 4276 140870
rect 4300 140868 4356 140870
rect 4380 140868 4436 140870
rect 4460 140868 4516 140870
rect 34940 140922 34996 140924
rect 35020 140922 35076 140924
rect 35100 140922 35156 140924
rect 35180 140922 35236 140924
rect 34940 140870 34986 140922
rect 34986 140870 34996 140922
rect 35020 140870 35050 140922
rect 35050 140870 35062 140922
rect 35062 140870 35076 140922
rect 35100 140870 35114 140922
rect 35114 140870 35126 140922
rect 35126 140870 35156 140922
rect 35180 140870 35190 140922
rect 35190 140870 35236 140922
rect 34940 140868 34996 140870
rect 35020 140868 35076 140870
rect 35100 140868 35156 140870
rect 35180 140868 35236 140870
rect 65660 140922 65716 140924
rect 65740 140922 65796 140924
rect 65820 140922 65876 140924
rect 65900 140922 65956 140924
rect 65660 140870 65706 140922
rect 65706 140870 65716 140922
rect 65740 140870 65770 140922
rect 65770 140870 65782 140922
rect 65782 140870 65796 140922
rect 65820 140870 65834 140922
rect 65834 140870 65846 140922
rect 65846 140870 65876 140922
rect 65900 140870 65910 140922
rect 65910 140870 65956 140922
rect 65660 140868 65716 140870
rect 65740 140868 65796 140870
rect 65820 140868 65876 140870
rect 65900 140868 65956 140870
rect 96380 140922 96436 140924
rect 96460 140922 96516 140924
rect 96540 140922 96596 140924
rect 96620 140922 96676 140924
rect 96380 140870 96426 140922
rect 96426 140870 96436 140922
rect 96460 140870 96490 140922
rect 96490 140870 96502 140922
rect 96502 140870 96516 140922
rect 96540 140870 96554 140922
rect 96554 140870 96566 140922
rect 96566 140870 96596 140922
rect 96620 140870 96630 140922
rect 96630 140870 96676 140922
rect 96380 140868 96436 140870
rect 96460 140868 96516 140870
rect 96540 140868 96596 140870
rect 96620 140868 96676 140870
rect 4880 140378 4936 140380
rect 4960 140378 5016 140380
rect 5040 140378 5096 140380
rect 5120 140378 5176 140380
rect 4880 140326 4926 140378
rect 4926 140326 4936 140378
rect 4960 140326 4990 140378
rect 4990 140326 5002 140378
rect 5002 140326 5016 140378
rect 5040 140326 5054 140378
rect 5054 140326 5066 140378
rect 5066 140326 5096 140378
rect 5120 140326 5130 140378
rect 5130 140326 5176 140378
rect 4880 140324 4936 140326
rect 4960 140324 5016 140326
rect 5040 140324 5096 140326
rect 5120 140324 5176 140326
rect 35600 140378 35656 140380
rect 35680 140378 35736 140380
rect 35760 140378 35816 140380
rect 35840 140378 35896 140380
rect 35600 140326 35646 140378
rect 35646 140326 35656 140378
rect 35680 140326 35710 140378
rect 35710 140326 35722 140378
rect 35722 140326 35736 140378
rect 35760 140326 35774 140378
rect 35774 140326 35786 140378
rect 35786 140326 35816 140378
rect 35840 140326 35850 140378
rect 35850 140326 35896 140378
rect 35600 140324 35656 140326
rect 35680 140324 35736 140326
rect 35760 140324 35816 140326
rect 35840 140324 35896 140326
rect 66320 140378 66376 140380
rect 66400 140378 66456 140380
rect 66480 140378 66536 140380
rect 66560 140378 66616 140380
rect 66320 140326 66366 140378
rect 66366 140326 66376 140378
rect 66400 140326 66430 140378
rect 66430 140326 66442 140378
rect 66442 140326 66456 140378
rect 66480 140326 66494 140378
rect 66494 140326 66506 140378
rect 66506 140326 66536 140378
rect 66560 140326 66570 140378
rect 66570 140326 66616 140378
rect 66320 140324 66376 140326
rect 66400 140324 66456 140326
rect 66480 140324 66536 140326
rect 66560 140324 66616 140326
rect 97040 140378 97096 140380
rect 97120 140378 97176 140380
rect 97200 140378 97256 140380
rect 97280 140378 97336 140380
rect 97040 140326 97086 140378
rect 97086 140326 97096 140378
rect 97120 140326 97150 140378
rect 97150 140326 97162 140378
rect 97162 140326 97176 140378
rect 97200 140326 97214 140378
rect 97214 140326 97226 140378
rect 97226 140326 97256 140378
rect 97280 140326 97290 140378
rect 97290 140326 97336 140378
rect 97040 140324 97096 140326
rect 97120 140324 97176 140326
rect 97200 140324 97256 140326
rect 97280 140324 97336 140326
rect 4220 139834 4276 139836
rect 4300 139834 4356 139836
rect 4380 139834 4436 139836
rect 4460 139834 4516 139836
rect 4220 139782 4266 139834
rect 4266 139782 4276 139834
rect 4300 139782 4330 139834
rect 4330 139782 4342 139834
rect 4342 139782 4356 139834
rect 4380 139782 4394 139834
rect 4394 139782 4406 139834
rect 4406 139782 4436 139834
rect 4460 139782 4470 139834
rect 4470 139782 4516 139834
rect 4220 139780 4276 139782
rect 4300 139780 4356 139782
rect 4380 139780 4436 139782
rect 4460 139780 4516 139782
rect 34940 139834 34996 139836
rect 35020 139834 35076 139836
rect 35100 139834 35156 139836
rect 35180 139834 35236 139836
rect 34940 139782 34986 139834
rect 34986 139782 34996 139834
rect 35020 139782 35050 139834
rect 35050 139782 35062 139834
rect 35062 139782 35076 139834
rect 35100 139782 35114 139834
rect 35114 139782 35126 139834
rect 35126 139782 35156 139834
rect 35180 139782 35190 139834
rect 35190 139782 35236 139834
rect 34940 139780 34996 139782
rect 35020 139780 35076 139782
rect 35100 139780 35156 139782
rect 35180 139780 35236 139782
rect 65660 139834 65716 139836
rect 65740 139834 65796 139836
rect 65820 139834 65876 139836
rect 65900 139834 65956 139836
rect 65660 139782 65706 139834
rect 65706 139782 65716 139834
rect 65740 139782 65770 139834
rect 65770 139782 65782 139834
rect 65782 139782 65796 139834
rect 65820 139782 65834 139834
rect 65834 139782 65846 139834
rect 65846 139782 65876 139834
rect 65900 139782 65910 139834
rect 65910 139782 65956 139834
rect 65660 139780 65716 139782
rect 65740 139780 65796 139782
rect 65820 139780 65876 139782
rect 65900 139780 65956 139782
rect 96380 139834 96436 139836
rect 96460 139834 96516 139836
rect 96540 139834 96596 139836
rect 96620 139834 96676 139836
rect 96380 139782 96426 139834
rect 96426 139782 96436 139834
rect 96460 139782 96490 139834
rect 96490 139782 96502 139834
rect 96502 139782 96516 139834
rect 96540 139782 96554 139834
rect 96554 139782 96566 139834
rect 96566 139782 96596 139834
rect 96620 139782 96630 139834
rect 96630 139782 96676 139834
rect 96380 139780 96436 139782
rect 96460 139780 96516 139782
rect 96540 139780 96596 139782
rect 96620 139780 96676 139782
rect 4880 139290 4936 139292
rect 4960 139290 5016 139292
rect 5040 139290 5096 139292
rect 5120 139290 5176 139292
rect 4880 139238 4926 139290
rect 4926 139238 4936 139290
rect 4960 139238 4990 139290
rect 4990 139238 5002 139290
rect 5002 139238 5016 139290
rect 5040 139238 5054 139290
rect 5054 139238 5066 139290
rect 5066 139238 5096 139290
rect 5120 139238 5130 139290
rect 5130 139238 5176 139290
rect 4880 139236 4936 139238
rect 4960 139236 5016 139238
rect 5040 139236 5096 139238
rect 5120 139236 5176 139238
rect 35600 139290 35656 139292
rect 35680 139290 35736 139292
rect 35760 139290 35816 139292
rect 35840 139290 35896 139292
rect 35600 139238 35646 139290
rect 35646 139238 35656 139290
rect 35680 139238 35710 139290
rect 35710 139238 35722 139290
rect 35722 139238 35736 139290
rect 35760 139238 35774 139290
rect 35774 139238 35786 139290
rect 35786 139238 35816 139290
rect 35840 139238 35850 139290
rect 35850 139238 35896 139290
rect 35600 139236 35656 139238
rect 35680 139236 35736 139238
rect 35760 139236 35816 139238
rect 35840 139236 35896 139238
rect 66320 139290 66376 139292
rect 66400 139290 66456 139292
rect 66480 139290 66536 139292
rect 66560 139290 66616 139292
rect 66320 139238 66366 139290
rect 66366 139238 66376 139290
rect 66400 139238 66430 139290
rect 66430 139238 66442 139290
rect 66442 139238 66456 139290
rect 66480 139238 66494 139290
rect 66494 139238 66506 139290
rect 66506 139238 66536 139290
rect 66560 139238 66570 139290
rect 66570 139238 66616 139290
rect 66320 139236 66376 139238
rect 66400 139236 66456 139238
rect 66480 139236 66536 139238
rect 66560 139236 66616 139238
rect 97040 139290 97096 139292
rect 97120 139290 97176 139292
rect 97200 139290 97256 139292
rect 97280 139290 97336 139292
rect 97040 139238 97086 139290
rect 97086 139238 97096 139290
rect 97120 139238 97150 139290
rect 97150 139238 97162 139290
rect 97162 139238 97176 139290
rect 97200 139238 97214 139290
rect 97214 139238 97226 139290
rect 97226 139238 97256 139290
rect 97280 139238 97290 139290
rect 97290 139238 97336 139290
rect 97040 139236 97096 139238
rect 97120 139236 97176 139238
rect 97200 139236 97256 139238
rect 97280 139236 97336 139238
rect 4220 138746 4276 138748
rect 4300 138746 4356 138748
rect 4380 138746 4436 138748
rect 4460 138746 4516 138748
rect 4220 138694 4266 138746
rect 4266 138694 4276 138746
rect 4300 138694 4330 138746
rect 4330 138694 4342 138746
rect 4342 138694 4356 138746
rect 4380 138694 4394 138746
rect 4394 138694 4406 138746
rect 4406 138694 4436 138746
rect 4460 138694 4470 138746
rect 4470 138694 4516 138746
rect 4220 138692 4276 138694
rect 4300 138692 4356 138694
rect 4380 138692 4436 138694
rect 4460 138692 4516 138694
rect 34940 138746 34996 138748
rect 35020 138746 35076 138748
rect 35100 138746 35156 138748
rect 35180 138746 35236 138748
rect 34940 138694 34986 138746
rect 34986 138694 34996 138746
rect 35020 138694 35050 138746
rect 35050 138694 35062 138746
rect 35062 138694 35076 138746
rect 35100 138694 35114 138746
rect 35114 138694 35126 138746
rect 35126 138694 35156 138746
rect 35180 138694 35190 138746
rect 35190 138694 35236 138746
rect 34940 138692 34996 138694
rect 35020 138692 35076 138694
rect 35100 138692 35156 138694
rect 35180 138692 35236 138694
rect 65660 138746 65716 138748
rect 65740 138746 65796 138748
rect 65820 138746 65876 138748
rect 65900 138746 65956 138748
rect 65660 138694 65706 138746
rect 65706 138694 65716 138746
rect 65740 138694 65770 138746
rect 65770 138694 65782 138746
rect 65782 138694 65796 138746
rect 65820 138694 65834 138746
rect 65834 138694 65846 138746
rect 65846 138694 65876 138746
rect 65900 138694 65910 138746
rect 65910 138694 65956 138746
rect 65660 138692 65716 138694
rect 65740 138692 65796 138694
rect 65820 138692 65876 138694
rect 65900 138692 65956 138694
rect 96380 138746 96436 138748
rect 96460 138746 96516 138748
rect 96540 138746 96596 138748
rect 96620 138746 96676 138748
rect 96380 138694 96426 138746
rect 96426 138694 96436 138746
rect 96460 138694 96490 138746
rect 96490 138694 96502 138746
rect 96502 138694 96516 138746
rect 96540 138694 96554 138746
rect 96554 138694 96566 138746
rect 96566 138694 96596 138746
rect 96620 138694 96630 138746
rect 96630 138694 96676 138746
rect 96380 138692 96436 138694
rect 96460 138692 96516 138694
rect 96540 138692 96596 138694
rect 96620 138692 96676 138694
rect 4880 138202 4936 138204
rect 4960 138202 5016 138204
rect 5040 138202 5096 138204
rect 5120 138202 5176 138204
rect 4880 138150 4926 138202
rect 4926 138150 4936 138202
rect 4960 138150 4990 138202
rect 4990 138150 5002 138202
rect 5002 138150 5016 138202
rect 5040 138150 5054 138202
rect 5054 138150 5066 138202
rect 5066 138150 5096 138202
rect 5120 138150 5130 138202
rect 5130 138150 5176 138202
rect 4880 138148 4936 138150
rect 4960 138148 5016 138150
rect 5040 138148 5096 138150
rect 5120 138148 5176 138150
rect 35600 138202 35656 138204
rect 35680 138202 35736 138204
rect 35760 138202 35816 138204
rect 35840 138202 35896 138204
rect 35600 138150 35646 138202
rect 35646 138150 35656 138202
rect 35680 138150 35710 138202
rect 35710 138150 35722 138202
rect 35722 138150 35736 138202
rect 35760 138150 35774 138202
rect 35774 138150 35786 138202
rect 35786 138150 35816 138202
rect 35840 138150 35850 138202
rect 35850 138150 35896 138202
rect 35600 138148 35656 138150
rect 35680 138148 35736 138150
rect 35760 138148 35816 138150
rect 35840 138148 35896 138150
rect 66320 138202 66376 138204
rect 66400 138202 66456 138204
rect 66480 138202 66536 138204
rect 66560 138202 66616 138204
rect 66320 138150 66366 138202
rect 66366 138150 66376 138202
rect 66400 138150 66430 138202
rect 66430 138150 66442 138202
rect 66442 138150 66456 138202
rect 66480 138150 66494 138202
rect 66494 138150 66506 138202
rect 66506 138150 66536 138202
rect 66560 138150 66570 138202
rect 66570 138150 66616 138202
rect 66320 138148 66376 138150
rect 66400 138148 66456 138150
rect 66480 138148 66536 138150
rect 66560 138148 66616 138150
rect 97040 138202 97096 138204
rect 97120 138202 97176 138204
rect 97200 138202 97256 138204
rect 97280 138202 97336 138204
rect 97040 138150 97086 138202
rect 97086 138150 97096 138202
rect 97120 138150 97150 138202
rect 97150 138150 97162 138202
rect 97162 138150 97176 138202
rect 97200 138150 97214 138202
rect 97214 138150 97226 138202
rect 97226 138150 97256 138202
rect 97280 138150 97290 138202
rect 97290 138150 97336 138202
rect 97040 138148 97096 138150
rect 97120 138148 97176 138150
rect 97200 138148 97256 138150
rect 97280 138148 97336 138150
rect 4220 137658 4276 137660
rect 4300 137658 4356 137660
rect 4380 137658 4436 137660
rect 4460 137658 4516 137660
rect 4220 137606 4266 137658
rect 4266 137606 4276 137658
rect 4300 137606 4330 137658
rect 4330 137606 4342 137658
rect 4342 137606 4356 137658
rect 4380 137606 4394 137658
rect 4394 137606 4406 137658
rect 4406 137606 4436 137658
rect 4460 137606 4470 137658
rect 4470 137606 4516 137658
rect 4220 137604 4276 137606
rect 4300 137604 4356 137606
rect 4380 137604 4436 137606
rect 4460 137604 4516 137606
rect 34940 137658 34996 137660
rect 35020 137658 35076 137660
rect 35100 137658 35156 137660
rect 35180 137658 35236 137660
rect 34940 137606 34986 137658
rect 34986 137606 34996 137658
rect 35020 137606 35050 137658
rect 35050 137606 35062 137658
rect 35062 137606 35076 137658
rect 35100 137606 35114 137658
rect 35114 137606 35126 137658
rect 35126 137606 35156 137658
rect 35180 137606 35190 137658
rect 35190 137606 35236 137658
rect 34940 137604 34996 137606
rect 35020 137604 35076 137606
rect 35100 137604 35156 137606
rect 35180 137604 35236 137606
rect 65660 137658 65716 137660
rect 65740 137658 65796 137660
rect 65820 137658 65876 137660
rect 65900 137658 65956 137660
rect 65660 137606 65706 137658
rect 65706 137606 65716 137658
rect 65740 137606 65770 137658
rect 65770 137606 65782 137658
rect 65782 137606 65796 137658
rect 65820 137606 65834 137658
rect 65834 137606 65846 137658
rect 65846 137606 65876 137658
rect 65900 137606 65910 137658
rect 65910 137606 65956 137658
rect 65660 137604 65716 137606
rect 65740 137604 65796 137606
rect 65820 137604 65876 137606
rect 65900 137604 65956 137606
rect 96380 137658 96436 137660
rect 96460 137658 96516 137660
rect 96540 137658 96596 137660
rect 96620 137658 96676 137660
rect 96380 137606 96426 137658
rect 96426 137606 96436 137658
rect 96460 137606 96490 137658
rect 96490 137606 96502 137658
rect 96502 137606 96516 137658
rect 96540 137606 96554 137658
rect 96554 137606 96566 137658
rect 96566 137606 96596 137658
rect 96620 137606 96630 137658
rect 96630 137606 96676 137658
rect 96380 137604 96436 137606
rect 96460 137604 96516 137606
rect 96540 137604 96596 137606
rect 96620 137604 96676 137606
rect 4880 137114 4936 137116
rect 4960 137114 5016 137116
rect 5040 137114 5096 137116
rect 5120 137114 5176 137116
rect 4880 137062 4926 137114
rect 4926 137062 4936 137114
rect 4960 137062 4990 137114
rect 4990 137062 5002 137114
rect 5002 137062 5016 137114
rect 5040 137062 5054 137114
rect 5054 137062 5066 137114
rect 5066 137062 5096 137114
rect 5120 137062 5130 137114
rect 5130 137062 5176 137114
rect 4880 137060 4936 137062
rect 4960 137060 5016 137062
rect 5040 137060 5096 137062
rect 5120 137060 5176 137062
rect 35600 137114 35656 137116
rect 35680 137114 35736 137116
rect 35760 137114 35816 137116
rect 35840 137114 35896 137116
rect 35600 137062 35646 137114
rect 35646 137062 35656 137114
rect 35680 137062 35710 137114
rect 35710 137062 35722 137114
rect 35722 137062 35736 137114
rect 35760 137062 35774 137114
rect 35774 137062 35786 137114
rect 35786 137062 35816 137114
rect 35840 137062 35850 137114
rect 35850 137062 35896 137114
rect 35600 137060 35656 137062
rect 35680 137060 35736 137062
rect 35760 137060 35816 137062
rect 35840 137060 35896 137062
rect 66320 137114 66376 137116
rect 66400 137114 66456 137116
rect 66480 137114 66536 137116
rect 66560 137114 66616 137116
rect 66320 137062 66366 137114
rect 66366 137062 66376 137114
rect 66400 137062 66430 137114
rect 66430 137062 66442 137114
rect 66442 137062 66456 137114
rect 66480 137062 66494 137114
rect 66494 137062 66506 137114
rect 66506 137062 66536 137114
rect 66560 137062 66570 137114
rect 66570 137062 66616 137114
rect 66320 137060 66376 137062
rect 66400 137060 66456 137062
rect 66480 137060 66536 137062
rect 66560 137060 66616 137062
rect 97040 137114 97096 137116
rect 97120 137114 97176 137116
rect 97200 137114 97256 137116
rect 97280 137114 97336 137116
rect 97040 137062 97086 137114
rect 97086 137062 97096 137114
rect 97120 137062 97150 137114
rect 97150 137062 97162 137114
rect 97162 137062 97176 137114
rect 97200 137062 97214 137114
rect 97214 137062 97226 137114
rect 97226 137062 97256 137114
rect 97280 137062 97290 137114
rect 97290 137062 97336 137114
rect 97040 137060 97096 137062
rect 97120 137060 97176 137062
rect 97200 137060 97256 137062
rect 97280 137060 97336 137062
rect 4220 136570 4276 136572
rect 4300 136570 4356 136572
rect 4380 136570 4436 136572
rect 4460 136570 4516 136572
rect 4220 136518 4266 136570
rect 4266 136518 4276 136570
rect 4300 136518 4330 136570
rect 4330 136518 4342 136570
rect 4342 136518 4356 136570
rect 4380 136518 4394 136570
rect 4394 136518 4406 136570
rect 4406 136518 4436 136570
rect 4460 136518 4470 136570
rect 4470 136518 4516 136570
rect 4220 136516 4276 136518
rect 4300 136516 4356 136518
rect 4380 136516 4436 136518
rect 4460 136516 4516 136518
rect 34940 136570 34996 136572
rect 35020 136570 35076 136572
rect 35100 136570 35156 136572
rect 35180 136570 35236 136572
rect 34940 136518 34986 136570
rect 34986 136518 34996 136570
rect 35020 136518 35050 136570
rect 35050 136518 35062 136570
rect 35062 136518 35076 136570
rect 35100 136518 35114 136570
rect 35114 136518 35126 136570
rect 35126 136518 35156 136570
rect 35180 136518 35190 136570
rect 35190 136518 35236 136570
rect 34940 136516 34996 136518
rect 35020 136516 35076 136518
rect 35100 136516 35156 136518
rect 35180 136516 35236 136518
rect 65660 136570 65716 136572
rect 65740 136570 65796 136572
rect 65820 136570 65876 136572
rect 65900 136570 65956 136572
rect 65660 136518 65706 136570
rect 65706 136518 65716 136570
rect 65740 136518 65770 136570
rect 65770 136518 65782 136570
rect 65782 136518 65796 136570
rect 65820 136518 65834 136570
rect 65834 136518 65846 136570
rect 65846 136518 65876 136570
rect 65900 136518 65910 136570
rect 65910 136518 65956 136570
rect 65660 136516 65716 136518
rect 65740 136516 65796 136518
rect 65820 136516 65876 136518
rect 65900 136516 65956 136518
rect 96380 136570 96436 136572
rect 96460 136570 96516 136572
rect 96540 136570 96596 136572
rect 96620 136570 96676 136572
rect 96380 136518 96426 136570
rect 96426 136518 96436 136570
rect 96460 136518 96490 136570
rect 96490 136518 96502 136570
rect 96502 136518 96516 136570
rect 96540 136518 96554 136570
rect 96554 136518 96566 136570
rect 96566 136518 96596 136570
rect 96620 136518 96630 136570
rect 96630 136518 96676 136570
rect 96380 136516 96436 136518
rect 96460 136516 96516 136518
rect 96540 136516 96596 136518
rect 96620 136516 96676 136518
rect 105928 136570 105984 136572
rect 106008 136570 106064 136572
rect 106088 136570 106144 136572
rect 106168 136570 106224 136572
rect 105928 136518 105974 136570
rect 105974 136518 105984 136570
rect 106008 136518 106038 136570
rect 106038 136518 106050 136570
rect 106050 136518 106064 136570
rect 106088 136518 106102 136570
rect 106102 136518 106114 136570
rect 106114 136518 106144 136570
rect 106168 136518 106178 136570
rect 106178 136518 106224 136570
rect 105928 136516 105984 136518
rect 106008 136516 106064 136518
rect 106088 136516 106144 136518
rect 106168 136516 106224 136518
rect 4880 136026 4936 136028
rect 4960 136026 5016 136028
rect 5040 136026 5096 136028
rect 5120 136026 5176 136028
rect 4880 135974 4926 136026
rect 4926 135974 4936 136026
rect 4960 135974 4990 136026
rect 4990 135974 5002 136026
rect 5002 135974 5016 136026
rect 5040 135974 5054 136026
rect 5054 135974 5066 136026
rect 5066 135974 5096 136026
rect 5120 135974 5130 136026
rect 5130 135974 5176 136026
rect 4880 135972 4936 135974
rect 4960 135972 5016 135974
rect 5040 135972 5096 135974
rect 5120 135972 5176 135974
rect 4220 135482 4276 135484
rect 4300 135482 4356 135484
rect 4380 135482 4436 135484
rect 4460 135482 4516 135484
rect 4220 135430 4266 135482
rect 4266 135430 4276 135482
rect 4300 135430 4330 135482
rect 4330 135430 4342 135482
rect 4342 135430 4356 135482
rect 4380 135430 4394 135482
rect 4394 135430 4406 135482
rect 4406 135430 4436 135482
rect 4460 135430 4470 135482
rect 4470 135430 4516 135482
rect 4220 135428 4276 135430
rect 4300 135428 4356 135430
rect 4380 135428 4436 135430
rect 4460 135428 4516 135430
rect 4880 134938 4936 134940
rect 4960 134938 5016 134940
rect 5040 134938 5096 134940
rect 5120 134938 5176 134940
rect 4880 134886 4926 134938
rect 4926 134886 4936 134938
rect 4960 134886 4990 134938
rect 4990 134886 5002 134938
rect 5002 134886 5016 134938
rect 5040 134886 5054 134938
rect 5054 134886 5066 134938
rect 5066 134886 5096 134938
rect 5120 134886 5130 134938
rect 5130 134886 5176 134938
rect 4880 134884 4936 134886
rect 4960 134884 5016 134886
rect 5040 134884 5096 134886
rect 5120 134884 5176 134886
rect 4220 134394 4276 134396
rect 4300 134394 4356 134396
rect 4380 134394 4436 134396
rect 4460 134394 4516 134396
rect 4220 134342 4266 134394
rect 4266 134342 4276 134394
rect 4300 134342 4330 134394
rect 4330 134342 4342 134394
rect 4342 134342 4356 134394
rect 4380 134342 4394 134394
rect 4394 134342 4406 134394
rect 4406 134342 4436 134394
rect 4460 134342 4470 134394
rect 4470 134342 4516 134394
rect 4220 134340 4276 134342
rect 4300 134340 4356 134342
rect 4380 134340 4436 134342
rect 4460 134340 4516 134342
rect 4880 133850 4936 133852
rect 4960 133850 5016 133852
rect 5040 133850 5096 133852
rect 5120 133850 5176 133852
rect 4880 133798 4926 133850
rect 4926 133798 4936 133850
rect 4960 133798 4990 133850
rect 4990 133798 5002 133850
rect 5002 133798 5016 133850
rect 5040 133798 5054 133850
rect 5054 133798 5066 133850
rect 5066 133798 5096 133850
rect 5120 133798 5130 133850
rect 5130 133798 5176 133850
rect 4880 133796 4936 133798
rect 4960 133796 5016 133798
rect 5040 133796 5096 133798
rect 5120 133796 5176 133798
rect 4220 133306 4276 133308
rect 4300 133306 4356 133308
rect 4380 133306 4436 133308
rect 4460 133306 4516 133308
rect 4220 133254 4266 133306
rect 4266 133254 4276 133306
rect 4300 133254 4330 133306
rect 4330 133254 4342 133306
rect 4342 133254 4356 133306
rect 4380 133254 4394 133306
rect 4394 133254 4406 133306
rect 4406 133254 4436 133306
rect 4460 133254 4470 133306
rect 4470 133254 4516 133306
rect 4220 133252 4276 133254
rect 4300 133252 4356 133254
rect 4380 133252 4436 133254
rect 4460 133252 4516 133254
rect 4880 132762 4936 132764
rect 4960 132762 5016 132764
rect 5040 132762 5096 132764
rect 5120 132762 5176 132764
rect 4880 132710 4926 132762
rect 4926 132710 4936 132762
rect 4960 132710 4990 132762
rect 4990 132710 5002 132762
rect 5002 132710 5016 132762
rect 5040 132710 5054 132762
rect 5054 132710 5066 132762
rect 5066 132710 5096 132762
rect 5120 132710 5130 132762
rect 5130 132710 5176 132762
rect 4880 132708 4936 132710
rect 4960 132708 5016 132710
rect 5040 132708 5096 132710
rect 5120 132708 5176 132710
rect 4220 132218 4276 132220
rect 4300 132218 4356 132220
rect 4380 132218 4436 132220
rect 4460 132218 4516 132220
rect 4220 132166 4266 132218
rect 4266 132166 4276 132218
rect 4300 132166 4330 132218
rect 4330 132166 4342 132218
rect 4342 132166 4356 132218
rect 4380 132166 4394 132218
rect 4394 132166 4406 132218
rect 4406 132166 4436 132218
rect 4460 132166 4470 132218
rect 4470 132166 4516 132218
rect 4220 132164 4276 132166
rect 4300 132164 4356 132166
rect 4380 132164 4436 132166
rect 4460 132164 4516 132166
rect 4880 131674 4936 131676
rect 4960 131674 5016 131676
rect 5040 131674 5096 131676
rect 5120 131674 5176 131676
rect 4880 131622 4926 131674
rect 4926 131622 4936 131674
rect 4960 131622 4990 131674
rect 4990 131622 5002 131674
rect 5002 131622 5016 131674
rect 5040 131622 5054 131674
rect 5054 131622 5066 131674
rect 5066 131622 5096 131674
rect 5120 131622 5130 131674
rect 5130 131622 5176 131674
rect 4880 131620 4936 131622
rect 4960 131620 5016 131622
rect 5040 131620 5096 131622
rect 5120 131620 5176 131622
rect 4220 131130 4276 131132
rect 4300 131130 4356 131132
rect 4380 131130 4436 131132
rect 4460 131130 4516 131132
rect 4220 131078 4266 131130
rect 4266 131078 4276 131130
rect 4300 131078 4330 131130
rect 4330 131078 4342 131130
rect 4342 131078 4356 131130
rect 4380 131078 4394 131130
rect 4394 131078 4406 131130
rect 4406 131078 4436 131130
rect 4460 131078 4470 131130
rect 4470 131078 4516 131130
rect 4220 131076 4276 131078
rect 4300 131076 4356 131078
rect 4380 131076 4436 131078
rect 4460 131076 4516 131078
rect 4880 130586 4936 130588
rect 4960 130586 5016 130588
rect 5040 130586 5096 130588
rect 5120 130586 5176 130588
rect 4880 130534 4926 130586
rect 4926 130534 4936 130586
rect 4960 130534 4990 130586
rect 4990 130534 5002 130586
rect 5002 130534 5016 130586
rect 5040 130534 5054 130586
rect 5054 130534 5066 130586
rect 5066 130534 5096 130586
rect 5120 130534 5130 130586
rect 5130 130534 5176 130586
rect 4880 130532 4936 130534
rect 4960 130532 5016 130534
rect 5040 130532 5096 130534
rect 5120 130532 5176 130534
rect 4220 130042 4276 130044
rect 4300 130042 4356 130044
rect 4380 130042 4436 130044
rect 4460 130042 4516 130044
rect 4220 129990 4266 130042
rect 4266 129990 4276 130042
rect 4300 129990 4330 130042
rect 4330 129990 4342 130042
rect 4342 129990 4356 130042
rect 4380 129990 4394 130042
rect 4394 129990 4406 130042
rect 4406 129990 4436 130042
rect 4460 129990 4470 130042
rect 4470 129990 4516 130042
rect 4220 129988 4276 129990
rect 4300 129988 4356 129990
rect 4380 129988 4436 129990
rect 4460 129988 4516 129990
rect 4880 129498 4936 129500
rect 4960 129498 5016 129500
rect 5040 129498 5096 129500
rect 5120 129498 5176 129500
rect 4880 129446 4926 129498
rect 4926 129446 4936 129498
rect 4960 129446 4990 129498
rect 4990 129446 5002 129498
rect 5002 129446 5016 129498
rect 5040 129446 5054 129498
rect 5054 129446 5066 129498
rect 5066 129446 5096 129498
rect 5120 129446 5130 129498
rect 5130 129446 5176 129498
rect 4880 129444 4936 129446
rect 4960 129444 5016 129446
rect 5040 129444 5096 129446
rect 5120 129444 5176 129446
rect 4220 128954 4276 128956
rect 4300 128954 4356 128956
rect 4380 128954 4436 128956
rect 4460 128954 4516 128956
rect 4220 128902 4266 128954
rect 4266 128902 4276 128954
rect 4300 128902 4330 128954
rect 4330 128902 4342 128954
rect 4342 128902 4356 128954
rect 4380 128902 4394 128954
rect 4394 128902 4406 128954
rect 4406 128902 4436 128954
rect 4460 128902 4470 128954
rect 4470 128902 4516 128954
rect 4220 128900 4276 128902
rect 4300 128900 4356 128902
rect 4380 128900 4436 128902
rect 4460 128900 4516 128902
rect 4880 128410 4936 128412
rect 4960 128410 5016 128412
rect 5040 128410 5096 128412
rect 5120 128410 5176 128412
rect 4880 128358 4926 128410
rect 4926 128358 4936 128410
rect 4960 128358 4990 128410
rect 4990 128358 5002 128410
rect 5002 128358 5016 128410
rect 5040 128358 5054 128410
rect 5054 128358 5066 128410
rect 5066 128358 5096 128410
rect 5120 128358 5130 128410
rect 5130 128358 5176 128410
rect 4880 128356 4936 128358
rect 4960 128356 5016 128358
rect 5040 128356 5096 128358
rect 5120 128356 5176 128358
rect 4220 127866 4276 127868
rect 4300 127866 4356 127868
rect 4380 127866 4436 127868
rect 4460 127866 4516 127868
rect 4220 127814 4266 127866
rect 4266 127814 4276 127866
rect 4300 127814 4330 127866
rect 4330 127814 4342 127866
rect 4342 127814 4356 127866
rect 4380 127814 4394 127866
rect 4394 127814 4406 127866
rect 4406 127814 4436 127866
rect 4460 127814 4470 127866
rect 4470 127814 4516 127866
rect 4220 127812 4276 127814
rect 4300 127812 4356 127814
rect 4380 127812 4436 127814
rect 4460 127812 4516 127814
rect 4880 127322 4936 127324
rect 4960 127322 5016 127324
rect 5040 127322 5096 127324
rect 5120 127322 5176 127324
rect 4880 127270 4926 127322
rect 4926 127270 4936 127322
rect 4960 127270 4990 127322
rect 4990 127270 5002 127322
rect 5002 127270 5016 127322
rect 5040 127270 5054 127322
rect 5054 127270 5066 127322
rect 5066 127270 5096 127322
rect 5120 127270 5130 127322
rect 5130 127270 5176 127322
rect 4880 127268 4936 127270
rect 4960 127268 5016 127270
rect 5040 127268 5096 127270
rect 5120 127268 5176 127270
rect 4220 126778 4276 126780
rect 4300 126778 4356 126780
rect 4380 126778 4436 126780
rect 4460 126778 4516 126780
rect 4220 126726 4266 126778
rect 4266 126726 4276 126778
rect 4300 126726 4330 126778
rect 4330 126726 4342 126778
rect 4342 126726 4356 126778
rect 4380 126726 4394 126778
rect 4394 126726 4406 126778
rect 4406 126726 4436 126778
rect 4460 126726 4470 126778
rect 4470 126726 4516 126778
rect 4220 126724 4276 126726
rect 4300 126724 4356 126726
rect 4380 126724 4436 126726
rect 4460 126724 4516 126726
rect 4880 126234 4936 126236
rect 4960 126234 5016 126236
rect 5040 126234 5096 126236
rect 5120 126234 5176 126236
rect 4880 126182 4926 126234
rect 4926 126182 4936 126234
rect 4960 126182 4990 126234
rect 4990 126182 5002 126234
rect 5002 126182 5016 126234
rect 5040 126182 5054 126234
rect 5054 126182 5066 126234
rect 5066 126182 5096 126234
rect 5120 126182 5130 126234
rect 5130 126182 5176 126234
rect 4880 126180 4936 126182
rect 4960 126180 5016 126182
rect 5040 126180 5096 126182
rect 5120 126180 5176 126182
rect 4220 125690 4276 125692
rect 4300 125690 4356 125692
rect 4380 125690 4436 125692
rect 4460 125690 4516 125692
rect 4220 125638 4266 125690
rect 4266 125638 4276 125690
rect 4300 125638 4330 125690
rect 4330 125638 4342 125690
rect 4342 125638 4356 125690
rect 4380 125638 4394 125690
rect 4394 125638 4406 125690
rect 4406 125638 4436 125690
rect 4460 125638 4470 125690
rect 4470 125638 4516 125690
rect 4220 125636 4276 125638
rect 4300 125636 4356 125638
rect 4380 125636 4436 125638
rect 4460 125636 4516 125638
rect 4880 125146 4936 125148
rect 4960 125146 5016 125148
rect 5040 125146 5096 125148
rect 5120 125146 5176 125148
rect 4880 125094 4926 125146
rect 4926 125094 4936 125146
rect 4960 125094 4990 125146
rect 4990 125094 5002 125146
rect 5002 125094 5016 125146
rect 5040 125094 5054 125146
rect 5054 125094 5066 125146
rect 5066 125094 5096 125146
rect 5120 125094 5130 125146
rect 5130 125094 5176 125146
rect 4880 125092 4936 125094
rect 4960 125092 5016 125094
rect 5040 125092 5096 125094
rect 5120 125092 5176 125094
rect 4220 124602 4276 124604
rect 4300 124602 4356 124604
rect 4380 124602 4436 124604
rect 4460 124602 4516 124604
rect 4220 124550 4266 124602
rect 4266 124550 4276 124602
rect 4300 124550 4330 124602
rect 4330 124550 4342 124602
rect 4342 124550 4356 124602
rect 4380 124550 4394 124602
rect 4394 124550 4406 124602
rect 4406 124550 4436 124602
rect 4460 124550 4470 124602
rect 4470 124550 4516 124602
rect 4220 124548 4276 124550
rect 4300 124548 4356 124550
rect 4380 124548 4436 124550
rect 4460 124548 4516 124550
rect 4880 124058 4936 124060
rect 4960 124058 5016 124060
rect 5040 124058 5096 124060
rect 5120 124058 5176 124060
rect 4880 124006 4926 124058
rect 4926 124006 4936 124058
rect 4960 124006 4990 124058
rect 4990 124006 5002 124058
rect 5002 124006 5016 124058
rect 5040 124006 5054 124058
rect 5054 124006 5066 124058
rect 5066 124006 5096 124058
rect 5120 124006 5130 124058
rect 5130 124006 5176 124058
rect 4880 124004 4936 124006
rect 4960 124004 5016 124006
rect 5040 124004 5096 124006
rect 5120 124004 5176 124006
rect 4220 123514 4276 123516
rect 4300 123514 4356 123516
rect 4380 123514 4436 123516
rect 4460 123514 4516 123516
rect 4220 123462 4266 123514
rect 4266 123462 4276 123514
rect 4300 123462 4330 123514
rect 4330 123462 4342 123514
rect 4342 123462 4356 123514
rect 4380 123462 4394 123514
rect 4394 123462 4406 123514
rect 4406 123462 4436 123514
rect 4460 123462 4470 123514
rect 4470 123462 4516 123514
rect 4220 123460 4276 123462
rect 4300 123460 4356 123462
rect 4380 123460 4436 123462
rect 4460 123460 4516 123462
rect 4880 122970 4936 122972
rect 4960 122970 5016 122972
rect 5040 122970 5096 122972
rect 5120 122970 5176 122972
rect 4880 122918 4926 122970
rect 4926 122918 4936 122970
rect 4960 122918 4990 122970
rect 4990 122918 5002 122970
rect 5002 122918 5016 122970
rect 5040 122918 5054 122970
rect 5054 122918 5066 122970
rect 5066 122918 5096 122970
rect 5120 122918 5130 122970
rect 5130 122918 5176 122970
rect 4880 122916 4936 122918
rect 4960 122916 5016 122918
rect 5040 122916 5096 122918
rect 5120 122916 5176 122918
rect 4220 122426 4276 122428
rect 4300 122426 4356 122428
rect 4380 122426 4436 122428
rect 4460 122426 4516 122428
rect 4220 122374 4266 122426
rect 4266 122374 4276 122426
rect 4300 122374 4330 122426
rect 4330 122374 4342 122426
rect 4342 122374 4356 122426
rect 4380 122374 4394 122426
rect 4394 122374 4406 122426
rect 4406 122374 4436 122426
rect 4460 122374 4470 122426
rect 4470 122374 4516 122426
rect 4220 122372 4276 122374
rect 4300 122372 4356 122374
rect 4380 122372 4436 122374
rect 4460 122372 4516 122374
rect 4880 121882 4936 121884
rect 4960 121882 5016 121884
rect 5040 121882 5096 121884
rect 5120 121882 5176 121884
rect 4880 121830 4926 121882
rect 4926 121830 4936 121882
rect 4960 121830 4990 121882
rect 4990 121830 5002 121882
rect 5002 121830 5016 121882
rect 5040 121830 5054 121882
rect 5054 121830 5066 121882
rect 5066 121830 5096 121882
rect 5120 121830 5130 121882
rect 5130 121830 5176 121882
rect 4880 121828 4936 121830
rect 4960 121828 5016 121830
rect 5040 121828 5096 121830
rect 5120 121828 5176 121830
rect 4220 121338 4276 121340
rect 4300 121338 4356 121340
rect 4380 121338 4436 121340
rect 4460 121338 4516 121340
rect 4220 121286 4266 121338
rect 4266 121286 4276 121338
rect 4300 121286 4330 121338
rect 4330 121286 4342 121338
rect 4342 121286 4356 121338
rect 4380 121286 4394 121338
rect 4394 121286 4406 121338
rect 4406 121286 4436 121338
rect 4460 121286 4470 121338
rect 4470 121286 4516 121338
rect 4220 121284 4276 121286
rect 4300 121284 4356 121286
rect 4380 121284 4436 121286
rect 4460 121284 4516 121286
rect 4880 120794 4936 120796
rect 4960 120794 5016 120796
rect 5040 120794 5096 120796
rect 5120 120794 5176 120796
rect 4880 120742 4926 120794
rect 4926 120742 4936 120794
rect 4960 120742 4990 120794
rect 4990 120742 5002 120794
rect 5002 120742 5016 120794
rect 5040 120742 5054 120794
rect 5054 120742 5066 120794
rect 5066 120742 5096 120794
rect 5120 120742 5130 120794
rect 5130 120742 5176 120794
rect 4880 120740 4936 120742
rect 4960 120740 5016 120742
rect 5040 120740 5096 120742
rect 5120 120740 5176 120742
rect 4220 120250 4276 120252
rect 4300 120250 4356 120252
rect 4380 120250 4436 120252
rect 4460 120250 4516 120252
rect 4220 120198 4266 120250
rect 4266 120198 4276 120250
rect 4300 120198 4330 120250
rect 4330 120198 4342 120250
rect 4342 120198 4356 120250
rect 4380 120198 4394 120250
rect 4394 120198 4406 120250
rect 4406 120198 4436 120250
rect 4460 120198 4470 120250
rect 4470 120198 4516 120250
rect 4220 120196 4276 120198
rect 4300 120196 4356 120198
rect 4380 120196 4436 120198
rect 4460 120196 4516 120198
rect 4880 119706 4936 119708
rect 4960 119706 5016 119708
rect 5040 119706 5096 119708
rect 5120 119706 5176 119708
rect 4880 119654 4926 119706
rect 4926 119654 4936 119706
rect 4960 119654 4990 119706
rect 4990 119654 5002 119706
rect 5002 119654 5016 119706
rect 5040 119654 5054 119706
rect 5054 119654 5066 119706
rect 5066 119654 5096 119706
rect 5120 119654 5130 119706
rect 5130 119654 5176 119706
rect 4880 119652 4936 119654
rect 4960 119652 5016 119654
rect 5040 119652 5096 119654
rect 5120 119652 5176 119654
rect 4220 119162 4276 119164
rect 4300 119162 4356 119164
rect 4380 119162 4436 119164
rect 4460 119162 4516 119164
rect 4220 119110 4266 119162
rect 4266 119110 4276 119162
rect 4300 119110 4330 119162
rect 4330 119110 4342 119162
rect 4342 119110 4356 119162
rect 4380 119110 4394 119162
rect 4394 119110 4406 119162
rect 4406 119110 4436 119162
rect 4460 119110 4470 119162
rect 4470 119110 4516 119162
rect 4220 119108 4276 119110
rect 4300 119108 4356 119110
rect 4380 119108 4436 119110
rect 4460 119108 4516 119110
rect 4880 118618 4936 118620
rect 4960 118618 5016 118620
rect 5040 118618 5096 118620
rect 5120 118618 5176 118620
rect 4880 118566 4926 118618
rect 4926 118566 4936 118618
rect 4960 118566 4990 118618
rect 4990 118566 5002 118618
rect 5002 118566 5016 118618
rect 5040 118566 5054 118618
rect 5054 118566 5066 118618
rect 5066 118566 5096 118618
rect 5120 118566 5130 118618
rect 5130 118566 5176 118618
rect 4880 118564 4936 118566
rect 4960 118564 5016 118566
rect 5040 118564 5096 118566
rect 5120 118564 5176 118566
rect 4220 118074 4276 118076
rect 4300 118074 4356 118076
rect 4380 118074 4436 118076
rect 4460 118074 4516 118076
rect 4220 118022 4266 118074
rect 4266 118022 4276 118074
rect 4300 118022 4330 118074
rect 4330 118022 4342 118074
rect 4342 118022 4356 118074
rect 4380 118022 4394 118074
rect 4394 118022 4406 118074
rect 4406 118022 4436 118074
rect 4460 118022 4470 118074
rect 4470 118022 4516 118074
rect 4220 118020 4276 118022
rect 4300 118020 4356 118022
rect 4380 118020 4436 118022
rect 4460 118020 4516 118022
rect 4880 117530 4936 117532
rect 4960 117530 5016 117532
rect 5040 117530 5096 117532
rect 5120 117530 5176 117532
rect 4880 117478 4926 117530
rect 4926 117478 4936 117530
rect 4960 117478 4990 117530
rect 4990 117478 5002 117530
rect 5002 117478 5016 117530
rect 5040 117478 5054 117530
rect 5054 117478 5066 117530
rect 5066 117478 5096 117530
rect 5120 117478 5130 117530
rect 5130 117478 5176 117530
rect 4880 117476 4936 117478
rect 4960 117476 5016 117478
rect 5040 117476 5096 117478
rect 5120 117476 5176 117478
rect 4220 116986 4276 116988
rect 4300 116986 4356 116988
rect 4380 116986 4436 116988
rect 4460 116986 4516 116988
rect 4220 116934 4266 116986
rect 4266 116934 4276 116986
rect 4300 116934 4330 116986
rect 4330 116934 4342 116986
rect 4342 116934 4356 116986
rect 4380 116934 4394 116986
rect 4394 116934 4406 116986
rect 4406 116934 4436 116986
rect 4460 116934 4470 116986
rect 4470 116934 4516 116986
rect 4220 116932 4276 116934
rect 4300 116932 4356 116934
rect 4380 116932 4436 116934
rect 4460 116932 4516 116934
rect 4880 116442 4936 116444
rect 4960 116442 5016 116444
rect 5040 116442 5096 116444
rect 5120 116442 5176 116444
rect 4880 116390 4926 116442
rect 4926 116390 4936 116442
rect 4960 116390 4990 116442
rect 4990 116390 5002 116442
rect 5002 116390 5016 116442
rect 5040 116390 5054 116442
rect 5054 116390 5066 116442
rect 5066 116390 5096 116442
rect 5120 116390 5130 116442
rect 5130 116390 5176 116442
rect 4880 116388 4936 116390
rect 4960 116388 5016 116390
rect 5040 116388 5096 116390
rect 5120 116388 5176 116390
rect 4220 115898 4276 115900
rect 4300 115898 4356 115900
rect 4380 115898 4436 115900
rect 4460 115898 4516 115900
rect 4220 115846 4266 115898
rect 4266 115846 4276 115898
rect 4300 115846 4330 115898
rect 4330 115846 4342 115898
rect 4342 115846 4356 115898
rect 4380 115846 4394 115898
rect 4394 115846 4406 115898
rect 4406 115846 4436 115898
rect 4460 115846 4470 115898
rect 4470 115846 4516 115898
rect 4220 115844 4276 115846
rect 4300 115844 4356 115846
rect 4380 115844 4436 115846
rect 4460 115844 4516 115846
rect 4880 115354 4936 115356
rect 4960 115354 5016 115356
rect 5040 115354 5096 115356
rect 5120 115354 5176 115356
rect 4880 115302 4926 115354
rect 4926 115302 4936 115354
rect 4960 115302 4990 115354
rect 4990 115302 5002 115354
rect 5002 115302 5016 115354
rect 5040 115302 5054 115354
rect 5054 115302 5066 115354
rect 5066 115302 5096 115354
rect 5120 115302 5130 115354
rect 5130 115302 5176 115354
rect 4880 115300 4936 115302
rect 4960 115300 5016 115302
rect 5040 115300 5096 115302
rect 5120 115300 5176 115302
rect 4220 114810 4276 114812
rect 4300 114810 4356 114812
rect 4380 114810 4436 114812
rect 4460 114810 4516 114812
rect 4220 114758 4266 114810
rect 4266 114758 4276 114810
rect 4300 114758 4330 114810
rect 4330 114758 4342 114810
rect 4342 114758 4356 114810
rect 4380 114758 4394 114810
rect 4394 114758 4406 114810
rect 4406 114758 4436 114810
rect 4460 114758 4470 114810
rect 4470 114758 4516 114810
rect 4220 114756 4276 114758
rect 4300 114756 4356 114758
rect 4380 114756 4436 114758
rect 4460 114756 4516 114758
rect 4880 114266 4936 114268
rect 4960 114266 5016 114268
rect 5040 114266 5096 114268
rect 5120 114266 5176 114268
rect 4880 114214 4926 114266
rect 4926 114214 4936 114266
rect 4960 114214 4990 114266
rect 4990 114214 5002 114266
rect 5002 114214 5016 114266
rect 5040 114214 5054 114266
rect 5054 114214 5066 114266
rect 5066 114214 5096 114266
rect 5120 114214 5130 114266
rect 5130 114214 5176 114266
rect 4880 114212 4936 114214
rect 4960 114212 5016 114214
rect 5040 114212 5096 114214
rect 5120 114212 5176 114214
rect 4220 113722 4276 113724
rect 4300 113722 4356 113724
rect 4380 113722 4436 113724
rect 4460 113722 4516 113724
rect 4220 113670 4266 113722
rect 4266 113670 4276 113722
rect 4300 113670 4330 113722
rect 4330 113670 4342 113722
rect 4342 113670 4356 113722
rect 4380 113670 4394 113722
rect 4394 113670 4406 113722
rect 4406 113670 4436 113722
rect 4460 113670 4470 113722
rect 4470 113670 4516 113722
rect 4220 113668 4276 113670
rect 4300 113668 4356 113670
rect 4380 113668 4436 113670
rect 4460 113668 4516 113670
rect 4880 113178 4936 113180
rect 4960 113178 5016 113180
rect 5040 113178 5096 113180
rect 5120 113178 5176 113180
rect 4880 113126 4926 113178
rect 4926 113126 4936 113178
rect 4960 113126 4990 113178
rect 4990 113126 5002 113178
rect 5002 113126 5016 113178
rect 5040 113126 5054 113178
rect 5054 113126 5066 113178
rect 5066 113126 5096 113178
rect 5120 113126 5130 113178
rect 5130 113126 5176 113178
rect 4880 113124 4936 113126
rect 4960 113124 5016 113126
rect 5040 113124 5096 113126
rect 5120 113124 5176 113126
rect 4220 112634 4276 112636
rect 4300 112634 4356 112636
rect 4380 112634 4436 112636
rect 4460 112634 4516 112636
rect 4220 112582 4266 112634
rect 4266 112582 4276 112634
rect 4300 112582 4330 112634
rect 4330 112582 4342 112634
rect 4342 112582 4356 112634
rect 4380 112582 4394 112634
rect 4394 112582 4406 112634
rect 4406 112582 4436 112634
rect 4460 112582 4470 112634
rect 4470 112582 4516 112634
rect 4220 112580 4276 112582
rect 4300 112580 4356 112582
rect 4380 112580 4436 112582
rect 4460 112580 4516 112582
rect 4880 112090 4936 112092
rect 4960 112090 5016 112092
rect 5040 112090 5096 112092
rect 5120 112090 5176 112092
rect 4880 112038 4926 112090
rect 4926 112038 4936 112090
rect 4960 112038 4990 112090
rect 4990 112038 5002 112090
rect 5002 112038 5016 112090
rect 5040 112038 5054 112090
rect 5054 112038 5066 112090
rect 5066 112038 5096 112090
rect 5120 112038 5130 112090
rect 5130 112038 5176 112090
rect 4880 112036 4936 112038
rect 4960 112036 5016 112038
rect 5040 112036 5096 112038
rect 5120 112036 5176 112038
rect 4220 111546 4276 111548
rect 4300 111546 4356 111548
rect 4380 111546 4436 111548
rect 4460 111546 4516 111548
rect 4220 111494 4266 111546
rect 4266 111494 4276 111546
rect 4300 111494 4330 111546
rect 4330 111494 4342 111546
rect 4342 111494 4356 111546
rect 4380 111494 4394 111546
rect 4394 111494 4406 111546
rect 4406 111494 4436 111546
rect 4460 111494 4470 111546
rect 4470 111494 4516 111546
rect 4220 111492 4276 111494
rect 4300 111492 4356 111494
rect 4380 111492 4436 111494
rect 4460 111492 4516 111494
rect 4880 111002 4936 111004
rect 4960 111002 5016 111004
rect 5040 111002 5096 111004
rect 5120 111002 5176 111004
rect 4880 110950 4926 111002
rect 4926 110950 4936 111002
rect 4960 110950 4990 111002
rect 4990 110950 5002 111002
rect 5002 110950 5016 111002
rect 5040 110950 5054 111002
rect 5054 110950 5066 111002
rect 5066 110950 5096 111002
rect 5120 110950 5130 111002
rect 5130 110950 5176 111002
rect 4880 110948 4936 110950
rect 4960 110948 5016 110950
rect 5040 110948 5096 110950
rect 5120 110948 5176 110950
rect 1306 110880 1362 110936
rect 4220 110458 4276 110460
rect 4300 110458 4356 110460
rect 4380 110458 4436 110460
rect 4460 110458 4516 110460
rect 4220 110406 4266 110458
rect 4266 110406 4276 110458
rect 4300 110406 4330 110458
rect 4330 110406 4342 110458
rect 4342 110406 4356 110458
rect 4380 110406 4394 110458
rect 4394 110406 4406 110458
rect 4406 110406 4436 110458
rect 4460 110406 4470 110458
rect 4470 110406 4516 110458
rect 4220 110404 4276 110406
rect 4300 110404 4356 110406
rect 4380 110404 4436 110406
rect 4460 110404 4516 110406
rect 4880 109914 4936 109916
rect 4960 109914 5016 109916
rect 5040 109914 5096 109916
rect 5120 109914 5176 109916
rect 4880 109862 4926 109914
rect 4926 109862 4936 109914
rect 4960 109862 4990 109914
rect 4990 109862 5002 109914
rect 5002 109862 5016 109914
rect 5040 109862 5054 109914
rect 5054 109862 5066 109914
rect 5066 109862 5096 109914
rect 5120 109862 5130 109914
rect 5130 109862 5176 109914
rect 4880 109860 4936 109862
rect 4960 109860 5016 109862
rect 5040 109860 5096 109862
rect 5120 109860 5176 109862
rect 1306 109520 1362 109576
rect 4220 109370 4276 109372
rect 4300 109370 4356 109372
rect 4380 109370 4436 109372
rect 4460 109370 4516 109372
rect 4220 109318 4266 109370
rect 4266 109318 4276 109370
rect 4300 109318 4330 109370
rect 4330 109318 4342 109370
rect 4342 109318 4356 109370
rect 4380 109318 4394 109370
rect 4394 109318 4406 109370
rect 4406 109318 4436 109370
rect 4460 109318 4470 109370
rect 4470 109318 4516 109370
rect 4220 109316 4276 109318
rect 4300 109316 4356 109318
rect 4380 109316 4436 109318
rect 4460 109316 4516 109318
rect 4880 108826 4936 108828
rect 4960 108826 5016 108828
rect 5040 108826 5096 108828
rect 5120 108826 5176 108828
rect 4880 108774 4926 108826
rect 4926 108774 4936 108826
rect 4960 108774 4990 108826
rect 4990 108774 5002 108826
rect 5002 108774 5016 108826
rect 5040 108774 5054 108826
rect 5054 108774 5066 108826
rect 5066 108774 5096 108826
rect 5120 108774 5130 108826
rect 5130 108774 5176 108826
rect 4880 108772 4936 108774
rect 4960 108772 5016 108774
rect 5040 108772 5096 108774
rect 5120 108772 5176 108774
rect 4220 108282 4276 108284
rect 4300 108282 4356 108284
rect 4380 108282 4436 108284
rect 4460 108282 4516 108284
rect 4220 108230 4266 108282
rect 4266 108230 4276 108282
rect 4300 108230 4330 108282
rect 4330 108230 4342 108282
rect 4342 108230 4356 108282
rect 4380 108230 4394 108282
rect 4394 108230 4406 108282
rect 4406 108230 4436 108282
rect 4460 108230 4470 108282
rect 4470 108230 4516 108282
rect 4220 108228 4276 108230
rect 4300 108228 4356 108230
rect 4380 108228 4436 108230
rect 4460 108228 4516 108230
rect 1306 108160 1362 108216
rect 4880 107738 4936 107740
rect 4960 107738 5016 107740
rect 5040 107738 5096 107740
rect 5120 107738 5176 107740
rect 4880 107686 4926 107738
rect 4926 107686 4936 107738
rect 4960 107686 4990 107738
rect 4990 107686 5002 107738
rect 5002 107686 5016 107738
rect 5040 107686 5054 107738
rect 5054 107686 5066 107738
rect 5066 107686 5096 107738
rect 5120 107686 5130 107738
rect 5130 107686 5176 107738
rect 4880 107684 4936 107686
rect 4960 107684 5016 107686
rect 5040 107684 5096 107686
rect 5120 107684 5176 107686
rect 4220 107194 4276 107196
rect 4300 107194 4356 107196
rect 4380 107194 4436 107196
rect 4460 107194 4516 107196
rect 4220 107142 4266 107194
rect 4266 107142 4276 107194
rect 4300 107142 4330 107194
rect 4330 107142 4342 107194
rect 4342 107142 4356 107194
rect 4380 107142 4394 107194
rect 4394 107142 4406 107194
rect 4406 107142 4436 107194
rect 4460 107142 4470 107194
rect 4470 107142 4516 107194
rect 4220 107140 4276 107142
rect 4300 107140 4356 107142
rect 4380 107140 4436 107142
rect 4460 107140 4516 107142
rect 1214 106836 1216 106856
rect 1216 106836 1268 106856
rect 1268 106836 1270 106856
rect 1214 106800 1270 106836
rect 4880 106650 4936 106652
rect 4960 106650 5016 106652
rect 5040 106650 5096 106652
rect 5120 106650 5176 106652
rect 4880 106598 4926 106650
rect 4926 106598 4936 106650
rect 4960 106598 4990 106650
rect 4990 106598 5002 106650
rect 5002 106598 5016 106650
rect 5040 106598 5054 106650
rect 5054 106598 5066 106650
rect 5066 106598 5096 106650
rect 5120 106598 5130 106650
rect 5130 106598 5176 106650
rect 4880 106596 4936 106598
rect 4960 106596 5016 106598
rect 5040 106596 5096 106598
rect 5120 106596 5176 106598
rect 4220 106106 4276 106108
rect 4300 106106 4356 106108
rect 4380 106106 4436 106108
rect 4460 106106 4516 106108
rect 4220 106054 4266 106106
rect 4266 106054 4276 106106
rect 4300 106054 4330 106106
rect 4330 106054 4342 106106
rect 4342 106054 4356 106106
rect 4380 106054 4394 106106
rect 4394 106054 4406 106106
rect 4406 106054 4436 106106
rect 4460 106054 4470 106106
rect 4470 106054 4516 106106
rect 4220 106052 4276 106054
rect 4300 106052 4356 106054
rect 4380 106052 4436 106054
rect 4460 106052 4516 106054
rect 4880 105562 4936 105564
rect 4960 105562 5016 105564
rect 5040 105562 5096 105564
rect 5120 105562 5176 105564
rect 4880 105510 4926 105562
rect 4926 105510 4936 105562
rect 4960 105510 4990 105562
rect 4990 105510 5002 105562
rect 5002 105510 5016 105562
rect 5040 105510 5054 105562
rect 5054 105510 5066 105562
rect 5066 105510 5096 105562
rect 5120 105510 5130 105562
rect 5130 105510 5176 105562
rect 4880 105508 4936 105510
rect 4960 105508 5016 105510
rect 5040 105508 5096 105510
rect 5120 105508 5176 105510
rect 1306 105440 1362 105496
rect 4220 105018 4276 105020
rect 4300 105018 4356 105020
rect 4380 105018 4436 105020
rect 4460 105018 4516 105020
rect 4220 104966 4266 105018
rect 4266 104966 4276 105018
rect 4300 104966 4330 105018
rect 4330 104966 4342 105018
rect 4342 104966 4356 105018
rect 4380 104966 4394 105018
rect 4394 104966 4406 105018
rect 4406 104966 4436 105018
rect 4460 104966 4470 105018
rect 4470 104966 4516 105018
rect 4220 104964 4276 104966
rect 4300 104964 4356 104966
rect 4380 104964 4436 104966
rect 4460 104964 4516 104966
rect 4880 104474 4936 104476
rect 4960 104474 5016 104476
rect 5040 104474 5096 104476
rect 5120 104474 5176 104476
rect 4880 104422 4926 104474
rect 4926 104422 4936 104474
rect 4960 104422 4990 104474
rect 4990 104422 5002 104474
rect 5002 104422 5016 104474
rect 5040 104422 5054 104474
rect 5054 104422 5066 104474
rect 5066 104422 5096 104474
rect 5120 104422 5130 104474
rect 5130 104422 5176 104474
rect 4880 104420 4936 104422
rect 4960 104420 5016 104422
rect 5040 104420 5096 104422
rect 5120 104420 5176 104422
rect 1306 104080 1362 104136
rect 4220 103930 4276 103932
rect 4300 103930 4356 103932
rect 4380 103930 4436 103932
rect 4460 103930 4516 103932
rect 4220 103878 4266 103930
rect 4266 103878 4276 103930
rect 4300 103878 4330 103930
rect 4330 103878 4342 103930
rect 4342 103878 4356 103930
rect 4380 103878 4394 103930
rect 4394 103878 4406 103930
rect 4406 103878 4436 103930
rect 4460 103878 4470 103930
rect 4470 103878 4516 103930
rect 4220 103876 4276 103878
rect 4300 103876 4356 103878
rect 4380 103876 4436 103878
rect 4460 103876 4516 103878
rect 4880 103386 4936 103388
rect 4960 103386 5016 103388
rect 5040 103386 5096 103388
rect 5120 103386 5176 103388
rect 4880 103334 4926 103386
rect 4926 103334 4936 103386
rect 4960 103334 4990 103386
rect 4990 103334 5002 103386
rect 5002 103334 5016 103386
rect 5040 103334 5054 103386
rect 5054 103334 5066 103386
rect 5066 103334 5096 103386
rect 5120 103334 5130 103386
rect 5130 103334 5176 103386
rect 4880 103332 4936 103334
rect 4960 103332 5016 103334
rect 5040 103332 5096 103334
rect 5120 103332 5176 103334
rect 4220 102842 4276 102844
rect 4300 102842 4356 102844
rect 4380 102842 4436 102844
rect 4460 102842 4516 102844
rect 4220 102790 4266 102842
rect 4266 102790 4276 102842
rect 4300 102790 4330 102842
rect 4330 102790 4342 102842
rect 4342 102790 4356 102842
rect 4380 102790 4394 102842
rect 4394 102790 4406 102842
rect 4406 102790 4436 102842
rect 4460 102790 4470 102842
rect 4470 102790 4516 102842
rect 4220 102788 4276 102790
rect 4300 102788 4356 102790
rect 4380 102788 4436 102790
rect 4460 102788 4516 102790
rect 4880 102298 4936 102300
rect 4960 102298 5016 102300
rect 5040 102298 5096 102300
rect 5120 102298 5176 102300
rect 4880 102246 4926 102298
rect 4926 102246 4936 102298
rect 4960 102246 4990 102298
rect 4990 102246 5002 102298
rect 5002 102246 5016 102298
rect 5040 102246 5054 102298
rect 5054 102246 5066 102298
rect 5066 102246 5096 102298
rect 5120 102246 5130 102298
rect 5130 102246 5176 102298
rect 4880 102244 4936 102246
rect 4960 102244 5016 102246
rect 5040 102244 5096 102246
rect 5120 102244 5176 102246
rect 4220 101754 4276 101756
rect 4300 101754 4356 101756
rect 4380 101754 4436 101756
rect 4460 101754 4516 101756
rect 4220 101702 4266 101754
rect 4266 101702 4276 101754
rect 4300 101702 4330 101754
rect 4330 101702 4342 101754
rect 4342 101702 4356 101754
rect 4380 101702 4394 101754
rect 4394 101702 4406 101754
rect 4406 101702 4436 101754
rect 4460 101702 4470 101754
rect 4470 101702 4516 101754
rect 4220 101700 4276 101702
rect 4300 101700 4356 101702
rect 4380 101700 4436 101702
rect 4460 101700 4516 101702
rect 4880 101210 4936 101212
rect 4960 101210 5016 101212
rect 5040 101210 5096 101212
rect 5120 101210 5176 101212
rect 4880 101158 4926 101210
rect 4926 101158 4936 101210
rect 4960 101158 4990 101210
rect 4990 101158 5002 101210
rect 5002 101158 5016 101210
rect 5040 101158 5054 101210
rect 5054 101158 5066 101210
rect 5066 101158 5096 101210
rect 5120 101158 5130 101210
rect 5130 101158 5176 101210
rect 4880 101156 4936 101158
rect 4960 101156 5016 101158
rect 5040 101156 5096 101158
rect 5120 101156 5176 101158
rect 4220 100666 4276 100668
rect 4300 100666 4356 100668
rect 4380 100666 4436 100668
rect 4460 100666 4516 100668
rect 4220 100614 4266 100666
rect 4266 100614 4276 100666
rect 4300 100614 4330 100666
rect 4330 100614 4342 100666
rect 4342 100614 4356 100666
rect 4380 100614 4394 100666
rect 4394 100614 4406 100666
rect 4406 100614 4436 100666
rect 4460 100614 4470 100666
rect 4470 100614 4516 100666
rect 4220 100612 4276 100614
rect 4300 100612 4356 100614
rect 4380 100612 4436 100614
rect 4460 100612 4516 100614
rect 4880 100122 4936 100124
rect 4960 100122 5016 100124
rect 5040 100122 5096 100124
rect 5120 100122 5176 100124
rect 4880 100070 4926 100122
rect 4926 100070 4936 100122
rect 4960 100070 4990 100122
rect 4990 100070 5002 100122
rect 5002 100070 5016 100122
rect 5040 100070 5054 100122
rect 5054 100070 5066 100122
rect 5066 100070 5096 100122
rect 5120 100070 5130 100122
rect 5130 100070 5176 100122
rect 4880 100068 4936 100070
rect 4960 100068 5016 100070
rect 5040 100068 5096 100070
rect 5120 100068 5176 100070
rect 4220 99578 4276 99580
rect 4300 99578 4356 99580
rect 4380 99578 4436 99580
rect 4460 99578 4516 99580
rect 4220 99526 4266 99578
rect 4266 99526 4276 99578
rect 4300 99526 4330 99578
rect 4330 99526 4342 99578
rect 4342 99526 4356 99578
rect 4380 99526 4394 99578
rect 4394 99526 4406 99578
rect 4406 99526 4436 99578
rect 4460 99526 4470 99578
rect 4470 99526 4516 99578
rect 4220 99524 4276 99526
rect 4300 99524 4356 99526
rect 4380 99524 4436 99526
rect 4460 99524 4516 99526
rect 4880 99034 4936 99036
rect 4960 99034 5016 99036
rect 5040 99034 5096 99036
rect 5120 99034 5176 99036
rect 4880 98982 4926 99034
rect 4926 98982 4936 99034
rect 4960 98982 4990 99034
rect 4990 98982 5002 99034
rect 5002 98982 5016 99034
rect 5040 98982 5054 99034
rect 5054 98982 5066 99034
rect 5066 98982 5096 99034
rect 5120 98982 5130 99034
rect 5130 98982 5176 99034
rect 4880 98980 4936 98982
rect 4960 98980 5016 98982
rect 5040 98980 5096 98982
rect 5120 98980 5176 98982
rect 4220 98490 4276 98492
rect 4300 98490 4356 98492
rect 4380 98490 4436 98492
rect 4460 98490 4516 98492
rect 4220 98438 4266 98490
rect 4266 98438 4276 98490
rect 4300 98438 4330 98490
rect 4330 98438 4342 98490
rect 4342 98438 4356 98490
rect 4380 98438 4394 98490
rect 4394 98438 4406 98490
rect 4406 98438 4436 98490
rect 4460 98438 4470 98490
rect 4470 98438 4516 98490
rect 4220 98436 4276 98438
rect 4300 98436 4356 98438
rect 4380 98436 4436 98438
rect 4460 98436 4516 98438
rect 4880 97946 4936 97948
rect 4960 97946 5016 97948
rect 5040 97946 5096 97948
rect 5120 97946 5176 97948
rect 4880 97894 4926 97946
rect 4926 97894 4936 97946
rect 4960 97894 4990 97946
rect 4990 97894 5002 97946
rect 5002 97894 5016 97946
rect 5040 97894 5054 97946
rect 5054 97894 5066 97946
rect 5066 97894 5096 97946
rect 5120 97894 5130 97946
rect 5130 97894 5176 97946
rect 4880 97892 4936 97894
rect 4960 97892 5016 97894
rect 5040 97892 5096 97894
rect 5120 97892 5176 97894
rect 4220 97402 4276 97404
rect 4300 97402 4356 97404
rect 4380 97402 4436 97404
rect 4460 97402 4516 97404
rect 4220 97350 4266 97402
rect 4266 97350 4276 97402
rect 4300 97350 4330 97402
rect 4330 97350 4342 97402
rect 4342 97350 4356 97402
rect 4380 97350 4394 97402
rect 4394 97350 4406 97402
rect 4406 97350 4436 97402
rect 4460 97350 4470 97402
rect 4470 97350 4516 97402
rect 4220 97348 4276 97350
rect 4300 97348 4356 97350
rect 4380 97348 4436 97350
rect 4460 97348 4516 97350
rect 4880 96858 4936 96860
rect 4960 96858 5016 96860
rect 5040 96858 5096 96860
rect 5120 96858 5176 96860
rect 4880 96806 4926 96858
rect 4926 96806 4936 96858
rect 4960 96806 4990 96858
rect 4990 96806 5002 96858
rect 5002 96806 5016 96858
rect 5040 96806 5054 96858
rect 5054 96806 5066 96858
rect 5066 96806 5096 96858
rect 5120 96806 5130 96858
rect 5130 96806 5176 96858
rect 4880 96804 4936 96806
rect 4960 96804 5016 96806
rect 5040 96804 5096 96806
rect 5120 96804 5176 96806
rect 4220 96314 4276 96316
rect 4300 96314 4356 96316
rect 4380 96314 4436 96316
rect 4460 96314 4516 96316
rect 4220 96262 4266 96314
rect 4266 96262 4276 96314
rect 4300 96262 4330 96314
rect 4330 96262 4342 96314
rect 4342 96262 4356 96314
rect 4380 96262 4394 96314
rect 4394 96262 4406 96314
rect 4406 96262 4436 96314
rect 4460 96262 4470 96314
rect 4470 96262 4516 96314
rect 4220 96260 4276 96262
rect 4300 96260 4356 96262
rect 4380 96260 4436 96262
rect 4460 96260 4516 96262
rect 4880 95770 4936 95772
rect 4960 95770 5016 95772
rect 5040 95770 5096 95772
rect 5120 95770 5176 95772
rect 4880 95718 4926 95770
rect 4926 95718 4936 95770
rect 4960 95718 4990 95770
rect 4990 95718 5002 95770
rect 5002 95718 5016 95770
rect 5040 95718 5054 95770
rect 5054 95718 5066 95770
rect 5066 95718 5096 95770
rect 5120 95718 5130 95770
rect 5130 95718 5176 95770
rect 4880 95716 4936 95718
rect 4960 95716 5016 95718
rect 5040 95716 5096 95718
rect 5120 95716 5176 95718
rect 4220 95226 4276 95228
rect 4300 95226 4356 95228
rect 4380 95226 4436 95228
rect 4460 95226 4516 95228
rect 4220 95174 4266 95226
rect 4266 95174 4276 95226
rect 4300 95174 4330 95226
rect 4330 95174 4342 95226
rect 4342 95174 4356 95226
rect 4380 95174 4394 95226
rect 4394 95174 4406 95226
rect 4406 95174 4436 95226
rect 4460 95174 4470 95226
rect 4470 95174 4516 95226
rect 4220 95172 4276 95174
rect 4300 95172 4356 95174
rect 4380 95172 4436 95174
rect 4460 95172 4516 95174
rect 4880 94682 4936 94684
rect 4960 94682 5016 94684
rect 5040 94682 5096 94684
rect 5120 94682 5176 94684
rect 4880 94630 4926 94682
rect 4926 94630 4936 94682
rect 4960 94630 4990 94682
rect 4990 94630 5002 94682
rect 5002 94630 5016 94682
rect 5040 94630 5054 94682
rect 5054 94630 5066 94682
rect 5066 94630 5096 94682
rect 5120 94630 5130 94682
rect 5130 94630 5176 94682
rect 4880 94628 4936 94630
rect 4960 94628 5016 94630
rect 5040 94628 5096 94630
rect 5120 94628 5176 94630
rect 4220 94138 4276 94140
rect 4300 94138 4356 94140
rect 4380 94138 4436 94140
rect 4460 94138 4516 94140
rect 4220 94086 4266 94138
rect 4266 94086 4276 94138
rect 4300 94086 4330 94138
rect 4330 94086 4342 94138
rect 4342 94086 4356 94138
rect 4380 94086 4394 94138
rect 4394 94086 4406 94138
rect 4406 94086 4436 94138
rect 4460 94086 4470 94138
rect 4470 94086 4516 94138
rect 4220 94084 4276 94086
rect 4300 94084 4356 94086
rect 4380 94084 4436 94086
rect 4460 94084 4516 94086
rect 4880 93594 4936 93596
rect 4960 93594 5016 93596
rect 5040 93594 5096 93596
rect 5120 93594 5176 93596
rect 4880 93542 4926 93594
rect 4926 93542 4936 93594
rect 4960 93542 4990 93594
rect 4990 93542 5002 93594
rect 5002 93542 5016 93594
rect 5040 93542 5054 93594
rect 5054 93542 5066 93594
rect 5066 93542 5096 93594
rect 5120 93542 5130 93594
rect 5130 93542 5176 93594
rect 4880 93540 4936 93542
rect 4960 93540 5016 93542
rect 5040 93540 5096 93542
rect 5120 93540 5176 93542
rect 4220 93050 4276 93052
rect 4300 93050 4356 93052
rect 4380 93050 4436 93052
rect 4460 93050 4516 93052
rect 4220 92998 4266 93050
rect 4266 92998 4276 93050
rect 4300 92998 4330 93050
rect 4330 92998 4342 93050
rect 4342 92998 4356 93050
rect 4380 92998 4394 93050
rect 4394 92998 4406 93050
rect 4406 92998 4436 93050
rect 4460 92998 4470 93050
rect 4470 92998 4516 93050
rect 4220 92996 4276 92998
rect 4300 92996 4356 92998
rect 4380 92996 4436 92998
rect 4460 92996 4516 92998
rect 4880 92506 4936 92508
rect 4960 92506 5016 92508
rect 5040 92506 5096 92508
rect 5120 92506 5176 92508
rect 4880 92454 4926 92506
rect 4926 92454 4936 92506
rect 4960 92454 4990 92506
rect 4990 92454 5002 92506
rect 5002 92454 5016 92506
rect 5040 92454 5054 92506
rect 5054 92454 5066 92506
rect 5066 92454 5096 92506
rect 5120 92454 5130 92506
rect 5130 92454 5176 92506
rect 4880 92452 4936 92454
rect 4960 92452 5016 92454
rect 5040 92452 5096 92454
rect 5120 92452 5176 92454
rect 4220 91962 4276 91964
rect 4300 91962 4356 91964
rect 4380 91962 4436 91964
rect 4460 91962 4516 91964
rect 4220 91910 4266 91962
rect 4266 91910 4276 91962
rect 4300 91910 4330 91962
rect 4330 91910 4342 91962
rect 4342 91910 4356 91962
rect 4380 91910 4394 91962
rect 4394 91910 4406 91962
rect 4406 91910 4436 91962
rect 4460 91910 4470 91962
rect 4470 91910 4516 91962
rect 4220 91908 4276 91910
rect 4300 91908 4356 91910
rect 4380 91908 4436 91910
rect 4460 91908 4516 91910
rect 4880 91418 4936 91420
rect 4960 91418 5016 91420
rect 5040 91418 5096 91420
rect 5120 91418 5176 91420
rect 4880 91366 4926 91418
rect 4926 91366 4936 91418
rect 4960 91366 4990 91418
rect 4990 91366 5002 91418
rect 5002 91366 5016 91418
rect 5040 91366 5054 91418
rect 5054 91366 5066 91418
rect 5066 91366 5096 91418
rect 5120 91366 5130 91418
rect 5130 91366 5176 91418
rect 4880 91364 4936 91366
rect 4960 91364 5016 91366
rect 5040 91364 5096 91366
rect 5120 91364 5176 91366
rect 4220 90874 4276 90876
rect 4300 90874 4356 90876
rect 4380 90874 4436 90876
rect 4460 90874 4516 90876
rect 4220 90822 4266 90874
rect 4266 90822 4276 90874
rect 4300 90822 4330 90874
rect 4330 90822 4342 90874
rect 4342 90822 4356 90874
rect 4380 90822 4394 90874
rect 4394 90822 4406 90874
rect 4406 90822 4436 90874
rect 4460 90822 4470 90874
rect 4470 90822 4516 90874
rect 4220 90820 4276 90822
rect 4300 90820 4356 90822
rect 4380 90820 4436 90822
rect 4460 90820 4516 90822
rect 4880 90330 4936 90332
rect 4960 90330 5016 90332
rect 5040 90330 5096 90332
rect 5120 90330 5176 90332
rect 4880 90278 4926 90330
rect 4926 90278 4936 90330
rect 4960 90278 4990 90330
rect 4990 90278 5002 90330
rect 5002 90278 5016 90330
rect 5040 90278 5054 90330
rect 5054 90278 5066 90330
rect 5066 90278 5096 90330
rect 5120 90278 5130 90330
rect 5130 90278 5176 90330
rect 4880 90276 4936 90278
rect 4960 90276 5016 90278
rect 5040 90276 5096 90278
rect 5120 90276 5176 90278
rect 4220 89786 4276 89788
rect 4300 89786 4356 89788
rect 4380 89786 4436 89788
rect 4460 89786 4516 89788
rect 4220 89734 4266 89786
rect 4266 89734 4276 89786
rect 4300 89734 4330 89786
rect 4330 89734 4342 89786
rect 4342 89734 4356 89786
rect 4380 89734 4394 89786
rect 4394 89734 4406 89786
rect 4406 89734 4436 89786
rect 4460 89734 4470 89786
rect 4470 89734 4516 89786
rect 4220 89732 4276 89734
rect 4300 89732 4356 89734
rect 4380 89732 4436 89734
rect 4460 89732 4516 89734
rect 4880 89242 4936 89244
rect 4960 89242 5016 89244
rect 5040 89242 5096 89244
rect 5120 89242 5176 89244
rect 4880 89190 4926 89242
rect 4926 89190 4936 89242
rect 4960 89190 4990 89242
rect 4990 89190 5002 89242
rect 5002 89190 5016 89242
rect 5040 89190 5054 89242
rect 5054 89190 5066 89242
rect 5066 89190 5096 89242
rect 5120 89190 5130 89242
rect 5130 89190 5176 89242
rect 4880 89188 4936 89190
rect 4960 89188 5016 89190
rect 5040 89188 5096 89190
rect 5120 89188 5176 89190
rect 4220 88698 4276 88700
rect 4300 88698 4356 88700
rect 4380 88698 4436 88700
rect 4460 88698 4516 88700
rect 4220 88646 4266 88698
rect 4266 88646 4276 88698
rect 4300 88646 4330 88698
rect 4330 88646 4342 88698
rect 4342 88646 4356 88698
rect 4380 88646 4394 88698
rect 4394 88646 4406 88698
rect 4406 88646 4436 88698
rect 4460 88646 4470 88698
rect 4470 88646 4516 88698
rect 4220 88644 4276 88646
rect 4300 88644 4356 88646
rect 4380 88644 4436 88646
rect 4460 88644 4516 88646
rect 1306 88440 1362 88496
rect 4880 88154 4936 88156
rect 4960 88154 5016 88156
rect 5040 88154 5096 88156
rect 5120 88154 5176 88156
rect 4880 88102 4926 88154
rect 4926 88102 4936 88154
rect 4960 88102 4990 88154
rect 4990 88102 5002 88154
rect 5002 88102 5016 88154
rect 5040 88102 5054 88154
rect 5054 88102 5066 88154
rect 5066 88102 5096 88154
rect 5120 88102 5130 88154
rect 5130 88102 5176 88154
rect 4880 88100 4936 88102
rect 4960 88100 5016 88102
rect 5040 88100 5096 88102
rect 5120 88100 5176 88102
rect 1214 87760 1270 87816
rect 4220 87610 4276 87612
rect 4300 87610 4356 87612
rect 4380 87610 4436 87612
rect 4460 87610 4516 87612
rect 4220 87558 4266 87610
rect 4266 87558 4276 87610
rect 4300 87558 4330 87610
rect 4330 87558 4342 87610
rect 4342 87558 4356 87610
rect 4380 87558 4394 87610
rect 4394 87558 4406 87610
rect 4406 87558 4436 87610
rect 4460 87558 4470 87610
rect 4470 87558 4516 87610
rect 4220 87556 4276 87558
rect 4300 87556 4356 87558
rect 4380 87556 4436 87558
rect 4460 87556 4516 87558
rect 1214 87080 1270 87136
rect 1306 86400 1362 86456
rect 4880 87066 4936 87068
rect 4960 87066 5016 87068
rect 5040 87066 5096 87068
rect 5120 87066 5176 87068
rect 4880 87014 4926 87066
rect 4926 87014 4936 87066
rect 4960 87014 4990 87066
rect 4990 87014 5002 87066
rect 5002 87014 5016 87066
rect 5040 87014 5054 87066
rect 5054 87014 5066 87066
rect 5066 87014 5096 87066
rect 5120 87014 5130 87066
rect 5130 87014 5176 87066
rect 4880 87012 4936 87014
rect 4960 87012 5016 87014
rect 5040 87012 5096 87014
rect 5120 87012 5176 87014
rect 4220 86522 4276 86524
rect 4300 86522 4356 86524
rect 4380 86522 4436 86524
rect 4460 86522 4516 86524
rect 4220 86470 4266 86522
rect 4266 86470 4276 86522
rect 4300 86470 4330 86522
rect 4330 86470 4342 86522
rect 4342 86470 4356 86522
rect 4380 86470 4394 86522
rect 4394 86470 4406 86522
rect 4406 86470 4436 86522
rect 4460 86470 4470 86522
rect 4470 86470 4516 86522
rect 4220 86468 4276 86470
rect 4300 86468 4356 86470
rect 4380 86468 4436 86470
rect 4460 86468 4516 86470
rect 4880 85978 4936 85980
rect 4960 85978 5016 85980
rect 5040 85978 5096 85980
rect 5120 85978 5176 85980
rect 4880 85926 4926 85978
rect 4926 85926 4936 85978
rect 4960 85926 4990 85978
rect 4990 85926 5002 85978
rect 5002 85926 5016 85978
rect 5040 85926 5054 85978
rect 5054 85926 5066 85978
rect 5066 85926 5096 85978
rect 5120 85926 5130 85978
rect 5130 85926 5176 85978
rect 4880 85924 4936 85926
rect 4960 85924 5016 85926
rect 5040 85924 5096 85926
rect 5120 85924 5176 85926
rect 1306 85720 1362 85776
rect 5998 85448 6054 85504
rect 4220 85434 4276 85436
rect 4300 85434 4356 85436
rect 4380 85434 4436 85436
rect 4460 85434 4516 85436
rect 4220 85382 4266 85434
rect 4266 85382 4276 85434
rect 4300 85382 4330 85434
rect 4330 85382 4342 85434
rect 4342 85382 4356 85434
rect 4380 85382 4394 85434
rect 4394 85382 4406 85434
rect 4406 85382 4436 85434
rect 4460 85382 4470 85434
rect 4470 85382 4516 85434
rect 4220 85380 4276 85382
rect 4300 85380 4356 85382
rect 4380 85380 4436 85382
rect 4460 85380 4516 85382
rect 1214 85060 1270 85096
rect 1214 85040 1216 85060
rect 1216 85040 1268 85060
rect 1268 85040 1270 85060
rect 1306 84360 1362 84416
rect 4880 84890 4936 84892
rect 4960 84890 5016 84892
rect 5040 84890 5096 84892
rect 5120 84890 5176 84892
rect 4880 84838 4926 84890
rect 4926 84838 4936 84890
rect 4960 84838 4990 84890
rect 4990 84838 5002 84890
rect 5002 84838 5016 84890
rect 5040 84838 5054 84890
rect 5054 84838 5066 84890
rect 5066 84838 5096 84890
rect 5120 84838 5130 84890
rect 5130 84838 5176 84890
rect 4880 84836 4936 84838
rect 4960 84836 5016 84838
rect 5040 84836 5096 84838
rect 5120 84836 5176 84838
rect 4220 84346 4276 84348
rect 4300 84346 4356 84348
rect 4380 84346 4436 84348
rect 4460 84346 4516 84348
rect 4220 84294 4266 84346
rect 4266 84294 4276 84346
rect 4300 84294 4330 84346
rect 4330 84294 4342 84346
rect 4342 84294 4356 84346
rect 4380 84294 4394 84346
rect 4394 84294 4406 84346
rect 4406 84294 4436 84346
rect 4460 84294 4470 84346
rect 4470 84294 4516 84346
rect 4220 84292 4276 84294
rect 4300 84292 4356 84294
rect 4380 84292 4436 84294
rect 4460 84292 4516 84294
rect 1306 83680 1362 83736
rect 1306 83000 1362 83056
rect 4880 83802 4936 83804
rect 4960 83802 5016 83804
rect 5040 83802 5096 83804
rect 5120 83802 5176 83804
rect 4880 83750 4926 83802
rect 4926 83750 4936 83802
rect 4960 83750 4990 83802
rect 4990 83750 5002 83802
rect 5002 83750 5016 83802
rect 5040 83750 5054 83802
rect 5054 83750 5066 83802
rect 5066 83750 5096 83802
rect 5120 83750 5130 83802
rect 5130 83750 5176 83802
rect 4880 83748 4936 83750
rect 4960 83748 5016 83750
rect 5040 83748 5096 83750
rect 5120 83748 5176 83750
rect 1214 82320 1270 82376
rect 1214 81640 1270 81696
rect 1306 80960 1362 81016
rect 4220 83258 4276 83260
rect 4300 83258 4356 83260
rect 4380 83258 4436 83260
rect 4460 83258 4516 83260
rect 4220 83206 4266 83258
rect 4266 83206 4276 83258
rect 4300 83206 4330 83258
rect 4330 83206 4342 83258
rect 4342 83206 4356 83258
rect 4380 83206 4394 83258
rect 4394 83206 4406 83258
rect 4406 83206 4436 83258
rect 4460 83206 4470 83258
rect 4470 83206 4516 83258
rect 4220 83204 4276 83206
rect 4300 83204 4356 83206
rect 4380 83204 4436 83206
rect 4460 83204 4516 83206
rect 4880 82714 4936 82716
rect 4960 82714 5016 82716
rect 5040 82714 5096 82716
rect 5120 82714 5176 82716
rect 4880 82662 4926 82714
rect 4926 82662 4936 82714
rect 4960 82662 4990 82714
rect 4990 82662 5002 82714
rect 5002 82662 5016 82714
rect 5040 82662 5054 82714
rect 5054 82662 5066 82714
rect 5066 82662 5096 82714
rect 5120 82662 5130 82714
rect 5130 82662 5176 82714
rect 4880 82660 4936 82662
rect 4960 82660 5016 82662
rect 5040 82660 5096 82662
rect 5120 82660 5176 82662
rect 4220 82170 4276 82172
rect 4300 82170 4356 82172
rect 4380 82170 4436 82172
rect 4460 82170 4516 82172
rect 4220 82118 4266 82170
rect 4266 82118 4276 82170
rect 4300 82118 4330 82170
rect 4330 82118 4342 82170
rect 4342 82118 4356 82170
rect 4380 82118 4394 82170
rect 4394 82118 4406 82170
rect 4406 82118 4436 82170
rect 4460 82118 4470 82170
rect 4470 82118 4516 82170
rect 4220 82116 4276 82118
rect 4300 82116 4356 82118
rect 4380 82116 4436 82118
rect 4460 82116 4516 82118
rect 4880 81626 4936 81628
rect 4960 81626 5016 81628
rect 5040 81626 5096 81628
rect 5120 81626 5176 81628
rect 4880 81574 4926 81626
rect 4926 81574 4936 81626
rect 4960 81574 4990 81626
rect 4990 81574 5002 81626
rect 5002 81574 5016 81626
rect 5040 81574 5054 81626
rect 5054 81574 5066 81626
rect 5066 81574 5096 81626
rect 5120 81574 5130 81626
rect 5130 81574 5176 81626
rect 4880 81572 4936 81574
rect 4960 81572 5016 81574
rect 5040 81572 5096 81574
rect 5120 81572 5176 81574
rect 4220 81082 4276 81084
rect 4300 81082 4356 81084
rect 4380 81082 4436 81084
rect 4460 81082 4516 81084
rect 4220 81030 4266 81082
rect 4266 81030 4276 81082
rect 4300 81030 4330 81082
rect 4330 81030 4342 81082
rect 4342 81030 4356 81082
rect 4380 81030 4394 81082
rect 4394 81030 4406 81082
rect 4406 81030 4436 81082
rect 4460 81030 4470 81082
rect 4470 81030 4516 81082
rect 4220 81028 4276 81030
rect 4300 81028 4356 81030
rect 4380 81028 4436 81030
rect 4460 81028 4516 81030
rect 4880 80538 4936 80540
rect 4960 80538 5016 80540
rect 5040 80538 5096 80540
rect 5120 80538 5176 80540
rect 4880 80486 4926 80538
rect 4926 80486 4936 80538
rect 4960 80486 4990 80538
rect 4990 80486 5002 80538
rect 5002 80486 5016 80538
rect 5040 80486 5054 80538
rect 5054 80486 5066 80538
rect 5066 80486 5096 80538
rect 5120 80486 5130 80538
rect 5130 80486 5176 80538
rect 4880 80484 4936 80486
rect 4960 80484 5016 80486
rect 5040 80484 5096 80486
rect 5120 80484 5176 80486
rect 1306 80316 1308 80336
rect 1308 80316 1360 80336
rect 1360 80316 1362 80336
rect 1306 80280 1362 80316
rect 4220 79994 4276 79996
rect 4300 79994 4356 79996
rect 4380 79994 4436 79996
rect 4460 79994 4516 79996
rect 4220 79942 4266 79994
rect 4266 79942 4276 79994
rect 4300 79942 4330 79994
rect 4330 79942 4342 79994
rect 4342 79942 4356 79994
rect 4380 79942 4394 79994
rect 4394 79942 4406 79994
rect 4406 79942 4436 79994
rect 4460 79942 4470 79994
rect 4470 79942 4516 79994
rect 4220 79940 4276 79942
rect 4300 79940 4356 79942
rect 4380 79940 4436 79942
rect 4460 79940 4516 79942
rect 1214 79620 1270 79656
rect 1214 79600 1216 79620
rect 1216 79600 1268 79620
rect 1268 79600 1270 79620
rect 5630 79600 5686 79656
rect 5538 79464 5594 79520
rect 4880 79450 4936 79452
rect 4960 79450 5016 79452
rect 5040 79450 5096 79452
rect 5120 79450 5176 79452
rect 4880 79398 4926 79450
rect 4926 79398 4936 79450
rect 4960 79398 4990 79450
rect 4990 79398 5002 79450
rect 5002 79398 5016 79450
rect 5040 79398 5054 79450
rect 5054 79398 5066 79450
rect 5066 79398 5096 79450
rect 5120 79398 5130 79450
rect 5130 79398 5176 79450
rect 4880 79396 4936 79398
rect 4960 79396 5016 79398
rect 5040 79396 5096 79398
rect 5120 79396 5176 79398
rect 7562 79192 7618 79248
rect 1306 78920 1362 78976
rect 4220 78906 4276 78908
rect 4300 78906 4356 78908
rect 4380 78906 4436 78908
rect 4460 78906 4516 78908
rect 4220 78854 4266 78906
rect 4266 78854 4276 78906
rect 4300 78854 4330 78906
rect 4330 78854 4342 78906
rect 4342 78854 4356 78906
rect 4380 78854 4394 78906
rect 4394 78854 4406 78906
rect 4406 78854 4436 78906
rect 4460 78854 4470 78906
rect 4470 78854 4516 78906
rect 4220 78852 4276 78854
rect 4300 78852 4356 78854
rect 4380 78852 4436 78854
rect 4460 78852 4516 78854
rect 4880 78362 4936 78364
rect 4960 78362 5016 78364
rect 5040 78362 5096 78364
rect 5120 78362 5176 78364
rect 4880 78310 4926 78362
rect 4926 78310 4936 78362
rect 4960 78310 4990 78362
rect 4990 78310 5002 78362
rect 5002 78310 5016 78362
rect 5040 78310 5054 78362
rect 5054 78310 5066 78362
rect 5066 78310 5096 78362
rect 5120 78310 5130 78362
rect 5130 78310 5176 78362
rect 4880 78308 4936 78310
rect 4960 78308 5016 78310
rect 5040 78308 5096 78310
rect 5120 78308 5176 78310
rect 1306 78240 1362 78296
rect 1306 77560 1362 77616
rect 1214 76880 1270 76936
rect 846 76336 902 76392
rect 1398 75520 1454 75576
rect 846 74976 902 75032
rect 846 74332 848 74352
rect 848 74332 900 74352
rect 900 74332 902 74352
rect 846 74296 902 74332
rect 846 73636 902 73672
rect 846 73616 848 73636
rect 848 73616 900 73636
rect 900 73616 902 73636
rect 4220 77818 4276 77820
rect 4300 77818 4356 77820
rect 4380 77818 4436 77820
rect 4460 77818 4516 77820
rect 4220 77766 4266 77818
rect 4266 77766 4276 77818
rect 4300 77766 4330 77818
rect 4330 77766 4342 77818
rect 4342 77766 4356 77818
rect 4380 77766 4394 77818
rect 4394 77766 4406 77818
rect 4406 77766 4436 77818
rect 4460 77766 4470 77818
rect 4470 77766 4516 77818
rect 4220 77764 4276 77766
rect 4300 77764 4356 77766
rect 4380 77764 4436 77766
rect 4460 77764 4516 77766
rect 8022 78512 8078 78568
rect 8390 111152 8446 111208
rect 8390 109540 8446 109576
rect 8390 109520 8392 109540
rect 8392 109520 8444 109540
rect 8444 109520 8446 109540
rect 8390 108452 8446 108488
rect 8390 108432 8392 108452
rect 8392 108432 8444 108452
rect 8444 108432 8446 108452
rect 8390 106664 8446 106720
rect 8390 105576 8446 105632
rect 8390 103944 8446 104000
rect 8482 79872 8538 79928
rect 8666 79736 8722 79792
rect 9402 79328 9458 79384
rect 8206 78104 8262 78160
rect 8114 77832 8170 77888
rect 7930 77696 7986 77752
rect 35600 136026 35656 136028
rect 35680 136026 35736 136028
rect 35760 136026 35816 136028
rect 35840 136026 35896 136028
rect 35600 135974 35646 136026
rect 35646 135974 35656 136026
rect 35680 135974 35710 136026
rect 35710 135974 35722 136026
rect 35722 135974 35736 136026
rect 35760 135974 35774 136026
rect 35774 135974 35786 136026
rect 35786 135974 35816 136026
rect 35840 135974 35850 136026
rect 35850 135974 35896 136026
rect 35600 135972 35656 135974
rect 35680 135972 35736 135974
rect 35760 135972 35816 135974
rect 35840 135972 35896 135974
rect 38198 134136 38254 134192
rect 40682 134136 40738 134192
rect 52366 134136 52422 134192
rect 60646 135224 60702 135280
rect 63130 135224 63186 135280
rect 66320 136026 66376 136028
rect 66400 136026 66456 136028
rect 66480 136026 66536 136028
rect 66560 136026 66616 136028
rect 66320 135974 66366 136026
rect 66366 135974 66376 136026
rect 66400 135974 66430 136026
rect 66430 135974 66442 136026
rect 66442 135974 66456 136026
rect 66480 135974 66494 136026
rect 66494 135974 66506 136026
rect 66506 135974 66536 136026
rect 66560 135974 66570 136026
rect 66570 135974 66616 136026
rect 66320 135972 66376 135974
rect 66400 135972 66456 135974
rect 66480 135972 66536 135974
rect 66560 135972 66616 135974
rect 67546 135224 67602 135280
rect 69754 135224 69810 135280
rect 72146 135224 72202 135280
rect 64418 135088 64474 135144
rect 58162 134136 58218 134192
rect 74170 134136 74226 134192
rect 55770 134000 55826 134056
rect 97040 136026 97096 136028
rect 97120 136026 97176 136028
rect 97200 136026 97256 136028
rect 97280 136026 97336 136028
rect 97040 135974 97086 136026
rect 97086 135974 97096 136026
rect 97120 135974 97150 136026
rect 97150 135974 97162 136026
rect 97162 135974 97176 136026
rect 97200 135974 97214 136026
rect 97214 135974 97226 136026
rect 97226 135974 97256 136026
rect 97280 135974 97290 136026
rect 97290 135974 97336 136026
rect 97040 135972 97096 135974
rect 97120 135972 97176 135974
rect 97200 135972 97256 135974
rect 97280 135972 97336 135974
rect 95974 134408 96030 134464
rect 36082 133900 36084 133920
rect 36084 133900 36136 133920
rect 36136 133900 36138 133920
rect 36082 133864 36138 133900
rect 42982 133864 43038 133920
rect 46018 133864 46074 133920
rect 48502 133864 48558 133920
rect 86130 133900 86132 133920
rect 86132 133900 86184 133920
rect 86184 133900 86186 133920
rect 86130 133864 86186 133900
rect 87326 133864 87382 133920
rect 36266 79872 36322 79928
rect 38658 79892 38714 79928
rect 38658 79872 38660 79892
rect 38660 79872 38712 79892
rect 38712 79872 38714 79892
rect 39762 79908 39764 79928
rect 39764 79908 39816 79928
rect 39816 79908 39818 79928
rect 39762 79872 39818 79908
rect 40958 79872 41014 79928
rect 90638 79872 90694 79928
rect 32310 79736 32366 79792
rect 27618 79600 27674 79656
rect 24674 79464 24730 79520
rect 9586 78240 9642 78296
rect 16026 77968 16082 78024
rect 9494 77560 9550 77616
rect 4880 77274 4936 77276
rect 4960 77274 5016 77276
rect 5040 77274 5096 77276
rect 5120 77274 5176 77276
rect 4880 77222 4926 77274
rect 4926 77222 4936 77274
rect 4960 77222 4990 77274
rect 4990 77222 5002 77274
rect 5002 77222 5016 77274
rect 5040 77222 5054 77274
rect 5054 77222 5066 77274
rect 5066 77222 5096 77274
rect 5120 77222 5130 77274
rect 5130 77222 5176 77274
rect 4880 77220 4936 77222
rect 4960 77220 5016 77222
rect 5040 77220 5096 77222
rect 5120 77220 5176 77222
rect 4220 76730 4276 76732
rect 4300 76730 4356 76732
rect 4380 76730 4436 76732
rect 4460 76730 4516 76732
rect 4220 76678 4266 76730
rect 4266 76678 4276 76730
rect 4300 76678 4330 76730
rect 4330 76678 4342 76730
rect 4342 76678 4356 76730
rect 4380 76678 4394 76730
rect 4394 76678 4406 76730
rect 4406 76678 4436 76730
rect 4460 76678 4470 76730
rect 4470 76678 4516 76730
rect 4220 76676 4276 76678
rect 4300 76676 4356 76678
rect 4380 76676 4436 76678
rect 4460 76676 4516 76678
rect 4880 76186 4936 76188
rect 4960 76186 5016 76188
rect 5040 76186 5096 76188
rect 5120 76186 5176 76188
rect 4880 76134 4926 76186
rect 4926 76134 4936 76186
rect 4960 76134 4990 76186
rect 4990 76134 5002 76186
rect 5002 76134 5016 76186
rect 5040 76134 5054 76186
rect 5054 76134 5066 76186
rect 5066 76134 5096 76186
rect 5120 76134 5130 76186
rect 5130 76134 5176 76186
rect 4880 76132 4936 76134
rect 4960 76132 5016 76134
rect 5040 76132 5096 76134
rect 5120 76132 5176 76134
rect 4220 75642 4276 75644
rect 4300 75642 4356 75644
rect 4380 75642 4436 75644
rect 4460 75642 4516 75644
rect 4220 75590 4266 75642
rect 4266 75590 4276 75642
rect 4300 75590 4330 75642
rect 4330 75590 4342 75642
rect 4342 75590 4356 75642
rect 4380 75590 4394 75642
rect 4394 75590 4406 75642
rect 4406 75590 4436 75642
rect 4460 75590 4470 75642
rect 4470 75590 4516 75642
rect 4220 75588 4276 75590
rect 4300 75588 4356 75590
rect 4380 75588 4436 75590
rect 4460 75588 4516 75590
rect 4880 75098 4936 75100
rect 4960 75098 5016 75100
rect 5040 75098 5096 75100
rect 5120 75098 5176 75100
rect 4880 75046 4926 75098
rect 4926 75046 4936 75098
rect 4960 75046 4990 75098
rect 4990 75046 5002 75098
rect 5002 75046 5016 75098
rect 5040 75046 5054 75098
rect 5054 75046 5066 75098
rect 5066 75046 5096 75098
rect 5120 75046 5130 75098
rect 5130 75046 5176 75098
rect 4880 75044 4936 75046
rect 4960 75044 5016 75046
rect 5040 75044 5096 75046
rect 5120 75044 5176 75046
rect 4220 74554 4276 74556
rect 4300 74554 4356 74556
rect 4380 74554 4436 74556
rect 4460 74554 4516 74556
rect 4220 74502 4266 74554
rect 4266 74502 4276 74554
rect 4300 74502 4330 74554
rect 4330 74502 4342 74554
rect 4342 74502 4356 74554
rect 4380 74502 4394 74554
rect 4394 74502 4406 74554
rect 4406 74502 4436 74554
rect 4460 74502 4470 74554
rect 4470 74502 4516 74554
rect 4220 74500 4276 74502
rect 4300 74500 4356 74502
rect 4380 74500 4436 74502
rect 4460 74500 4516 74502
rect 4880 74010 4936 74012
rect 4960 74010 5016 74012
rect 5040 74010 5096 74012
rect 5120 74010 5176 74012
rect 4880 73958 4926 74010
rect 4926 73958 4936 74010
rect 4960 73958 4990 74010
rect 4990 73958 5002 74010
rect 5002 73958 5016 74010
rect 5040 73958 5054 74010
rect 5054 73958 5066 74010
rect 5066 73958 5096 74010
rect 5120 73958 5130 74010
rect 5130 73958 5176 74010
rect 4880 73956 4936 73958
rect 4960 73956 5016 73958
rect 5040 73956 5096 73958
rect 5120 73956 5176 73958
rect 4220 73466 4276 73468
rect 4300 73466 4356 73468
rect 4380 73466 4436 73468
rect 4460 73466 4516 73468
rect 4220 73414 4266 73466
rect 4266 73414 4276 73466
rect 4300 73414 4330 73466
rect 4330 73414 4342 73466
rect 4342 73414 4356 73466
rect 4380 73414 4394 73466
rect 4394 73414 4406 73466
rect 4406 73414 4436 73466
rect 4460 73414 4470 73466
rect 4470 73414 4516 73466
rect 4220 73412 4276 73414
rect 4300 73412 4356 73414
rect 4380 73412 4436 73414
rect 4460 73412 4516 73414
rect 846 72972 848 72992
rect 848 72972 900 72992
rect 900 72972 902 72992
rect 846 72936 902 72972
rect 4880 72922 4936 72924
rect 4960 72922 5016 72924
rect 5040 72922 5096 72924
rect 5120 72922 5176 72924
rect 4880 72870 4926 72922
rect 4926 72870 4936 72922
rect 4960 72870 4990 72922
rect 4990 72870 5002 72922
rect 5002 72870 5016 72922
rect 5040 72870 5054 72922
rect 5054 72870 5066 72922
rect 5066 72870 5096 72922
rect 5120 72870 5130 72922
rect 5130 72870 5176 72922
rect 4880 72868 4936 72870
rect 4960 72868 5016 72870
rect 5040 72868 5096 72870
rect 5120 72868 5176 72870
rect 4220 72378 4276 72380
rect 4300 72378 4356 72380
rect 4380 72378 4436 72380
rect 4460 72378 4516 72380
rect 4220 72326 4266 72378
rect 4266 72326 4276 72378
rect 4300 72326 4330 72378
rect 4330 72326 4342 72378
rect 4342 72326 4356 72378
rect 4380 72326 4394 72378
rect 4394 72326 4406 72378
rect 4406 72326 4436 72378
rect 4460 72326 4470 72378
rect 4470 72326 4516 72378
rect 4220 72324 4276 72326
rect 4300 72324 4356 72326
rect 4380 72324 4436 72326
rect 4460 72324 4516 72326
rect 1122 72120 1178 72176
rect 4880 71834 4936 71836
rect 4960 71834 5016 71836
rect 5040 71834 5096 71836
rect 5120 71834 5176 71836
rect 4880 71782 4926 71834
rect 4926 71782 4936 71834
rect 4960 71782 4990 71834
rect 4990 71782 5002 71834
rect 5002 71782 5016 71834
rect 5040 71782 5054 71834
rect 5054 71782 5066 71834
rect 5066 71782 5096 71834
rect 5120 71782 5130 71834
rect 5130 71782 5176 71834
rect 4880 71780 4936 71782
rect 4960 71780 5016 71782
rect 5040 71780 5096 71782
rect 5120 71780 5176 71782
rect 4220 71290 4276 71292
rect 4300 71290 4356 71292
rect 4380 71290 4436 71292
rect 4460 71290 4516 71292
rect 4220 71238 4266 71290
rect 4266 71238 4276 71290
rect 4300 71238 4330 71290
rect 4330 71238 4342 71290
rect 4342 71238 4356 71290
rect 4380 71238 4394 71290
rect 4394 71238 4406 71290
rect 4406 71238 4436 71290
rect 4460 71238 4470 71290
rect 4470 71238 4516 71290
rect 4220 71236 4276 71238
rect 4300 71236 4356 71238
rect 4380 71236 4436 71238
rect 4460 71236 4516 71238
rect 4880 70746 4936 70748
rect 4960 70746 5016 70748
rect 5040 70746 5096 70748
rect 5120 70746 5176 70748
rect 4880 70694 4926 70746
rect 4926 70694 4936 70746
rect 4960 70694 4990 70746
rect 4990 70694 5002 70746
rect 5002 70694 5016 70746
rect 5040 70694 5054 70746
rect 5054 70694 5066 70746
rect 5066 70694 5096 70746
rect 5120 70694 5130 70746
rect 5130 70694 5176 70746
rect 4880 70692 4936 70694
rect 4960 70692 5016 70694
rect 5040 70692 5096 70694
rect 5120 70692 5176 70694
rect 4220 70202 4276 70204
rect 4300 70202 4356 70204
rect 4380 70202 4436 70204
rect 4460 70202 4516 70204
rect 4220 70150 4266 70202
rect 4266 70150 4276 70202
rect 4300 70150 4330 70202
rect 4330 70150 4342 70202
rect 4342 70150 4356 70202
rect 4380 70150 4394 70202
rect 4394 70150 4406 70202
rect 4406 70150 4436 70202
rect 4460 70150 4470 70202
rect 4470 70150 4516 70202
rect 4220 70148 4276 70150
rect 4300 70148 4356 70150
rect 4380 70148 4436 70150
rect 4460 70148 4516 70150
rect 4880 69658 4936 69660
rect 4960 69658 5016 69660
rect 5040 69658 5096 69660
rect 5120 69658 5176 69660
rect 4880 69606 4926 69658
rect 4926 69606 4936 69658
rect 4960 69606 4990 69658
rect 4990 69606 5002 69658
rect 5002 69606 5016 69658
rect 5040 69606 5054 69658
rect 5054 69606 5066 69658
rect 5066 69606 5096 69658
rect 5120 69606 5130 69658
rect 5130 69606 5176 69658
rect 4880 69604 4936 69606
rect 4960 69604 5016 69606
rect 5040 69604 5096 69606
rect 5120 69604 5176 69606
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 4880 68570 4936 68572
rect 4960 68570 5016 68572
rect 5040 68570 5096 68572
rect 5120 68570 5176 68572
rect 4880 68518 4926 68570
rect 4926 68518 4936 68570
rect 4960 68518 4990 68570
rect 4990 68518 5002 68570
rect 5002 68518 5016 68570
rect 5040 68518 5054 68570
rect 5054 68518 5066 68570
rect 5066 68518 5096 68570
rect 5120 68518 5130 68570
rect 5130 68518 5176 68570
rect 4880 68516 4936 68518
rect 4960 68516 5016 68518
rect 5040 68516 5096 68518
rect 5120 68516 5176 68518
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 4880 67482 4936 67484
rect 4960 67482 5016 67484
rect 5040 67482 5096 67484
rect 5120 67482 5176 67484
rect 4880 67430 4926 67482
rect 4926 67430 4936 67482
rect 4960 67430 4990 67482
rect 4990 67430 5002 67482
rect 5002 67430 5016 67482
rect 5040 67430 5054 67482
rect 5054 67430 5066 67482
rect 5066 67430 5096 67482
rect 5120 67430 5130 67482
rect 5130 67430 5176 67482
rect 4880 67428 4936 67430
rect 4960 67428 5016 67430
rect 5040 67428 5096 67430
rect 5120 67428 5176 67430
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 4880 66394 4936 66396
rect 4960 66394 5016 66396
rect 5040 66394 5096 66396
rect 5120 66394 5176 66396
rect 4880 66342 4926 66394
rect 4926 66342 4936 66394
rect 4960 66342 4990 66394
rect 4990 66342 5002 66394
rect 5002 66342 5016 66394
rect 5040 66342 5054 66394
rect 5054 66342 5066 66394
rect 5066 66342 5096 66394
rect 5120 66342 5130 66394
rect 5130 66342 5176 66394
rect 4880 66340 4936 66342
rect 4960 66340 5016 66342
rect 5040 66340 5096 66342
rect 5120 66340 5176 66342
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 4880 65306 4936 65308
rect 4960 65306 5016 65308
rect 5040 65306 5096 65308
rect 5120 65306 5176 65308
rect 4880 65254 4926 65306
rect 4926 65254 4936 65306
rect 4960 65254 4990 65306
rect 4990 65254 5002 65306
rect 5002 65254 5016 65306
rect 5040 65254 5054 65306
rect 5054 65254 5066 65306
rect 5066 65254 5096 65306
rect 5120 65254 5130 65306
rect 5130 65254 5176 65306
rect 4880 65252 4936 65254
rect 4960 65252 5016 65254
rect 5040 65252 5096 65254
rect 5120 65252 5176 65254
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 4880 64218 4936 64220
rect 4960 64218 5016 64220
rect 5040 64218 5096 64220
rect 5120 64218 5176 64220
rect 4880 64166 4926 64218
rect 4926 64166 4936 64218
rect 4960 64166 4990 64218
rect 4990 64166 5002 64218
rect 5002 64166 5016 64218
rect 5040 64166 5054 64218
rect 5054 64166 5066 64218
rect 5066 64166 5096 64218
rect 5120 64166 5130 64218
rect 5130 64166 5176 64218
rect 4880 64164 4936 64166
rect 4960 64164 5016 64166
rect 5040 64164 5096 64166
rect 5120 64164 5176 64166
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 4880 63130 4936 63132
rect 4960 63130 5016 63132
rect 5040 63130 5096 63132
rect 5120 63130 5176 63132
rect 4880 63078 4926 63130
rect 4926 63078 4936 63130
rect 4960 63078 4990 63130
rect 4990 63078 5002 63130
rect 5002 63078 5016 63130
rect 5040 63078 5054 63130
rect 5054 63078 5066 63130
rect 5066 63078 5096 63130
rect 5120 63078 5130 63130
rect 5130 63078 5176 63130
rect 4880 63076 4936 63078
rect 4960 63076 5016 63078
rect 5040 63076 5096 63078
rect 5120 63076 5176 63078
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 4880 62042 4936 62044
rect 4960 62042 5016 62044
rect 5040 62042 5096 62044
rect 5120 62042 5176 62044
rect 4880 61990 4926 62042
rect 4926 61990 4936 62042
rect 4960 61990 4990 62042
rect 4990 61990 5002 62042
rect 5002 61990 5016 62042
rect 5040 61990 5054 62042
rect 5054 61990 5066 62042
rect 5066 61990 5096 62042
rect 5120 61990 5130 62042
rect 5130 61990 5176 62042
rect 4880 61988 4936 61990
rect 4960 61988 5016 61990
rect 5040 61988 5096 61990
rect 5120 61988 5176 61990
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 4880 60954 4936 60956
rect 4960 60954 5016 60956
rect 5040 60954 5096 60956
rect 5120 60954 5176 60956
rect 4880 60902 4926 60954
rect 4926 60902 4936 60954
rect 4960 60902 4990 60954
rect 4990 60902 5002 60954
rect 5002 60902 5016 60954
rect 5040 60902 5054 60954
rect 5054 60902 5066 60954
rect 5066 60902 5096 60954
rect 5120 60902 5130 60954
rect 5130 60902 5176 60954
rect 4880 60900 4936 60902
rect 4960 60900 5016 60902
rect 5040 60900 5096 60902
rect 5120 60900 5176 60902
rect 26790 79328 26846 79384
rect 24766 78784 24822 78840
rect 29550 79464 29606 79520
rect 30470 79464 30526 79520
rect 31574 79464 31630 79520
rect 28170 77716 28226 77752
rect 28170 77696 28172 77716
rect 28172 77696 28224 77716
rect 28224 77696 28226 77716
rect 31206 77832 31262 77888
rect 33966 79464 34022 79520
rect 34702 79464 34758 79520
rect 32954 78512 33010 78568
rect 35346 78240 35402 78296
rect 34940 77818 34996 77820
rect 35020 77818 35076 77820
rect 35100 77818 35156 77820
rect 35180 77818 35236 77820
rect 34940 77766 34986 77818
rect 34986 77766 34996 77818
rect 35020 77766 35050 77818
rect 35050 77766 35062 77818
rect 35062 77766 35076 77818
rect 35100 77766 35114 77818
rect 35114 77766 35126 77818
rect 35126 77766 35156 77818
rect 35180 77766 35190 77818
rect 35190 77766 35236 77818
rect 34940 77764 34996 77766
rect 35020 77764 35076 77766
rect 35100 77764 35156 77766
rect 35180 77764 35236 77766
rect 35990 77324 35992 77344
rect 35992 77324 36044 77344
rect 36044 77324 36046 77344
rect 35990 77288 36046 77324
rect 35600 77274 35656 77276
rect 35680 77274 35736 77276
rect 35760 77274 35816 77276
rect 35840 77274 35896 77276
rect 35600 77222 35646 77274
rect 35646 77222 35656 77274
rect 35680 77222 35710 77274
rect 35710 77222 35722 77274
rect 35722 77222 35736 77274
rect 35760 77222 35774 77274
rect 35774 77222 35786 77274
rect 35786 77222 35816 77274
rect 35840 77222 35850 77274
rect 35850 77222 35896 77274
rect 35600 77220 35656 77222
rect 35680 77220 35736 77222
rect 35760 77220 35816 77222
rect 35840 77220 35896 77222
rect 34940 76730 34996 76732
rect 35020 76730 35076 76732
rect 35100 76730 35156 76732
rect 35180 76730 35236 76732
rect 34940 76678 34986 76730
rect 34986 76678 34996 76730
rect 35020 76678 35050 76730
rect 35050 76678 35062 76730
rect 35062 76678 35076 76730
rect 35100 76678 35114 76730
rect 35114 76678 35126 76730
rect 35126 76678 35156 76730
rect 35180 76678 35190 76730
rect 35190 76678 35236 76730
rect 34940 76676 34996 76678
rect 35020 76676 35076 76678
rect 35100 76676 35156 76678
rect 35180 76676 35236 76678
rect 35600 76186 35656 76188
rect 35680 76186 35736 76188
rect 35760 76186 35816 76188
rect 35840 76186 35896 76188
rect 35600 76134 35646 76186
rect 35646 76134 35656 76186
rect 35680 76134 35710 76186
rect 35710 76134 35722 76186
rect 35722 76134 35736 76186
rect 35760 76134 35774 76186
rect 35774 76134 35786 76186
rect 35786 76134 35816 76186
rect 35840 76134 35850 76186
rect 35850 76134 35896 76186
rect 35600 76132 35656 76134
rect 35680 76132 35736 76134
rect 35760 76132 35816 76134
rect 35840 76132 35896 76134
rect 34940 75642 34996 75644
rect 35020 75642 35076 75644
rect 35100 75642 35156 75644
rect 35180 75642 35236 75644
rect 34940 75590 34986 75642
rect 34986 75590 34996 75642
rect 35020 75590 35050 75642
rect 35050 75590 35062 75642
rect 35062 75590 35076 75642
rect 35100 75590 35114 75642
rect 35114 75590 35126 75642
rect 35126 75590 35156 75642
rect 35180 75590 35190 75642
rect 35190 75590 35236 75642
rect 34940 75588 34996 75590
rect 35020 75588 35076 75590
rect 35100 75588 35156 75590
rect 35180 75588 35236 75590
rect 35600 75098 35656 75100
rect 35680 75098 35736 75100
rect 35760 75098 35816 75100
rect 35840 75098 35896 75100
rect 35600 75046 35646 75098
rect 35646 75046 35656 75098
rect 35680 75046 35710 75098
rect 35710 75046 35722 75098
rect 35722 75046 35736 75098
rect 35760 75046 35774 75098
rect 35774 75046 35786 75098
rect 35786 75046 35816 75098
rect 35840 75046 35850 75098
rect 35850 75046 35896 75098
rect 35600 75044 35656 75046
rect 35680 75044 35736 75046
rect 35760 75044 35816 75046
rect 35840 75044 35896 75046
rect 34940 74554 34996 74556
rect 35020 74554 35076 74556
rect 35100 74554 35156 74556
rect 35180 74554 35236 74556
rect 34940 74502 34986 74554
rect 34986 74502 34996 74554
rect 35020 74502 35050 74554
rect 35050 74502 35062 74554
rect 35062 74502 35076 74554
rect 35100 74502 35114 74554
rect 35114 74502 35126 74554
rect 35126 74502 35156 74554
rect 35180 74502 35190 74554
rect 35190 74502 35236 74554
rect 34940 74500 34996 74502
rect 35020 74500 35076 74502
rect 35100 74500 35156 74502
rect 35180 74500 35236 74502
rect 35600 74010 35656 74012
rect 35680 74010 35736 74012
rect 35760 74010 35816 74012
rect 35840 74010 35896 74012
rect 35600 73958 35646 74010
rect 35646 73958 35656 74010
rect 35680 73958 35710 74010
rect 35710 73958 35722 74010
rect 35722 73958 35736 74010
rect 35760 73958 35774 74010
rect 35774 73958 35786 74010
rect 35786 73958 35816 74010
rect 35840 73958 35850 74010
rect 35850 73958 35896 74010
rect 35600 73956 35656 73958
rect 35680 73956 35736 73958
rect 35760 73956 35816 73958
rect 35840 73956 35896 73958
rect 34940 73466 34996 73468
rect 35020 73466 35076 73468
rect 35100 73466 35156 73468
rect 35180 73466 35236 73468
rect 34940 73414 34986 73466
rect 34986 73414 34996 73466
rect 35020 73414 35050 73466
rect 35050 73414 35062 73466
rect 35062 73414 35076 73466
rect 35100 73414 35114 73466
rect 35114 73414 35126 73466
rect 35126 73414 35156 73466
rect 35180 73414 35190 73466
rect 35190 73414 35236 73466
rect 34940 73412 34996 73414
rect 35020 73412 35076 73414
rect 35100 73412 35156 73414
rect 35180 73412 35236 73414
rect 35600 72922 35656 72924
rect 35680 72922 35736 72924
rect 35760 72922 35816 72924
rect 35840 72922 35896 72924
rect 35600 72870 35646 72922
rect 35646 72870 35656 72922
rect 35680 72870 35710 72922
rect 35710 72870 35722 72922
rect 35722 72870 35736 72922
rect 35760 72870 35774 72922
rect 35774 72870 35786 72922
rect 35786 72870 35816 72922
rect 35840 72870 35850 72922
rect 35850 72870 35896 72922
rect 35600 72868 35656 72870
rect 35680 72868 35736 72870
rect 35760 72868 35816 72870
rect 35840 72868 35896 72870
rect 34940 72378 34996 72380
rect 35020 72378 35076 72380
rect 35100 72378 35156 72380
rect 35180 72378 35236 72380
rect 34940 72326 34986 72378
rect 34986 72326 34996 72378
rect 35020 72326 35050 72378
rect 35050 72326 35062 72378
rect 35062 72326 35076 72378
rect 35100 72326 35114 72378
rect 35114 72326 35126 72378
rect 35126 72326 35156 72378
rect 35180 72326 35190 72378
rect 35190 72326 35236 72378
rect 34940 72324 34996 72326
rect 35020 72324 35076 72326
rect 35100 72324 35156 72326
rect 35180 72324 35236 72326
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 4880 59866 4936 59868
rect 4960 59866 5016 59868
rect 5040 59866 5096 59868
rect 5120 59866 5176 59868
rect 4880 59814 4926 59866
rect 4926 59814 4936 59866
rect 4960 59814 4990 59866
rect 4990 59814 5002 59866
rect 5002 59814 5016 59866
rect 5040 59814 5054 59866
rect 5054 59814 5066 59866
rect 5066 59814 5096 59866
rect 5120 59814 5130 59866
rect 5130 59814 5176 59866
rect 4880 59812 4936 59814
rect 4960 59812 5016 59814
rect 5040 59812 5096 59814
rect 5120 59812 5176 59814
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4880 58778 4936 58780
rect 4960 58778 5016 58780
rect 5040 58778 5096 58780
rect 5120 58778 5176 58780
rect 4880 58726 4926 58778
rect 4926 58726 4936 58778
rect 4960 58726 4990 58778
rect 4990 58726 5002 58778
rect 5002 58726 5016 58778
rect 5040 58726 5054 58778
rect 5054 58726 5066 58778
rect 5066 58726 5096 58778
rect 5120 58726 5130 58778
rect 5130 58726 5176 58778
rect 4880 58724 4936 58726
rect 4960 58724 5016 58726
rect 5040 58724 5096 58726
rect 5120 58724 5176 58726
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4880 57690 4936 57692
rect 4960 57690 5016 57692
rect 5040 57690 5096 57692
rect 5120 57690 5176 57692
rect 4880 57638 4926 57690
rect 4926 57638 4936 57690
rect 4960 57638 4990 57690
rect 4990 57638 5002 57690
rect 5002 57638 5016 57690
rect 5040 57638 5054 57690
rect 5054 57638 5066 57690
rect 5066 57638 5096 57690
rect 5120 57638 5130 57690
rect 5130 57638 5176 57690
rect 4880 57636 4936 57638
rect 4960 57636 5016 57638
rect 5040 57636 5096 57638
rect 5120 57636 5176 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4880 56602 4936 56604
rect 4960 56602 5016 56604
rect 5040 56602 5096 56604
rect 5120 56602 5176 56604
rect 4880 56550 4926 56602
rect 4926 56550 4936 56602
rect 4960 56550 4990 56602
rect 4990 56550 5002 56602
rect 5002 56550 5016 56602
rect 5040 56550 5054 56602
rect 5054 56550 5066 56602
rect 5066 56550 5096 56602
rect 5120 56550 5130 56602
rect 5130 56550 5176 56602
rect 4880 56548 4936 56550
rect 4960 56548 5016 56550
rect 5040 56548 5096 56550
rect 5120 56548 5176 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4880 55514 4936 55516
rect 4960 55514 5016 55516
rect 5040 55514 5096 55516
rect 5120 55514 5176 55516
rect 4880 55462 4926 55514
rect 4926 55462 4936 55514
rect 4960 55462 4990 55514
rect 4990 55462 5002 55514
rect 5002 55462 5016 55514
rect 5040 55462 5054 55514
rect 5054 55462 5066 55514
rect 5066 55462 5096 55514
rect 5120 55462 5130 55514
rect 5130 55462 5176 55514
rect 4880 55460 4936 55462
rect 4960 55460 5016 55462
rect 5040 55460 5096 55462
rect 5120 55460 5176 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4880 54426 4936 54428
rect 4960 54426 5016 54428
rect 5040 54426 5096 54428
rect 5120 54426 5176 54428
rect 4880 54374 4926 54426
rect 4926 54374 4936 54426
rect 4960 54374 4990 54426
rect 4990 54374 5002 54426
rect 5002 54374 5016 54426
rect 5040 54374 5054 54426
rect 5054 54374 5066 54426
rect 5066 54374 5096 54426
rect 5120 54374 5130 54426
rect 5130 54374 5176 54426
rect 4880 54372 4936 54374
rect 4960 54372 5016 54374
rect 5040 54372 5096 54374
rect 5120 54372 5176 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4880 53338 4936 53340
rect 4960 53338 5016 53340
rect 5040 53338 5096 53340
rect 5120 53338 5176 53340
rect 4880 53286 4926 53338
rect 4926 53286 4936 53338
rect 4960 53286 4990 53338
rect 4990 53286 5002 53338
rect 5002 53286 5016 53338
rect 5040 53286 5054 53338
rect 5054 53286 5066 53338
rect 5066 53286 5096 53338
rect 5120 53286 5130 53338
rect 5130 53286 5176 53338
rect 4880 53284 4936 53286
rect 4960 53284 5016 53286
rect 5040 53284 5096 53286
rect 5120 53284 5176 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4880 52250 4936 52252
rect 4960 52250 5016 52252
rect 5040 52250 5096 52252
rect 5120 52250 5176 52252
rect 4880 52198 4926 52250
rect 4926 52198 4936 52250
rect 4960 52198 4990 52250
rect 4990 52198 5002 52250
rect 5002 52198 5016 52250
rect 5040 52198 5054 52250
rect 5054 52198 5066 52250
rect 5066 52198 5096 52250
rect 5120 52198 5130 52250
rect 5130 52198 5176 52250
rect 4880 52196 4936 52198
rect 4960 52196 5016 52198
rect 5040 52196 5096 52198
rect 5120 52196 5176 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4880 51162 4936 51164
rect 4960 51162 5016 51164
rect 5040 51162 5096 51164
rect 5120 51162 5176 51164
rect 4880 51110 4926 51162
rect 4926 51110 4936 51162
rect 4960 51110 4990 51162
rect 4990 51110 5002 51162
rect 5002 51110 5016 51162
rect 5040 51110 5054 51162
rect 5054 51110 5066 51162
rect 5066 51110 5096 51162
rect 5120 51110 5130 51162
rect 5130 51110 5176 51162
rect 4880 51108 4936 51110
rect 4960 51108 5016 51110
rect 5040 51108 5096 51110
rect 5120 51108 5176 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4880 50074 4936 50076
rect 4960 50074 5016 50076
rect 5040 50074 5096 50076
rect 5120 50074 5176 50076
rect 4880 50022 4926 50074
rect 4926 50022 4936 50074
rect 4960 50022 4990 50074
rect 4990 50022 5002 50074
rect 5002 50022 5016 50074
rect 5040 50022 5054 50074
rect 5054 50022 5066 50074
rect 5066 50022 5096 50074
rect 5120 50022 5130 50074
rect 5130 50022 5176 50074
rect 4880 50020 4936 50022
rect 4960 50020 5016 50022
rect 5040 50020 5096 50022
rect 5120 50020 5176 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4880 48986 4936 48988
rect 4960 48986 5016 48988
rect 5040 48986 5096 48988
rect 5120 48986 5176 48988
rect 4880 48934 4926 48986
rect 4926 48934 4936 48986
rect 4960 48934 4990 48986
rect 4990 48934 5002 48986
rect 5002 48934 5016 48986
rect 5040 48934 5054 48986
rect 5054 48934 5066 48986
rect 5066 48934 5096 48986
rect 5120 48934 5130 48986
rect 5130 48934 5176 48986
rect 4880 48932 4936 48934
rect 4960 48932 5016 48934
rect 5040 48932 5096 48934
rect 5120 48932 5176 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4880 47898 4936 47900
rect 4960 47898 5016 47900
rect 5040 47898 5096 47900
rect 5120 47898 5176 47900
rect 4880 47846 4926 47898
rect 4926 47846 4936 47898
rect 4960 47846 4990 47898
rect 4990 47846 5002 47898
rect 5002 47846 5016 47898
rect 5040 47846 5054 47898
rect 5054 47846 5066 47898
rect 5066 47846 5096 47898
rect 5120 47846 5130 47898
rect 5130 47846 5176 47898
rect 4880 47844 4936 47846
rect 4960 47844 5016 47846
rect 5040 47844 5096 47846
rect 5120 47844 5176 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 1490 13640 1546 13696
rect 1306 12960 1362 13016
rect 1490 12280 1546 12336
rect 1214 11600 1270 11656
rect 1490 10920 1546 10976
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1306 10240 1362 10296
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 1490 9560 1546 9616
rect 7562 41248 7618 41304
rect 7286 39480 7342 39536
rect 7562 38392 7618 38448
rect 7562 36644 7618 36680
rect 7562 36624 7564 36644
rect 7564 36624 7616 36644
rect 7616 36624 7618 36644
rect 7470 35536 7526 35592
rect 7562 33924 7618 33960
rect 7562 33904 7564 33924
rect 7564 33904 7616 33924
rect 7616 33904 7618 33924
rect 7470 15408 7526 15464
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 1306 8900 1362 8936
rect 1306 8880 1308 8900
rect 1308 8880 1360 8900
rect 1360 8880 1362 8900
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 1950 8200 2006 8256
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 1306 7520 1362 7576
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1306 6840 1362 6896
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 1214 6160 1270 6216
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 35600 71834 35656 71836
rect 35680 71834 35736 71836
rect 35760 71834 35816 71836
rect 35840 71834 35896 71836
rect 35600 71782 35646 71834
rect 35646 71782 35656 71834
rect 35680 71782 35710 71834
rect 35710 71782 35722 71834
rect 35722 71782 35736 71834
rect 35760 71782 35774 71834
rect 35774 71782 35786 71834
rect 35786 71782 35816 71834
rect 35840 71782 35850 71834
rect 35850 71782 35896 71834
rect 35600 71780 35656 71782
rect 35680 71780 35736 71782
rect 35760 71780 35816 71782
rect 35840 71780 35896 71782
rect 34940 71290 34996 71292
rect 35020 71290 35076 71292
rect 35100 71290 35156 71292
rect 35180 71290 35236 71292
rect 34940 71238 34986 71290
rect 34986 71238 34996 71290
rect 35020 71238 35050 71290
rect 35050 71238 35062 71290
rect 35062 71238 35076 71290
rect 35100 71238 35114 71290
rect 35114 71238 35126 71290
rect 35126 71238 35156 71290
rect 35180 71238 35190 71290
rect 35190 71238 35236 71290
rect 34940 71236 34996 71238
rect 35020 71236 35076 71238
rect 35100 71236 35156 71238
rect 35180 71236 35236 71238
rect 35600 70746 35656 70748
rect 35680 70746 35736 70748
rect 35760 70746 35816 70748
rect 35840 70746 35896 70748
rect 35600 70694 35646 70746
rect 35646 70694 35656 70746
rect 35680 70694 35710 70746
rect 35710 70694 35722 70746
rect 35722 70694 35736 70746
rect 35760 70694 35774 70746
rect 35774 70694 35786 70746
rect 35786 70694 35816 70746
rect 35840 70694 35850 70746
rect 35850 70694 35896 70746
rect 35600 70692 35656 70694
rect 35680 70692 35736 70694
rect 35760 70692 35816 70694
rect 35840 70692 35896 70694
rect 34940 70202 34996 70204
rect 35020 70202 35076 70204
rect 35100 70202 35156 70204
rect 35180 70202 35236 70204
rect 34940 70150 34986 70202
rect 34986 70150 34996 70202
rect 35020 70150 35050 70202
rect 35050 70150 35062 70202
rect 35062 70150 35076 70202
rect 35100 70150 35114 70202
rect 35114 70150 35126 70202
rect 35126 70150 35156 70202
rect 35180 70150 35190 70202
rect 35190 70150 35236 70202
rect 34940 70148 34996 70150
rect 35020 70148 35076 70150
rect 35100 70148 35156 70150
rect 35180 70148 35236 70150
rect 35600 69658 35656 69660
rect 35680 69658 35736 69660
rect 35760 69658 35816 69660
rect 35840 69658 35896 69660
rect 35600 69606 35646 69658
rect 35646 69606 35656 69658
rect 35680 69606 35710 69658
rect 35710 69606 35722 69658
rect 35722 69606 35736 69658
rect 35760 69606 35774 69658
rect 35774 69606 35786 69658
rect 35786 69606 35816 69658
rect 35840 69606 35850 69658
rect 35850 69606 35896 69658
rect 35600 69604 35656 69606
rect 35680 69604 35736 69606
rect 35760 69604 35816 69606
rect 35840 69604 35896 69606
rect 34940 69114 34996 69116
rect 35020 69114 35076 69116
rect 35100 69114 35156 69116
rect 35180 69114 35236 69116
rect 34940 69062 34986 69114
rect 34986 69062 34996 69114
rect 35020 69062 35050 69114
rect 35050 69062 35062 69114
rect 35062 69062 35076 69114
rect 35100 69062 35114 69114
rect 35114 69062 35126 69114
rect 35126 69062 35156 69114
rect 35180 69062 35190 69114
rect 35190 69062 35236 69114
rect 34940 69060 34996 69062
rect 35020 69060 35076 69062
rect 35100 69060 35156 69062
rect 35180 69060 35236 69062
rect 35600 68570 35656 68572
rect 35680 68570 35736 68572
rect 35760 68570 35816 68572
rect 35840 68570 35896 68572
rect 35600 68518 35646 68570
rect 35646 68518 35656 68570
rect 35680 68518 35710 68570
rect 35710 68518 35722 68570
rect 35722 68518 35736 68570
rect 35760 68518 35774 68570
rect 35774 68518 35786 68570
rect 35786 68518 35816 68570
rect 35840 68518 35850 68570
rect 35850 68518 35896 68570
rect 35600 68516 35656 68518
rect 35680 68516 35736 68518
rect 35760 68516 35816 68518
rect 35840 68516 35896 68518
rect 34940 68026 34996 68028
rect 35020 68026 35076 68028
rect 35100 68026 35156 68028
rect 35180 68026 35236 68028
rect 34940 67974 34986 68026
rect 34986 67974 34996 68026
rect 35020 67974 35050 68026
rect 35050 67974 35062 68026
rect 35062 67974 35076 68026
rect 35100 67974 35114 68026
rect 35114 67974 35126 68026
rect 35126 67974 35156 68026
rect 35180 67974 35190 68026
rect 35190 67974 35236 68026
rect 34940 67972 34996 67974
rect 35020 67972 35076 67974
rect 35100 67972 35156 67974
rect 35180 67972 35236 67974
rect 35600 67482 35656 67484
rect 35680 67482 35736 67484
rect 35760 67482 35816 67484
rect 35840 67482 35896 67484
rect 35600 67430 35646 67482
rect 35646 67430 35656 67482
rect 35680 67430 35710 67482
rect 35710 67430 35722 67482
rect 35722 67430 35736 67482
rect 35760 67430 35774 67482
rect 35774 67430 35786 67482
rect 35786 67430 35816 67482
rect 35840 67430 35850 67482
rect 35850 67430 35896 67482
rect 35600 67428 35656 67430
rect 35680 67428 35736 67430
rect 35760 67428 35816 67430
rect 35840 67428 35896 67430
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 35600 66394 35656 66396
rect 35680 66394 35736 66396
rect 35760 66394 35816 66396
rect 35840 66394 35896 66396
rect 35600 66342 35646 66394
rect 35646 66342 35656 66394
rect 35680 66342 35710 66394
rect 35710 66342 35722 66394
rect 35722 66342 35736 66394
rect 35760 66342 35774 66394
rect 35774 66342 35786 66394
rect 35786 66342 35816 66394
rect 35840 66342 35850 66394
rect 35850 66342 35896 66394
rect 35600 66340 35656 66342
rect 35680 66340 35736 66342
rect 35760 66340 35816 66342
rect 35840 66340 35896 66342
rect 37002 79600 37058 79656
rect 37738 78104 37794 78160
rect 40130 77968 40186 78024
rect 40866 77968 40922 78024
rect 40038 77460 40040 77480
rect 40040 77460 40092 77480
rect 40092 77460 40094 77480
rect 40038 77424 40094 77460
rect 37922 77288 37978 77344
rect 39946 77288 40002 77344
rect 42154 79464 42210 79520
rect 43258 79464 43314 79520
rect 42890 77560 42946 77616
rect 43626 77424 43682 77480
rect 42430 77324 42432 77344
rect 42432 77324 42484 77344
rect 42484 77324 42486 77344
rect 42430 77288 42486 77324
rect 63314 78512 63370 78568
rect 65660 77818 65716 77820
rect 65740 77818 65796 77820
rect 65820 77818 65876 77820
rect 65900 77818 65956 77820
rect 65660 77766 65706 77818
rect 65706 77766 65716 77818
rect 65740 77766 65770 77818
rect 65770 77766 65782 77818
rect 65782 77766 65796 77818
rect 65820 77766 65834 77818
rect 65834 77766 65846 77818
rect 65846 77766 65876 77818
rect 65900 77766 65910 77818
rect 65910 77766 65956 77818
rect 65660 77764 65716 77766
rect 65740 77764 65796 77766
rect 65820 77764 65876 77766
rect 65900 77764 65956 77766
rect 65890 77460 65892 77480
rect 65892 77460 65944 77480
rect 65944 77460 65946 77480
rect 65890 77424 65946 77460
rect 65660 76730 65716 76732
rect 65740 76730 65796 76732
rect 65820 76730 65876 76732
rect 65900 76730 65956 76732
rect 65660 76678 65706 76730
rect 65706 76678 65716 76730
rect 65740 76678 65770 76730
rect 65770 76678 65782 76730
rect 65782 76678 65796 76730
rect 65820 76678 65834 76730
rect 65834 76678 65846 76730
rect 65846 76678 65876 76730
rect 65900 76678 65910 76730
rect 65910 76678 65956 76730
rect 65660 76676 65716 76678
rect 65740 76676 65796 76678
rect 65820 76676 65876 76678
rect 65900 76676 65956 76678
rect 65660 75642 65716 75644
rect 65740 75642 65796 75644
rect 65820 75642 65876 75644
rect 65900 75642 65956 75644
rect 65660 75590 65706 75642
rect 65706 75590 65716 75642
rect 65740 75590 65770 75642
rect 65770 75590 65782 75642
rect 65782 75590 65796 75642
rect 65820 75590 65834 75642
rect 65834 75590 65846 75642
rect 65846 75590 65876 75642
rect 65900 75590 65910 75642
rect 65910 75590 65956 75642
rect 65660 75588 65716 75590
rect 65740 75588 65796 75590
rect 65820 75588 65876 75590
rect 65900 75588 65956 75590
rect 65660 74554 65716 74556
rect 65740 74554 65796 74556
rect 65820 74554 65876 74556
rect 65900 74554 65956 74556
rect 65660 74502 65706 74554
rect 65706 74502 65716 74554
rect 65740 74502 65770 74554
rect 65770 74502 65782 74554
rect 65782 74502 65796 74554
rect 65820 74502 65834 74554
rect 65834 74502 65846 74554
rect 65846 74502 65876 74554
rect 65900 74502 65910 74554
rect 65910 74502 65956 74554
rect 65660 74500 65716 74502
rect 65740 74500 65796 74502
rect 65820 74500 65876 74502
rect 65900 74500 65956 74502
rect 65660 73466 65716 73468
rect 65740 73466 65796 73468
rect 65820 73466 65876 73468
rect 65900 73466 65956 73468
rect 65660 73414 65706 73466
rect 65706 73414 65716 73466
rect 65740 73414 65770 73466
rect 65770 73414 65782 73466
rect 65782 73414 65796 73466
rect 65820 73414 65834 73466
rect 65834 73414 65846 73466
rect 65846 73414 65876 73466
rect 65900 73414 65910 73466
rect 65910 73414 65956 73466
rect 65660 73412 65716 73414
rect 65740 73412 65796 73414
rect 65820 73412 65876 73414
rect 65900 73412 65956 73414
rect 65660 72378 65716 72380
rect 65740 72378 65796 72380
rect 65820 72378 65876 72380
rect 65900 72378 65956 72380
rect 65660 72326 65706 72378
rect 65706 72326 65716 72378
rect 65740 72326 65770 72378
rect 65770 72326 65782 72378
rect 65782 72326 65796 72378
rect 65820 72326 65834 72378
rect 65834 72326 65846 72378
rect 65846 72326 65876 72378
rect 65900 72326 65910 72378
rect 65910 72326 65956 72378
rect 65660 72324 65716 72326
rect 65740 72324 65796 72326
rect 65820 72324 65876 72326
rect 65900 72324 65956 72326
rect 65660 71290 65716 71292
rect 65740 71290 65796 71292
rect 65820 71290 65876 71292
rect 65900 71290 65956 71292
rect 65660 71238 65706 71290
rect 65706 71238 65716 71290
rect 65740 71238 65770 71290
rect 65770 71238 65782 71290
rect 65782 71238 65796 71290
rect 65820 71238 65834 71290
rect 65834 71238 65846 71290
rect 65846 71238 65876 71290
rect 65900 71238 65910 71290
rect 65910 71238 65956 71290
rect 65660 71236 65716 71238
rect 65740 71236 65796 71238
rect 65820 71236 65876 71238
rect 65900 71236 65956 71238
rect 65660 70202 65716 70204
rect 65740 70202 65796 70204
rect 65820 70202 65876 70204
rect 65900 70202 65956 70204
rect 65660 70150 65706 70202
rect 65706 70150 65716 70202
rect 65740 70150 65770 70202
rect 65770 70150 65782 70202
rect 65782 70150 65796 70202
rect 65820 70150 65834 70202
rect 65834 70150 65846 70202
rect 65846 70150 65876 70202
rect 65900 70150 65910 70202
rect 65910 70150 65956 70202
rect 65660 70148 65716 70150
rect 65740 70148 65796 70150
rect 65820 70148 65876 70150
rect 65900 70148 65956 70150
rect 65660 69114 65716 69116
rect 65740 69114 65796 69116
rect 65820 69114 65876 69116
rect 65900 69114 65956 69116
rect 65660 69062 65706 69114
rect 65706 69062 65716 69114
rect 65740 69062 65770 69114
rect 65770 69062 65782 69114
rect 65782 69062 65796 69114
rect 65820 69062 65834 69114
rect 65834 69062 65846 69114
rect 65846 69062 65876 69114
rect 65900 69062 65910 69114
rect 65910 69062 65956 69114
rect 65660 69060 65716 69062
rect 65740 69060 65796 69062
rect 65820 69060 65876 69062
rect 65900 69060 65956 69062
rect 65660 68026 65716 68028
rect 65740 68026 65796 68028
rect 65820 68026 65876 68028
rect 65900 68026 65956 68028
rect 65660 67974 65706 68026
rect 65706 67974 65716 68026
rect 65740 67974 65770 68026
rect 65770 67974 65782 68026
rect 65782 67974 65796 68026
rect 65820 67974 65834 68026
rect 65834 67974 65846 68026
rect 65846 67974 65876 68026
rect 65900 67974 65910 68026
rect 65910 67974 65956 68026
rect 65660 67972 65716 67974
rect 65740 67972 65796 67974
rect 65820 67972 65876 67974
rect 65900 67972 65956 67974
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 68466 77580 68522 77616
rect 70950 77968 71006 78024
rect 68466 77560 68468 77580
rect 68468 77560 68520 77580
rect 68520 77560 68522 77580
rect 66320 77274 66376 77276
rect 66400 77274 66456 77276
rect 66480 77274 66536 77276
rect 66560 77274 66616 77276
rect 66320 77222 66366 77274
rect 66366 77222 66376 77274
rect 66400 77222 66430 77274
rect 66430 77222 66442 77274
rect 66442 77222 66456 77274
rect 66480 77222 66494 77274
rect 66494 77222 66506 77274
rect 66506 77222 66536 77274
rect 66560 77222 66570 77274
rect 66570 77222 66616 77274
rect 66320 77220 66376 77222
rect 66400 77220 66456 77222
rect 66480 77220 66536 77222
rect 66560 77220 66616 77222
rect 66320 76186 66376 76188
rect 66400 76186 66456 76188
rect 66480 76186 66536 76188
rect 66560 76186 66616 76188
rect 66320 76134 66366 76186
rect 66366 76134 66376 76186
rect 66400 76134 66430 76186
rect 66430 76134 66442 76186
rect 66442 76134 66456 76186
rect 66480 76134 66494 76186
rect 66494 76134 66506 76186
rect 66506 76134 66536 76186
rect 66560 76134 66570 76186
rect 66570 76134 66616 76186
rect 66320 76132 66376 76134
rect 66400 76132 66456 76134
rect 66480 76132 66536 76134
rect 66560 76132 66616 76134
rect 66320 75098 66376 75100
rect 66400 75098 66456 75100
rect 66480 75098 66536 75100
rect 66560 75098 66616 75100
rect 66320 75046 66366 75098
rect 66366 75046 66376 75098
rect 66400 75046 66430 75098
rect 66430 75046 66442 75098
rect 66442 75046 66456 75098
rect 66480 75046 66494 75098
rect 66494 75046 66506 75098
rect 66506 75046 66536 75098
rect 66560 75046 66570 75098
rect 66570 75046 66616 75098
rect 66320 75044 66376 75046
rect 66400 75044 66456 75046
rect 66480 75044 66536 75046
rect 66560 75044 66616 75046
rect 66320 74010 66376 74012
rect 66400 74010 66456 74012
rect 66480 74010 66536 74012
rect 66560 74010 66616 74012
rect 66320 73958 66366 74010
rect 66366 73958 66376 74010
rect 66400 73958 66430 74010
rect 66430 73958 66442 74010
rect 66442 73958 66456 74010
rect 66480 73958 66494 74010
rect 66494 73958 66506 74010
rect 66506 73958 66536 74010
rect 66560 73958 66570 74010
rect 66570 73958 66616 74010
rect 66320 73956 66376 73958
rect 66400 73956 66456 73958
rect 66480 73956 66536 73958
rect 66560 73956 66616 73958
rect 66320 72922 66376 72924
rect 66400 72922 66456 72924
rect 66480 72922 66536 72924
rect 66560 72922 66616 72924
rect 66320 72870 66366 72922
rect 66366 72870 66376 72922
rect 66400 72870 66430 72922
rect 66430 72870 66442 72922
rect 66442 72870 66456 72922
rect 66480 72870 66494 72922
rect 66494 72870 66506 72922
rect 66506 72870 66536 72922
rect 66560 72870 66570 72922
rect 66570 72870 66616 72922
rect 66320 72868 66376 72870
rect 66400 72868 66456 72870
rect 66480 72868 66536 72870
rect 66560 72868 66616 72870
rect 66320 71834 66376 71836
rect 66400 71834 66456 71836
rect 66480 71834 66536 71836
rect 66560 71834 66616 71836
rect 66320 71782 66366 71834
rect 66366 71782 66376 71834
rect 66400 71782 66430 71834
rect 66430 71782 66442 71834
rect 66442 71782 66456 71834
rect 66480 71782 66494 71834
rect 66494 71782 66506 71834
rect 66506 71782 66536 71834
rect 66560 71782 66570 71834
rect 66570 71782 66616 71834
rect 66320 71780 66376 71782
rect 66400 71780 66456 71782
rect 66480 71780 66536 71782
rect 66560 71780 66616 71782
rect 66320 70746 66376 70748
rect 66400 70746 66456 70748
rect 66480 70746 66536 70748
rect 66560 70746 66616 70748
rect 66320 70694 66366 70746
rect 66366 70694 66376 70746
rect 66400 70694 66430 70746
rect 66430 70694 66442 70746
rect 66442 70694 66456 70746
rect 66480 70694 66494 70746
rect 66494 70694 66506 70746
rect 66506 70694 66536 70746
rect 66560 70694 66570 70746
rect 66570 70694 66616 70746
rect 66320 70692 66376 70694
rect 66400 70692 66456 70694
rect 66480 70692 66536 70694
rect 66560 70692 66616 70694
rect 66320 69658 66376 69660
rect 66400 69658 66456 69660
rect 66480 69658 66536 69660
rect 66560 69658 66616 69660
rect 66320 69606 66366 69658
rect 66366 69606 66376 69658
rect 66400 69606 66430 69658
rect 66430 69606 66442 69658
rect 66442 69606 66456 69658
rect 66480 69606 66494 69658
rect 66494 69606 66506 69658
rect 66506 69606 66536 69658
rect 66560 69606 66570 69658
rect 66570 69606 66616 69658
rect 66320 69604 66376 69606
rect 66400 69604 66456 69606
rect 66480 69604 66536 69606
rect 66560 69604 66616 69606
rect 66320 68570 66376 68572
rect 66400 68570 66456 68572
rect 66480 68570 66536 68572
rect 66560 68570 66616 68572
rect 66320 68518 66366 68570
rect 66366 68518 66376 68570
rect 66400 68518 66430 68570
rect 66430 68518 66442 68570
rect 66442 68518 66456 68570
rect 66480 68518 66494 68570
rect 66494 68518 66506 68570
rect 66506 68518 66536 68570
rect 66560 68518 66570 68570
rect 66570 68518 66616 68570
rect 66320 68516 66376 68518
rect 66400 68516 66456 68518
rect 66480 68516 66536 68518
rect 66560 68516 66616 68518
rect 66320 67482 66376 67484
rect 66400 67482 66456 67484
rect 66480 67482 66536 67484
rect 66560 67482 66616 67484
rect 66320 67430 66366 67482
rect 66366 67430 66376 67482
rect 66400 67430 66430 67482
rect 66430 67430 66442 67482
rect 66442 67430 66456 67482
rect 66480 67430 66494 67482
rect 66494 67430 66506 67482
rect 66506 67430 66536 67482
rect 66560 67430 66570 67482
rect 66570 67430 66616 67482
rect 66320 67428 66376 67430
rect 66400 67428 66456 67430
rect 66480 67428 66536 67430
rect 66560 67428 66616 67430
rect 66320 66394 66376 66396
rect 66400 66394 66456 66396
rect 66480 66394 66536 66396
rect 66560 66394 66616 66396
rect 66320 66342 66366 66394
rect 66366 66342 66376 66394
rect 66400 66342 66430 66394
rect 66430 66342 66442 66394
rect 66442 66342 66456 66394
rect 66480 66342 66494 66394
rect 66494 66342 66506 66394
rect 66506 66342 66536 66394
rect 66560 66342 66570 66394
rect 66570 66342 66616 66394
rect 66320 66340 66376 66342
rect 66400 66340 66456 66342
rect 66480 66340 66536 66342
rect 66560 66340 66616 66342
rect 71686 77968 71742 78024
rect 76194 78240 76250 78296
rect 73986 78104 74042 78160
rect 78770 78376 78826 78432
rect 36082 66172 36084 66192
rect 36084 66172 36136 66192
rect 36136 66172 36138 66192
rect 36082 66136 36138 66172
rect 38474 66172 38476 66192
rect 38476 66172 38528 66192
rect 38528 66172 38530 66192
rect 38474 66136 38530 66172
rect 41142 66172 41144 66192
rect 41144 66172 41196 66192
rect 41196 66172 41198 66192
rect 41142 66136 41198 66172
rect 43626 66172 43628 66192
rect 43628 66172 43680 66192
rect 43680 66172 43682 66192
rect 43626 66136 43682 66172
rect 46110 66172 46112 66192
rect 46112 66172 46164 66192
rect 46164 66172 46166 66192
rect 46110 66136 46166 66172
rect 48594 66172 48596 66192
rect 48596 66172 48648 66192
rect 48648 66172 48650 66192
rect 48594 66136 48650 66172
rect 51078 66172 51080 66192
rect 51080 66172 51132 66192
rect 51132 66172 51134 66192
rect 51078 66136 51134 66172
rect 53562 66172 53564 66192
rect 53564 66172 53616 66192
rect 53616 66172 53618 66192
rect 53562 66136 53618 66172
rect 56138 66172 56140 66192
rect 56140 66172 56192 66192
rect 56192 66172 56194 66192
rect 56138 66136 56194 66172
rect 58622 66172 58624 66192
rect 58624 66172 58676 66192
rect 58676 66172 58678 66192
rect 58622 66136 58678 66172
rect 61106 66172 61108 66192
rect 61108 66172 61160 66192
rect 61160 66172 61162 66192
rect 61106 66136 61162 66172
rect 63590 66172 63592 66192
rect 63592 66172 63644 66192
rect 63644 66172 63646 66192
rect 63590 66136 63646 66172
rect 66074 66172 66076 66192
rect 66076 66172 66128 66192
rect 66128 66172 66130 66192
rect 66074 66136 66130 66172
rect 68558 66172 68560 66192
rect 68560 66172 68612 66192
rect 68612 66172 68614 66192
rect 68558 66136 68614 66172
rect 71042 66172 71044 66192
rect 71044 66172 71096 66192
rect 71096 66172 71098 66192
rect 71042 66136 71098 66172
rect 73526 66172 73528 66192
rect 73528 66172 73580 66192
rect 73580 66172 73582 66192
rect 73526 66136 73582 66172
rect 90546 77152 90602 77208
rect 87694 68992 87750 69048
rect 86314 66136 86370 66192
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 89442 66292 89498 66328
rect 89442 66272 89444 66292
rect 89444 66272 89496 66292
rect 89496 66272 89498 66292
rect 89350 66136 89406 66192
rect 90914 79464 90970 79520
rect 106664 136026 106720 136028
rect 106744 136026 106800 136028
rect 106824 136026 106880 136028
rect 106904 136026 106960 136028
rect 106664 135974 106710 136026
rect 106710 135974 106720 136026
rect 106744 135974 106774 136026
rect 106774 135974 106786 136026
rect 106786 135974 106800 136026
rect 106824 135974 106838 136026
rect 106838 135974 106850 136026
rect 106850 135974 106880 136026
rect 106904 135974 106914 136026
rect 106914 135974 106960 136026
rect 106664 135972 106720 135974
rect 106744 135972 106800 135974
rect 106824 135972 106880 135974
rect 106904 135972 106960 135974
rect 96526 78548 96528 78568
rect 96528 78548 96580 78568
rect 96580 78548 96582 78568
rect 96526 78512 96582 78548
rect 96380 77818 96436 77820
rect 96460 77818 96516 77820
rect 96540 77818 96596 77820
rect 96620 77818 96676 77820
rect 96380 77766 96426 77818
rect 96426 77766 96436 77818
rect 96460 77766 96490 77818
rect 96490 77766 96502 77818
rect 96502 77766 96516 77818
rect 96540 77766 96554 77818
rect 96554 77766 96566 77818
rect 96566 77766 96596 77818
rect 96620 77766 96630 77818
rect 96630 77766 96676 77818
rect 96380 77764 96436 77766
rect 96460 77764 96516 77766
rect 96540 77764 96596 77766
rect 96620 77764 96676 77766
rect 97040 77274 97096 77276
rect 97120 77274 97176 77276
rect 97200 77274 97256 77276
rect 97280 77274 97336 77276
rect 97040 77222 97086 77274
rect 97086 77222 97096 77274
rect 97120 77222 97150 77274
rect 97150 77222 97162 77274
rect 97162 77222 97176 77274
rect 97200 77222 97214 77274
rect 97214 77222 97226 77274
rect 97226 77222 97256 77274
rect 97280 77222 97290 77274
rect 97290 77222 97336 77274
rect 97040 77220 97096 77222
rect 97120 77220 97176 77222
rect 97200 77220 97256 77222
rect 97280 77220 97336 77222
rect 96380 76730 96436 76732
rect 96460 76730 96516 76732
rect 96540 76730 96596 76732
rect 96620 76730 96676 76732
rect 96380 76678 96426 76730
rect 96426 76678 96436 76730
rect 96460 76678 96490 76730
rect 96490 76678 96502 76730
rect 96502 76678 96516 76730
rect 96540 76678 96554 76730
rect 96554 76678 96566 76730
rect 96566 76678 96596 76730
rect 96620 76678 96630 76730
rect 96630 76678 96676 76730
rect 96380 76676 96436 76678
rect 96460 76676 96516 76678
rect 96540 76676 96596 76678
rect 96620 76676 96676 76678
rect 102506 78240 102562 78296
rect 102690 94968 102746 95024
rect 102322 77560 102378 77616
rect 97040 76186 97096 76188
rect 97120 76186 97176 76188
rect 97200 76186 97256 76188
rect 97280 76186 97336 76188
rect 97040 76134 97086 76186
rect 97086 76134 97096 76186
rect 97120 76134 97150 76186
rect 97150 76134 97162 76186
rect 97162 76134 97176 76186
rect 97200 76134 97214 76186
rect 97214 76134 97226 76186
rect 97226 76134 97256 76186
rect 97280 76134 97290 76186
rect 97290 76134 97336 76186
rect 97040 76132 97096 76134
rect 97120 76132 97176 76134
rect 97200 76132 97256 76134
rect 97280 76132 97336 76134
rect 102874 93336 102930 93392
rect 96380 75642 96436 75644
rect 96460 75642 96516 75644
rect 96540 75642 96596 75644
rect 96620 75642 96676 75644
rect 96380 75590 96426 75642
rect 96426 75590 96436 75642
rect 96460 75590 96490 75642
rect 96490 75590 96502 75642
rect 96502 75590 96516 75642
rect 96540 75590 96554 75642
rect 96554 75590 96566 75642
rect 96566 75590 96596 75642
rect 96620 75590 96630 75642
rect 96630 75590 96676 75642
rect 96380 75588 96436 75590
rect 96460 75588 96516 75590
rect 96540 75588 96596 75590
rect 96620 75588 96676 75590
rect 97040 75098 97096 75100
rect 97120 75098 97176 75100
rect 97200 75098 97256 75100
rect 97280 75098 97336 75100
rect 97040 75046 97086 75098
rect 97086 75046 97096 75098
rect 97120 75046 97150 75098
rect 97150 75046 97162 75098
rect 97162 75046 97176 75098
rect 97200 75046 97214 75098
rect 97214 75046 97226 75098
rect 97226 75046 97256 75098
rect 97280 75046 97290 75098
rect 97290 75046 97336 75098
rect 97040 75044 97096 75046
rect 97120 75044 97176 75046
rect 97200 75044 97256 75046
rect 97280 75044 97336 75046
rect 96380 74554 96436 74556
rect 96460 74554 96516 74556
rect 96540 74554 96596 74556
rect 96620 74554 96676 74556
rect 96380 74502 96426 74554
rect 96426 74502 96436 74554
rect 96460 74502 96490 74554
rect 96490 74502 96502 74554
rect 96502 74502 96516 74554
rect 96540 74502 96554 74554
rect 96554 74502 96566 74554
rect 96566 74502 96596 74554
rect 96620 74502 96630 74554
rect 96630 74502 96676 74554
rect 96380 74500 96436 74502
rect 96460 74500 96516 74502
rect 96540 74500 96596 74502
rect 96620 74500 96676 74502
rect 97040 74010 97096 74012
rect 97120 74010 97176 74012
rect 97200 74010 97256 74012
rect 97280 74010 97336 74012
rect 97040 73958 97086 74010
rect 97086 73958 97096 74010
rect 97120 73958 97150 74010
rect 97150 73958 97162 74010
rect 97162 73958 97176 74010
rect 97200 73958 97214 74010
rect 97214 73958 97226 74010
rect 97226 73958 97256 74010
rect 97280 73958 97290 74010
rect 97290 73958 97336 74010
rect 97040 73956 97096 73958
rect 97120 73956 97176 73958
rect 97200 73956 97256 73958
rect 97280 73956 97336 73958
rect 96380 73466 96436 73468
rect 96460 73466 96516 73468
rect 96540 73466 96596 73468
rect 96620 73466 96676 73468
rect 96380 73414 96426 73466
rect 96426 73414 96436 73466
rect 96460 73414 96490 73466
rect 96490 73414 96502 73466
rect 96502 73414 96516 73466
rect 96540 73414 96554 73466
rect 96554 73414 96566 73466
rect 96566 73414 96596 73466
rect 96620 73414 96630 73466
rect 96630 73414 96676 73466
rect 96380 73412 96436 73414
rect 96460 73412 96516 73414
rect 96540 73412 96596 73414
rect 96620 73412 96676 73414
rect 97040 72922 97096 72924
rect 97120 72922 97176 72924
rect 97200 72922 97256 72924
rect 97280 72922 97336 72924
rect 97040 72870 97086 72922
rect 97086 72870 97096 72922
rect 97120 72870 97150 72922
rect 97150 72870 97162 72922
rect 97162 72870 97176 72922
rect 97200 72870 97214 72922
rect 97214 72870 97226 72922
rect 97226 72870 97256 72922
rect 97280 72870 97290 72922
rect 97290 72870 97336 72922
rect 97040 72868 97096 72870
rect 97120 72868 97176 72870
rect 97200 72868 97256 72870
rect 97280 72868 97336 72870
rect 96380 72378 96436 72380
rect 96460 72378 96516 72380
rect 96540 72378 96596 72380
rect 96620 72378 96676 72380
rect 96380 72326 96426 72378
rect 96426 72326 96436 72378
rect 96460 72326 96490 72378
rect 96490 72326 96502 72378
rect 96502 72326 96516 72378
rect 96540 72326 96554 72378
rect 96554 72326 96566 72378
rect 96566 72326 96596 72378
rect 96620 72326 96630 72378
rect 96630 72326 96676 72378
rect 96380 72324 96436 72326
rect 96460 72324 96516 72326
rect 96540 72324 96596 72326
rect 96620 72324 96676 72326
rect 91006 66292 91062 66328
rect 91006 66272 91008 66292
rect 91008 66272 91060 66292
rect 91060 66272 91062 66292
rect 102966 92248 103022 92304
rect 97040 71834 97096 71836
rect 97120 71834 97176 71836
rect 97200 71834 97256 71836
rect 97280 71834 97336 71836
rect 97040 71782 97086 71834
rect 97086 71782 97096 71834
rect 97120 71782 97150 71834
rect 97150 71782 97162 71834
rect 97162 71782 97176 71834
rect 97200 71782 97214 71834
rect 97214 71782 97226 71834
rect 97226 71782 97256 71834
rect 97280 71782 97290 71834
rect 97290 71782 97336 71834
rect 97040 71780 97096 71782
rect 97120 71780 97176 71782
rect 97200 71780 97256 71782
rect 97280 71780 97336 71782
rect 96380 71290 96436 71292
rect 96460 71290 96516 71292
rect 96540 71290 96596 71292
rect 96620 71290 96676 71292
rect 96380 71238 96426 71290
rect 96426 71238 96436 71290
rect 96460 71238 96490 71290
rect 96490 71238 96502 71290
rect 96502 71238 96516 71290
rect 96540 71238 96554 71290
rect 96554 71238 96566 71290
rect 96566 71238 96596 71290
rect 96620 71238 96630 71290
rect 96630 71238 96676 71290
rect 96380 71236 96436 71238
rect 96460 71236 96516 71238
rect 96540 71236 96596 71238
rect 96620 71236 96676 71238
rect 97040 70746 97096 70748
rect 97120 70746 97176 70748
rect 97200 70746 97256 70748
rect 97280 70746 97336 70748
rect 97040 70694 97086 70746
rect 97086 70694 97096 70746
rect 97120 70694 97150 70746
rect 97150 70694 97162 70746
rect 97162 70694 97176 70746
rect 97200 70694 97214 70746
rect 97214 70694 97226 70746
rect 97226 70694 97256 70746
rect 97280 70694 97290 70746
rect 97290 70694 97336 70746
rect 97040 70692 97096 70694
rect 97120 70692 97176 70694
rect 97200 70692 97256 70694
rect 97280 70692 97336 70694
rect 96380 70202 96436 70204
rect 96460 70202 96516 70204
rect 96540 70202 96596 70204
rect 96620 70202 96676 70204
rect 96380 70150 96426 70202
rect 96426 70150 96436 70202
rect 96460 70150 96490 70202
rect 96490 70150 96502 70202
rect 96502 70150 96516 70202
rect 96540 70150 96554 70202
rect 96554 70150 96566 70202
rect 96566 70150 96596 70202
rect 96620 70150 96630 70202
rect 96630 70150 96676 70202
rect 96380 70148 96436 70150
rect 96460 70148 96516 70150
rect 96540 70148 96596 70150
rect 96620 70148 96676 70150
rect 97040 69658 97096 69660
rect 97120 69658 97176 69660
rect 97200 69658 97256 69660
rect 97280 69658 97336 69660
rect 97040 69606 97086 69658
rect 97086 69606 97096 69658
rect 97120 69606 97150 69658
rect 97150 69606 97162 69658
rect 97162 69606 97176 69658
rect 97200 69606 97214 69658
rect 97214 69606 97226 69658
rect 97226 69606 97256 69658
rect 97280 69606 97290 69658
rect 97290 69606 97336 69658
rect 97040 69604 97096 69606
rect 97120 69604 97176 69606
rect 97200 69604 97256 69606
rect 97280 69604 97336 69606
rect 96380 69114 96436 69116
rect 96460 69114 96516 69116
rect 96540 69114 96596 69116
rect 96620 69114 96676 69116
rect 96380 69062 96426 69114
rect 96426 69062 96436 69114
rect 96460 69062 96490 69114
rect 96490 69062 96502 69114
rect 96502 69062 96516 69114
rect 96540 69062 96554 69114
rect 96554 69062 96566 69114
rect 96566 69062 96596 69114
rect 96620 69062 96630 69114
rect 96630 69062 96676 69114
rect 96380 69060 96436 69062
rect 96460 69060 96516 69062
rect 96540 69060 96596 69062
rect 96620 69060 96676 69062
rect 97040 68570 97096 68572
rect 97120 68570 97176 68572
rect 97200 68570 97256 68572
rect 97280 68570 97336 68572
rect 97040 68518 97086 68570
rect 97086 68518 97096 68570
rect 97120 68518 97150 68570
rect 97150 68518 97162 68570
rect 97162 68518 97176 68570
rect 97200 68518 97214 68570
rect 97214 68518 97226 68570
rect 97226 68518 97256 68570
rect 97280 68518 97290 68570
rect 97290 68518 97336 68570
rect 97040 68516 97096 68518
rect 97120 68516 97176 68518
rect 97200 68516 97256 68518
rect 97280 68516 97336 68518
rect 96380 68026 96436 68028
rect 96460 68026 96516 68028
rect 96540 68026 96596 68028
rect 96620 68026 96676 68028
rect 96380 67974 96426 68026
rect 96426 67974 96436 68026
rect 96460 67974 96490 68026
rect 96490 67974 96502 68026
rect 96502 67974 96516 68026
rect 96540 67974 96554 68026
rect 96554 67974 96566 68026
rect 96566 67974 96596 68026
rect 96620 67974 96630 68026
rect 96630 67974 96676 68026
rect 96380 67972 96436 67974
rect 96460 67972 96516 67974
rect 96540 67972 96596 67974
rect 96620 67972 96676 67974
rect 97040 67482 97096 67484
rect 97120 67482 97176 67484
rect 97200 67482 97256 67484
rect 97280 67482 97336 67484
rect 97040 67430 97086 67482
rect 97086 67430 97096 67482
rect 97120 67430 97150 67482
rect 97150 67430 97162 67482
rect 97162 67430 97176 67482
rect 97200 67430 97214 67482
rect 97214 67430 97226 67482
rect 97226 67430 97256 67482
rect 97280 67430 97290 67482
rect 97290 67430 97336 67482
rect 97040 67428 97096 67430
rect 97120 67428 97176 67430
rect 97200 67428 97256 67430
rect 97280 67428 97336 67430
rect 91926 66156 91982 66192
rect 91926 66136 91928 66156
rect 91928 66136 91980 66156
rect 91980 66136 91982 66156
rect 96380 66938 96436 66940
rect 96460 66938 96516 66940
rect 96540 66938 96596 66940
rect 96620 66938 96676 66940
rect 96380 66886 96426 66938
rect 96426 66886 96436 66938
rect 96460 66886 96490 66938
rect 96490 66886 96502 66938
rect 96502 66886 96516 66938
rect 96540 66886 96554 66938
rect 96554 66886 96566 66938
rect 96566 66886 96596 66938
rect 96620 66886 96630 66938
rect 96630 66886 96676 66938
rect 96380 66884 96436 66886
rect 96460 66884 96516 66886
rect 96540 66884 96596 66886
rect 96620 66884 96676 66886
rect 97040 66394 97096 66396
rect 97120 66394 97176 66396
rect 97200 66394 97256 66396
rect 97280 66394 97336 66396
rect 97040 66342 97086 66394
rect 97086 66342 97096 66394
rect 97120 66342 97150 66394
rect 97150 66342 97162 66394
rect 97162 66342 97176 66394
rect 97200 66342 97214 66394
rect 97214 66342 97226 66394
rect 97226 66342 97256 66394
rect 97280 66342 97290 66394
rect 97290 66342 97336 66394
rect 97040 66340 97096 66342
rect 97120 66340 97176 66342
rect 97200 66340 97256 66342
rect 97280 66340 97336 66342
rect 96380 65850 96436 65852
rect 96460 65850 96516 65852
rect 96540 65850 96596 65852
rect 96620 65850 96676 65852
rect 96380 65798 96426 65850
rect 96426 65798 96436 65850
rect 96460 65798 96490 65850
rect 96490 65798 96502 65850
rect 96502 65798 96516 65850
rect 96540 65798 96554 65850
rect 96554 65798 96566 65850
rect 96566 65798 96596 65850
rect 96620 65798 96630 65850
rect 96630 65798 96676 65850
rect 96380 65796 96436 65798
rect 96460 65796 96516 65798
rect 96540 65796 96596 65798
rect 96620 65796 96676 65798
rect 95882 64096 95938 64152
rect 102046 23332 102102 23388
rect 23478 9696 23534 9752
rect 25778 9696 25834 9752
rect 28170 9696 28226 9752
rect 29550 9696 29606 9752
rect 30470 9696 30526 9752
rect 90546 9696 90602 9752
rect 90914 9696 90970 9752
rect 16026 9580 16082 9616
rect 16026 9560 16028 9580
rect 16028 9560 16080 9580
rect 16080 9560 16082 9580
rect 1398 5480 1454 5536
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 1306 4800 1362 4856
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 24674 9560 24730 9616
rect 26698 8880 26754 8936
rect 31666 8200 31722 8256
rect 32954 8200 33010 8256
rect 34242 8200 34298 8256
rect 35438 8200 35494 8256
rect 36358 8200 36414 8256
rect 37462 8200 37518 8256
rect 38750 8200 38806 8256
rect 41326 8200 41382 8256
rect 42154 8200 42210 8256
rect 43442 8200 43498 8256
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 39946 4528 40002 4584
rect 66320 7642 66376 7644
rect 66400 7642 66456 7644
rect 66480 7642 66536 7644
rect 66560 7642 66616 7644
rect 66320 7590 66366 7642
rect 66366 7590 66376 7642
rect 66400 7590 66430 7642
rect 66430 7590 66442 7642
rect 66442 7590 66456 7642
rect 66480 7590 66494 7642
rect 66494 7590 66506 7642
rect 66506 7590 66536 7642
rect 66560 7590 66570 7642
rect 66570 7590 66616 7642
rect 66320 7588 66376 7590
rect 66400 7588 66456 7590
rect 66480 7588 66536 7590
rect 66560 7588 66616 7590
rect 90730 9560 90786 9616
rect 103702 78104 103758 78160
rect 103610 77968 103666 78024
rect 103886 78376 103942 78432
rect 105928 135482 105984 135484
rect 106008 135482 106064 135484
rect 106088 135482 106144 135484
rect 106168 135482 106224 135484
rect 105928 135430 105974 135482
rect 105974 135430 105984 135482
rect 106008 135430 106038 135482
rect 106038 135430 106050 135482
rect 106050 135430 106064 135482
rect 106088 135430 106102 135482
rect 106102 135430 106114 135482
rect 106114 135430 106144 135482
rect 106168 135430 106178 135482
rect 106178 135430 106224 135482
rect 105928 135428 105984 135430
rect 106008 135428 106064 135430
rect 106088 135428 106144 135430
rect 106168 135428 106224 135430
rect 106664 134938 106720 134940
rect 106744 134938 106800 134940
rect 106824 134938 106880 134940
rect 106904 134938 106960 134940
rect 106664 134886 106710 134938
rect 106710 134886 106720 134938
rect 106744 134886 106774 134938
rect 106774 134886 106786 134938
rect 106786 134886 106800 134938
rect 106824 134886 106838 134938
rect 106838 134886 106850 134938
rect 106850 134886 106880 134938
rect 106904 134886 106914 134938
rect 106914 134886 106960 134938
rect 106664 134884 106720 134886
rect 106744 134884 106800 134886
rect 106824 134884 106880 134886
rect 106904 134884 106960 134886
rect 105928 134394 105984 134396
rect 106008 134394 106064 134396
rect 106088 134394 106144 134396
rect 106168 134394 106224 134396
rect 105928 134342 105974 134394
rect 105974 134342 105984 134394
rect 106008 134342 106038 134394
rect 106038 134342 106050 134394
rect 106050 134342 106064 134394
rect 106088 134342 106102 134394
rect 106102 134342 106114 134394
rect 106114 134342 106144 134394
rect 106168 134342 106178 134394
rect 106178 134342 106224 134394
rect 105928 134340 105984 134342
rect 106008 134340 106064 134342
rect 106088 134340 106144 134342
rect 106168 134340 106224 134342
rect 106664 133850 106720 133852
rect 106744 133850 106800 133852
rect 106824 133850 106880 133852
rect 106904 133850 106960 133852
rect 106664 133798 106710 133850
rect 106710 133798 106720 133850
rect 106744 133798 106774 133850
rect 106774 133798 106786 133850
rect 106786 133798 106800 133850
rect 106824 133798 106838 133850
rect 106838 133798 106850 133850
rect 106850 133798 106880 133850
rect 106904 133798 106914 133850
rect 106914 133798 106960 133850
rect 106664 133796 106720 133798
rect 106744 133796 106800 133798
rect 106824 133796 106880 133798
rect 106904 133796 106960 133798
rect 105928 133306 105984 133308
rect 106008 133306 106064 133308
rect 106088 133306 106144 133308
rect 106168 133306 106224 133308
rect 105928 133254 105974 133306
rect 105974 133254 105984 133306
rect 106008 133254 106038 133306
rect 106038 133254 106050 133306
rect 106050 133254 106064 133306
rect 106088 133254 106102 133306
rect 106102 133254 106114 133306
rect 106114 133254 106144 133306
rect 106168 133254 106178 133306
rect 106178 133254 106224 133306
rect 105928 133252 105984 133254
rect 106008 133252 106064 133254
rect 106088 133252 106144 133254
rect 106168 133252 106224 133254
rect 106664 132762 106720 132764
rect 106744 132762 106800 132764
rect 106824 132762 106880 132764
rect 106904 132762 106960 132764
rect 106664 132710 106710 132762
rect 106710 132710 106720 132762
rect 106744 132710 106774 132762
rect 106774 132710 106786 132762
rect 106786 132710 106800 132762
rect 106824 132710 106838 132762
rect 106838 132710 106850 132762
rect 106850 132710 106880 132762
rect 106904 132710 106914 132762
rect 106914 132710 106960 132762
rect 106664 132708 106720 132710
rect 106744 132708 106800 132710
rect 106824 132708 106880 132710
rect 106904 132708 106960 132710
rect 105928 132218 105984 132220
rect 106008 132218 106064 132220
rect 106088 132218 106144 132220
rect 106168 132218 106224 132220
rect 105928 132166 105974 132218
rect 105974 132166 105984 132218
rect 106008 132166 106038 132218
rect 106038 132166 106050 132218
rect 106050 132166 106064 132218
rect 106088 132166 106102 132218
rect 106102 132166 106114 132218
rect 106114 132166 106144 132218
rect 106168 132166 106178 132218
rect 106178 132166 106224 132218
rect 105928 132164 105984 132166
rect 106008 132164 106064 132166
rect 106088 132164 106144 132166
rect 106168 132164 106224 132166
rect 106664 131674 106720 131676
rect 106744 131674 106800 131676
rect 106824 131674 106880 131676
rect 106904 131674 106960 131676
rect 106664 131622 106710 131674
rect 106710 131622 106720 131674
rect 106744 131622 106774 131674
rect 106774 131622 106786 131674
rect 106786 131622 106800 131674
rect 106824 131622 106838 131674
rect 106838 131622 106850 131674
rect 106850 131622 106880 131674
rect 106904 131622 106914 131674
rect 106914 131622 106960 131674
rect 106664 131620 106720 131622
rect 106744 131620 106800 131622
rect 106824 131620 106880 131622
rect 106904 131620 106960 131622
rect 105928 131130 105984 131132
rect 106008 131130 106064 131132
rect 106088 131130 106144 131132
rect 106168 131130 106224 131132
rect 105928 131078 105974 131130
rect 105974 131078 105984 131130
rect 106008 131078 106038 131130
rect 106038 131078 106050 131130
rect 106050 131078 106064 131130
rect 106088 131078 106102 131130
rect 106102 131078 106114 131130
rect 106114 131078 106144 131130
rect 106168 131078 106178 131130
rect 106178 131078 106224 131130
rect 105928 131076 105984 131078
rect 106008 131076 106064 131078
rect 106088 131076 106144 131078
rect 106168 131076 106224 131078
rect 106664 130586 106720 130588
rect 106744 130586 106800 130588
rect 106824 130586 106880 130588
rect 106904 130586 106960 130588
rect 106664 130534 106710 130586
rect 106710 130534 106720 130586
rect 106744 130534 106774 130586
rect 106774 130534 106786 130586
rect 106786 130534 106800 130586
rect 106824 130534 106838 130586
rect 106838 130534 106850 130586
rect 106850 130534 106880 130586
rect 106904 130534 106914 130586
rect 106914 130534 106960 130586
rect 106664 130532 106720 130534
rect 106744 130532 106800 130534
rect 106824 130532 106880 130534
rect 106904 130532 106960 130534
rect 105928 130042 105984 130044
rect 106008 130042 106064 130044
rect 106088 130042 106144 130044
rect 106168 130042 106224 130044
rect 105928 129990 105974 130042
rect 105974 129990 105984 130042
rect 106008 129990 106038 130042
rect 106038 129990 106050 130042
rect 106050 129990 106064 130042
rect 106088 129990 106102 130042
rect 106102 129990 106114 130042
rect 106114 129990 106144 130042
rect 106168 129990 106178 130042
rect 106178 129990 106224 130042
rect 105928 129988 105984 129990
rect 106008 129988 106064 129990
rect 106088 129988 106144 129990
rect 106168 129988 106224 129990
rect 104346 129820 104348 129840
rect 104348 129820 104400 129840
rect 104400 129820 104402 129840
rect 104346 129784 104402 129820
rect 106664 129498 106720 129500
rect 106744 129498 106800 129500
rect 106824 129498 106880 129500
rect 106904 129498 106960 129500
rect 106664 129446 106710 129498
rect 106710 129446 106720 129498
rect 106744 129446 106774 129498
rect 106774 129446 106786 129498
rect 106786 129446 106800 129498
rect 106824 129446 106838 129498
rect 106838 129446 106850 129498
rect 106850 129446 106880 129498
rect 106904 129446 106914 129498
rect 106914 129446 106960 129498
rect 106664 129444 106720 129446
rect 106744 129444 106800 129446
rect 106824 129444 106880 129446
rect 106904 129444 106960 129446
rect 105928 128954 105984 128956
rect 106008 128954 106064 128956
rect 106088 128954 106144 128956
rect 106168 128954 106224 128956
rect 105928 128902 105974 128954
rect 105974 128902 105984 128954
rect 106008 128902 106038 128954
rect 106038 128902 106050 128954
rect 106050 128902 106064 128954
rect 106088 128902 106102 128954
rect 106102 128902 106114 128954
rect 106114 128902 106144 128954
rect 106168 128902 106178 128954
rect 106178 128902 106224 128954
rect 105928 128900 105984 128902
rect 106008 128900 106064 128902
rect 106088 128900 106144 128902
rect 106168 128900 106224 128902
rect 106664 128410 106720 128412
rect 106744 128410 106800 128412
rect 106824 128410 106880 128412
rect 106904 128410 106960 128412
rect 106664 128358 106710 128410
rect 106710 128358 106720 128410
rect 106744 128358 106774 128410
rect 106774 128358 106786 128410
rect 106786 128358 106800 128410
rect 106824 128358 106838 128410
rect 106838 128358 106850 128410
rect 106850 128358 106880 128410
rect 106904 128358 106914 128410
rect 106914 128358 106960 128410
rect 106664 128356 106720 128358
rect 106744 128356 106800 128358
rect 106824 128356 106880 128358
rect 106904 128356 106960 128358
rect 105928 127866 105984 127868
rect 106008 127866 106064 127868
rect 106088 127866 106144 127868
rect 106168 127866 106224 127868
rect 105928 127814 105974 127866
rect 105974 127814 105984 127866
rect 106008 127814 106038 127866
rect 106038 127814 106050 127866
rect 106050 127814 106064 127866
rect 106088 127814 106102 127866
rect 106102 127814 106114 127866
rect 106114 127814 106144 127866
rect 106168 127814 106178 127866
rect 106178 127814 106224 127866
rect 105928 127812 105984 127814
rect 106008 127812 106064 127814
rect 106088 127812 106144 127814
rect 106168 127812 106224 127814
rect 106664 127322 106720 127324
rect 106744 127322 106800 127324
rect 106824 127322 106880 127324
rect 106904 127322 106960 127324
rect 106664 127270 106710 127322
rect 106710 127270 106720 127322
rect 106744 127270 106774 127322
rect 106774 127270 106786 127322
rect 106786 127270 106800 127322
rect 106824 127270 106838 127322
rect 106838 127270 106850 127322
rect 106850 127270 106880 127322
rect 106904 127270 106914 127322
rect 106914 127270 106960 127322
rect 106664 127268 106720 127270
rect 106744 127268 106800 127270
rect 106824 127268 106880 127270
rect 106904 127268 106960 127270
rect 105928 126778 105984 126780
rect 106008 126778 106064 126780
rect 106088 126778 106144 126780
rect 106168 126778 106224 126780
rect 105928 126726 105974 126778
rect 105974 126726 105984 126778
rect 106008 126726 106038 126778
rect 106038 126726 106050 126778
rect 106050 126726 106064 126778
rect 106088 126726 106102 126778
rect 106102 126726 106114 126778
rect 106114 126726 106144 126778
rect 106168 126726 106178 126778
rect 106178 126726 106224 126778
rect 105928 126724 105984 126726
rect 106008 126724 106064 126726
rect 106088 126724 106144 126726
rect 106168 126724 106224 126726
rect 106664 126234 106720 126236
rect 106744 126234 106800 126236
rect 106824 126234 106880 126236
rect 106904 126234 106960 126236
rect 106664 126182 106710 126234
rect 106710 126182 106720 126234
rect 106744 126182 106774 126234
rect 106774 126182 106786 126234
rect 106786 126182 106800 126234
rect 106824 126182 106838 126234
rect 106838 126182 106850 126234
rect 106850 126182 106880 126234
rect 106904 126182 106914 126234
rect 106914 126182 106960 126234
rect 106664 126180 106720 126182
rect 106744 126180 106800 126182
rect 106824 126180 106880 126182
rect 106904 126180 106960 126182
rect 105928 125690 105984 125692
rect 106008 125690 106064 125692
rect 106088 125690 106144 125692
rect 106168 125690 106224 125692
rect 105928 125638 105974 125690
rect 105974 125638 105984 125690
rect 106008 125638 106038 125690
rect 106038 125638 106050 125690
rect 106050 125638 106064 125690
rect 106088 125638 106102 125690
rect 106102 125638 106114 125690
rect 106114 125638 106144 125690
rect 106168 125638 106178 125690
rect 106178 125638 106224 125690
rect 105928 125636 105984 125638
rect 106008 125636 106064 125638
rect 106088 125636 106144 125638
rect 106168 125636 106224 125638
rect 106664 125146 106720 125148
rect 106744 125146 106800 125148
rect 106824 125146 106880 125148
rect 106904 125146 106960 125148
rect 106664 125094 106710 125146
rect 106710 125094 106720 125146
rect 106744 125094 106774 125146
rect 106774 125094 106786 125146
rect 106786 125094 106800 125146
rect 106824 125094 106838 125146
rect 106838 125094 106850 125146
rect 106850 125094 106880 125146
rect 106904 125094 106914 125146
rect 106914 125094 106960 125146
rect 106664 125092 106720 125094
rect 106744 125092 106800 125094
rect 106824 125092 106880 125094
rect 106904 125092 106960 125094
rect 105928 124602 105984 124604
rect 106008 124602 106064 124604
rect 106088 124602 106144 124604
rect 106168 124602 106224 124604
rect 105928 124550 105974 124602
rect 105974 124550 105984 124602
rect 106008 124550 106038 124602
rect 106038 124550 106050 124602
rect 106050 124550 106064 124602
rect 106088 124550 106102 124602
rect 106102 124550 106114 124602
rect 106114 124550 106144 124602
rect 106168 124550 106178 124602
rect 106178 124550 106224 124602
rect 105928 124548 105984 124550
rect 106008 124548 106064 124550
rect 106088 124548 106144 124550
rect 106168 124548 106224 124550
rect 106664 124058 106720 124060
rect 106744 124058 106800 124060
rect 106824 124058 106880 124060
rect 106904 124058 106960 124060
rect 106664 124006 106710 124058
rect 106710 124006 106720 124058
rect 106744 124006 106774 124058
rect 106774 124006 106786 124058
rect 106786 124006 106800 124058
rect 106824 124006 106838 124058
rect 106838 124006 106850 124058
rect 106850 124006 106880 124058
rect 106904 124006 106914 124058
rect 106914 124006 106960 124058
rect 106664 124004 106720 124006
rect 106744 124004 106800 124006
rect 106824 124004 106880 124006
rect 106904 124004 106960 124006
rect 105928 123514 105984 123516
rect 106008 123514 106064 123516
rect 106088 123514 106144 123516
rect 106168 123514 106224 123516
rect 105928 123462 105974 123514
rect 105974 123462 105984 123514
rect 106008 123462 106038 123514
rect 106038 123462 106050 123514
rect 106050 123462 106064 123514
rect 106088 123462 106102 123514
rect 106102 123462 106114 123514
rect 106114 123462 106144 123514
rect 106168 123462 106178 123514
rect 106178 123462 106224 123514
rect 105928 123460 105984 123462
rect 106008 123460 106064 123462
rect 106088 123460 106144 123462
rect 106168 123460 106224 123462
rect 106664 122970 106720 122972
rect 106744 122970 106800 122972
rect 106824 122970 106880 122972
rect 106904 122970 106960 122972
rect 106664 122918 106710 122970
rect 106710 122918 106720 122970
rect 106744 122918 106774 122970
rect 106774 122918 106786 122970
rect 106786 122918 106800 122970
rect 106824 122918 106838 122970
rect 106838 122918 106850 122970
rect 106850 122918 106880 122970
rect 106904 122918 106914 122970
rect 106914 122918 106960 122970
rect 106664 122916 106720 122918
rect 106744 122916 106800 122918
rect 106824 122916 106880 122918
rect 106904 122916 106960 122918
rect 105928 122426 105984 122428
rect 106008 122426 106064 122428
rect 106088 122426 106144 122428
rect 106168 122426 106224 122428
rect 105928 122374 105974 122426
rect 105974 122374 105984 122426
rect 106008 122374 106038 122426
rect 106038 122374 106050 122426
rect 106050 122374 106064 122426
rect 106088 122374 106102 122426
rect 106102 122374 106114 122426
rect 106114 122374 106144 122426
rect 106168 122374 106178 122426
rect 106178 122374 106224 122426
rect 105928 122372 105984 122374
rect 106008 122372 106064 122374
rect 106088 122372 106144 122374
rect 106168 122372 106224 122374
rect 106664 121882 106720 121884
rect 106744 121882 106800 121884
rect 106824 121882 106880 121884
rect 106904 121882 106960 121884
rect 106664 121830 106710 121882
rect 106710 121830 106720 121882
rect 106744 121830 106774 121882
rect 106774 121830 106786 121882
rect 106786 121830 106800 121882
rect 106824 121830 106838 121882
rect 106838 121830 106850 121882
rect 106850 121830 106880 121882
rect 106904 121830 106914 121882
rect 106914 121830 106960 121882
rect 106664 121828 106720 121830
rect 106744 121828 106800 121830
rect 106824 121828 106880 121830
rect 106904 121828 106960 121830
rect 105928 121338 105984 121340
rect 106008 121338 106064 121340
rect 106088 121338 106144 121340
rect 106168 121338 106224 121340
rect 105928 121286 105974 121338
rect 105974 121286 105984 121338
rect 106008 121286 106038 121338
rect 106038 121286 106050 121338
rect 106050 121286 106064 121338
rect 106088 121286 106102 121338
rect 106102 121286 106114 121338
rect 106114 121286 106144 121338
rect 106168 121286 106178 121338
rect 106178 121286 106224 121338
rect 105928 121284 105984 121286
rect 106008 121284 106064 121286
rect 106088 121284 106144 121286
rect 106168 121284 106224 121286
rect 106664 120794 106720 120796
rect 106744 120794 106800 120796
rect 106824 120794 106880 120796
rect 106904 120794 106960 120796
rect 106664 120742 106710 120794
rect 106710 120742 106720 120794
rect 106744 120742 106774 120794
rect 106774 120742 106786 120794
rect 106786 120742 106800 120794
rect 106824 120742 106838 120794
rect 106838 120742 106850 120794
rect 106850 120742 106880 120794
rect 106904 120742 106914 120794
rect 106914 120742 106960 120794
rect 106664 120740 106720 120742
rect 106744 120740 106800 120742
rect 106824 120740 106880 120742
rect 106904 120740 106960 120742
rect 105928 120250 105984 120252
rect 106008 120250 106064 120252
rect 106088 120250 106144 120252
rect 106168 120250 106224 120252
rect 105928 120198 105974 120250
rect 105974 120198 105984 120250
rect 106008 120198 106038 120250
rect 106038 120198 106050 120250
rect 106050 120198 106064 120250
rect 106088 120198 106102 120250
rect 106102 120198 106114 120250
rect 106114 120198 106144 120250
rect 106168 120198 106178 120250
rect 106178 120198 106224 120250
rect 105928 120196 105984 120198
rect 106008 120196 106064 120198
rect 106088 120196 106144 120198
rect 106168 120196 106224 120198
rect 106664 119706 106720 119708
rect 106744 119706 106800 119708
rect 106824 119706 106880 119708
rect 106904 119706 106960 119708
rect 106664 119654 106710 119706
rect 106710 119654 106720 119706
rect 106744 119654 106774 119706
rect 106774 119654 106786 119706
rect 106786 119654 106800 119706
rect 106824 119654 106838 119706
rect 106838 119654 106850 119706
rect 106850 119654 106880 119706
rect 106904 119654 106914 119706
rect 106914 119654 106960 119706
rect 106664 119652 106720 119654
rect 106744 119652 106800 119654
rect 106824 119652 106880 119654
rect 106904 119652 106960 119654
rect 105928 119162 105984 119164
rect 106008 119162 106064 119164
rect 106088 119162 106144 119164
rect 106168 119162 106224 119164
rect 105928 119110 105974 119162
rect 105974 119110 105984 119162
rect 106008 119110 106038 119162
rect 106038 119110 106050 119162
rect 106050 119110 106064 119162
rect 106088 119110 106102 119162
rect 106102 119110 106114 119162
rect 106114 119110 106144 119162
rect 106168 119110 106178 119162
rect 106178 119110 106224 119162
rect 105928 119108 105984 119110
rect 106008 119108 106064 119110
rect 106088 119108 106144 119110
rect 106168 119108 106224 119110
rect 106664 118618 106720 118620
rect 106744 118618 106800 118620
rect 106824 118618 106880 118620
rect 106904 118618 106960 118620
rect 106664 118566 106710 118618
rect 106710 118566 106720 118618
rect 106744 118566 106774 118618
rect 106774 118566 106786 118618
rect 106786 118566 106800 118618
rect 106824 118566 106838 118618
rect 106838 118566 106850 118618
rect 106850 118566 106880 118618
rect 106904 118566 106914 118618
rect 106914 118566 106960 118618
rect 106664 118564 106720 118566
rect 106744 118564 106800 118566
rect 106824 118564 106880 118566
rect 106904 118564 106960 118566
rect 105928 118074 105984 118076
rect 106008 118074 106064 118076
rect 106088 118074 106144 118076
rect 106168 118074 106224 118076
rect 105928 118022 105974 118074
rect 105974 118022 105984 118074
rect 106008 118022 106038 118074
rect 106038 118022 106050 118074
rect 106050 118022 106064 118074
rect 106088 118022 106102 118074
rect 106102 118022 106114 118074
rect 106114 118022 106144 118074
rect 106168 118022 106178 118074
rect 106178 118022 106224 118074
rect 105928 118020 105984 118022
rect 106008 118020 106064 118022
rect 106088 118020 106144 118022
rect 106168 118020 106224 118022
rect 106664 117530 106720 117532
rect 106744 117530 106800 117532
rect 106824 117530 106880 117532
rect 106904 117530 106960 117532
rect 106664 117478 106710 117530
rect 106710 117478 106720 117530
rect 106744 117478 106774 117530
rect 106774 117478 106786 117530
rect 106786 117478 106800 117530
rect 106824 117478 106838 117530
rect 106838 117478 106850 117530
rect 106850 117478 106880 117530
rect 106904 117478 106914 117530
rect 106914 117478 106960 117530
rect 106664 117476 106720 117478
rect 106744 117476 106800 117478
rect 106824 117476 106880 117478
rect 106904 117476 106960 117478
rect 105928 116986 105984 116988
rect 106008 116986 106064 116988
rect 106088 116986 106144 116988
rect 106168 116986 106224 116988
rect 105928 116934 105974 116986
rect 105974 116934 105984 116986
rect 106008 116934 106038 116986
rect 106038 116934 106050 116986
rect 106050 116934 106064 116986
rect 106088 116934 106102 116986
rect 106102 116934 106114 116986
rect 106114 116934 106144 116986
rect 106168 116934 106178 116986
rect 106178 116934 106224 116986
rect 105928 116932 105984 116934
rect 106008 116932 106064 116934
rect 106088 116932 106144 116934
rect 106168 116932 106224 116934
rect 106664 116442 106720 116444
rect 106744 116442 106800 116444
rect 106824 116442 106880 116444
rect 106904 116442 106960 116444
rect 106664 116390 106710 116442
rect 106710 116390 106720 116442
rect 106744 116390 106774 116442
rect 106774 116390 106786 116442
rect 106786 116390 106800 116442
rect 106824 116390 106838 116442
rect 106838 116390 106850 116442
rect 106850 116390 106880 116442
rect 106904 116390 106914 116442
rect 106914 116390 106960 116442
rect 106664 116388 106720 116390
rect 106744 116388 106800 116390
rect 106824 116388 106880 116390
rect 106904 116388 106960 116390
rect 105928 115898 105984 115900
rect 106008 115898 106064 115900
rect 106088 115898 106144 115900
rect 106168 115898 106224 115900
rect 105928 115846 105974 115898
rect 105974 115846 105984 115898
rect 106008 115846 106038 115898
rect 106038 115846 106050 115898
rect 106050 115846 106064 115898
rect 106088 115846 106102 115898
rect 106102 115846 106114 115898
rect 106114 115846 106144 115898
rect 106168 115846 106178 115898
rect 106178 115846 106224 115898
rect 105928 115844 105984 115846
rect 106008 115844 106064 115846
rect 106088 115844 106144 115846
rect 106168 115844 106224 115846
rect 106664 115354 106720 115356
rect 106744 115354 106800 115356
rect 106824 115354 106880 115356
rect 106904 115354 106960 115356
rect 106664 115302 106710 115354
rect 106710 115302 106720 115354
rect 106744 115302 106774 115354
rect 106774 115302 106786 115354
rect 106786 115302 106800 115354
rect 106824 115302 106838 115354
rect 106838 115302 106850 115354
rect 106850 115302 106880 115354
rect 106904 115302 106914 115354
rect 106914 115302 106960 115354
rect 106664 115300 106720 115302
rect 106744 115300 106800 115302
rect 106824 115300 106880 115302
rect 106904 115300 106960 115302
rect 105928 114810 105984 114812
rect 106008 114810 106064 114812
rect 106088 114810 106144 114812
rect 106168 114810 106224 114812
rect 105928 114758 105974 114810
rect 105974 114758 105984 114810
rect 106008 114758 106038 114810
rect 106038 114758 106050 114810
rect 106050 114758 106064 114810
rect 106088 114758 106102 114810
rect 106102 114758 106114 114810
rect 106114 114758 106144 114810
rect 106168 114758 106178 114810
rect 106178 114758 106224 114810
rect 105928 114756 105984 114758
rect 106008 114756 106064 114758
rect 106088 114756 106144 114758
rect 106168 114756 106224 114758
rect 106664 114266 106720 114268
rect 106744 114266 106800 114268
rect 106824 114266 106880 114268
rect 106904 114266 106960 114268
rect 106664 114214 106710 114266
rect 106710 114214 106720 114266
rect 106744 114214 106774 114266
rect 106774 114214 106786 114266
rect 106786 114214 106800 114266
rect 106824 114214 106838 114266
rect 106838 114214 106850 114266
rect 106850 114214 106880 114266
rect 106904 114214 106914 114266
rect 106914 114214 106960 114266
rect 106664 114212 106720 114214
rect 106744 114212 106800 114214
rect 106824 114212 106880 114214
rect 106904 114212 106960 114214
rect 105928 113722 105984 113724
rect 106008 113722 106064 113724
rect 106088 113722 106144 113724
rect 106168 113722 106224 113724
rect 105928 113670 105974 113722
rect 105974 113670 105984 113722
rect 106008 113670 106038 113722
rect 106038 113670 106050 113722
rect 106050 113670 106064 113722
rect 106088 113670 106102 113722
rect 106102 113670 106114 113722
rect 106114 113670 106144 113722
rect 106168 113670 106178 113722
rect 106178 113670 106224 113722
rect 105928 113668 105984 113670
rect 106008 113668 106064 113670
rect 106088 113668 106144 113670
rect 106168 113668 106224 113670
rect 106664 113178 106720 113180
rect 106744 113178 106800 113180
rect 106824 113178 106880 113180
rect 106904 113178 106960 113180
rect 106664 113126 106710 113178
rect 106710 113126 106720 113178
rect 106744 113126 106774 113178
rect 106774 113126 106786 113178
rect 106786 113126 106800 113178
rect 106824 113126 106838 113178
rect 106838 113126 106850 113178
rect 106850 113126 106880 113178
rect 106904 113126 106914 113178
rect 106914 113126 106960 113178
rect 106664 113124 106720 113126
rect 106744 113124 106800 113126
rect 106824 113124 106880 113126
rect 106904 113124 106960 113126
rect 105928 112634 105984 112636
rect 106008 112634 106064 112636
rect 106088 112634 106144 112636
rect 106168 112634 106224 112636
rect 105928 112582 105974 112634
rect 105974 112582 105984 112634
rect 106008 112582 106038 112634
rect 106038 112582 106050 112634
rect 106050 112582 106064 112634
rect 106088 112582 106102 112634
rect 106102 112582 106114 112634
rect 106114 112582 106144 112634
rect 106168 112582 106178 112634
rect 106178 112582 106224 112634
rect 105928 112580 105984 112582
rect 106008 112580 106064 112582
rect 106088 112580 106144 112582
rect 106168 112580 106224 112582
rect 106664 112090 106720 112092
rect 106744 112090 106800 112092
rect 106824 112090 106880 112092
rect 106904 112090 106960 112092
rect 106664 112038 106710 112090
rect 106710 112038 106720 112090
rect 106744 112038 106774 112090
rect 106774 112038 106786 112090
rect 106786 112038 106800 112090
rect 106824 112038 106838 112090
rect 106838 112038 106850 112090
rect 106850 112038 106880 112090
rect 106904 112038 106914 112090
rect 106914 112038 106960 112090
rect 106664 112036 106720 112038
rect 106744 112036 106800 112038
rect 106824 112036 106880 112038
rect 106904 112036 106960 112038
rect 105928 111546 105984 111548
rect 106008 111546 106064 111548
rect 106088 111546 106144 111548
rect 106168 111546 106224 111548
rect 105928 111494 105974 111546
rect 105974 111494 105984 111546
rect 106008 111494 106038 111546
rect 106038 111494 106050 111546
rect 106050 111494 106064 111546
rect 106088 111494 106102 111546
rect 106102 111494 106114 111546
rect 106114 111494 106144 111546
rect 106168 111494 106178 111546
rect 106178 111494 106224 111546
rect 105928 111492 105984 111494
rect 106008 111492 106064 111494
rect 106088 111492 106144 111494
rect 106168 111492 106224 111494
rect 106664 111002 106720 111004
rect 106744 111002 106800 111004
rect 106824 111002 106880 111004
rect 106904 111002 106960 111004
rect 106664 110950 106710 111002
rect 106710 110950 106720 111002
rect 106744 110950 106774 111002
rect 106774 110950 106786 111002
rect 106786 110950 106800 111002
rect 106824 110950 106838 111002
rect 106838 110950 106850 111002
rect 106850 110950 106880 111002
rect 106904 110950 106914 111002
rect 106914 110950 106960 111002
rect 106664 110948 106720 110950
rect 106744 110948 106800 110950
rect 106824 110948 106880 110950
rect 106904 110948 106960 110950
rect 105928 110458 105984 110460
rect 106008 110458 106064 110460
rect 106088 110458 106144 110460
rect 106168 110458 106224 110460
rect 105928 110406 105974 110458
rect 105974 110406 105984 110458
rect 106008 110406 106038 110458
rect 106038 110406 106050 110458
rect 106050 110406 106064 110458
rect 106088 110406 106102 110458
rect 106102 110406 106114 110458
rect 106114 110406 106144 110458
rect 106168 110406 106178 110458
rect 106178 110406 106224 110458
rect 105928 110404 105984 110406
rect 106008 110404 106064 110406
rect 106088 110404 106144 110406
rect 106168 110404 106224 110406
rect 106664 109914 106720 109916
rect 106744 109914 106800 109916
rect 106824 109914 106880 109916
rect 106904 109914 106960 109916
rect 106664 109862 106710 109914
rect 106710 109862 106720 109914
rect 106744 109862 106774 109914
rect 106774 109862 106786 109914
rect 106786 109862 106800 109914
rect 106824 109862 106838 109914
rect 106838 109862 106850 109914
rect 106850 109862 106880 109914
rect 106904 109862 106914 109914
rect 106914 109862 106960 109914
rect 106664 109860 106720 109862
rect 106744 109860 106800 109862
rect 106824 109860 106880 109862
rect 106904 109860 106960 109862
rect 105928 109370 105984 109372
rect 106008 109370 106064 109372
rect 106088 109370 106144 109372
rect 106168 109370 106224 109372
rect 105928 109318 105974 109370
rect 105974 109318 105984 109370
rect 106008 109318 106038 109370
rect 106038 109318 106050 109370
rect 106050 109318 106064 109370
rect 106088 109318 106102 109370
rect 106102 109318 106114 109370
rect 106114 109318 106144 109370
rect 106168 109318 106178 109370
rect 106178 109318 106224 109370
rect 105928 109316 105984 109318
rect 106008 109316 106064 109318
rect 106088 109316 106144 109318
rect 106168 109316 106224 109318
rect 106664 108826 106720 108828
rect 106744 108826 106800 108828
rect 106824 108826 106880 108828
rect 106904 108826 106960 108828
rect 106664 108774 106710 108826
rect 106710 108774 106720 108826
rect 106744 108774 106774 108826
rect 106774 108774 106786 108826
rect 106786 108774 106800 108826
rect 106824 108774 106838 108826
rect 106838 108774 106850 108826
rect 106850 108774 106880 108826
rect 106904 108774 106914 108826
rect 106914 108774 106960 108826
rect 106664 108772 106720 108774
rect 106744 108772 106800 108774
rect 106824 108772 106880 108774
rect 106904 108772 106960 108774
rect 105928 108282 105984 108284
rect 106008 108282 106064 108284
rect 106088 108282 106144 108284
rect 106168 108282 106224 108284
rect 105928 108230 105974 108282
rect 105974 108230 105984 108282
rect 106008 108230 106038 108282
rect 106038 108230 106050 108282
rect 106050 108230 106064 108282
rect 106088 108230 106102 108282
rect 106102 108230 106114 108282
rect 106114 108230 106144 108282
rect 106168 108230 106178 108282
rect 106178 108230 106224 108282
rect 105928 108228 105984 108230
rect 106008 108228 106064 108230
rect 106088 108228 106144 108230
rect 106168 108228 106224 108230
rect 106664 107738 106720 107740
rect 106744 107738 106800 107740
rect 106824 107738 106880 107740
rect 106904 107738 106960 107740
rect 106664 107686 106710 107738
rect 106710 107686 106720 107738
rect 106744 107686 106774 107738
rect 106774 107686 106786 107738
rect 106786 107686 106800 107738
rect 106824 107686 106838 107738
rect 106838 107686 106850 107738
rect 106850 107686 106880 107738
rect 106904 107686 106914 107738
rect 106914 107686 106960 107738
rect 106664 107684 106720 107686
rect 106744 107684 106800 107686
rect 106824 107684 106880 107686
rect 106904 107684 106960 107686
rect 105928 107194 105984 107196
rect 106008 107194 106064 107196
rect 106088 107194 106144 107196
rect 106168 107194 106224 107196
rect 105928 107142 105974 107194
rect 105974 107142 105984 107194
rect 106008 107142 106038 107194
rect 106038 107142 106050 107194
rect 106050 107142 106064 107194
rect 106088 107142 106102 107194
rect 106102 107142 106114 107194
rect 106114 107142 106144 107194
rect 106168 107142 106178 107194
rect 106178 107142 106224 107194
rect 105928 107140 105984 107142
rect 106008 107140 106064 107142
rect 106088 107140 106144 107142
rect 106168 107140 106224 107142
rect 106664 106650 106720 106652
rect 106744 106650 106800 106652
rect 106824 106650 106880 106652
rect 106904 106650 106960 106652
rect 106664 106598 106710 106650
rect 106710 106598 106720 106650
rect 106744 106598 106774 106650
rect 106774 106598 106786 106650
rect 106786 106598 106800 106650
rect 106824 106598 106838 106650
rect 106838 106598 106850 106650
rect 106850 106598 106880 106650
rect 106904 106598 106914 106650
rect 106914 106598 106960 106650
rect 106664 106596 106720 106598
rect 106744 106596 106800 106598
rect 106824 106596 106880 106598
rect 106904 106596 106960 106598
rect 105928 106106 105984 106108
rect 106008 106106 106064 106108
rect 106088 106106 106144 106108
rect 106168 106106 106224 106108
rect 105928 106054 105974 106106
rect 105974 106054 105984 106106
rect 106008 106054 106038 106106
rect 106038 106054 106050 106106
rect 106050 106054 106064 106106
rect 106088 106054 106102 106106
rect 106102 106054 106114 106106
rect 106114 106054 106144 106106
rect 106168 106054 106178 106106
rect 106178 106054 106224 106106
rect 105928 106052 105984 106054
rect 106008 106052 106064 106054
rect 106088 106052 106144 106054
rect 106168 106052 106224 106054
rect 106664 105562 106720 105564
rect 106744 105562 106800 105564
rect 106824 105562 106880 105564
rect 106904 105562 106960 105564
rect 106664 105510 106710 105562
rect 106710 105510 106720 105562
rect 106744 105510 106774 105562
rect 106774 105510 106786 105562
rect 106786 105510 106800 105562
rect 106824 105510 106838 105562
rect 106838 105510 106850 105562
rect 106850 105510 106880 105562
rect 106904 105510 106914 105562
rect 106914 105510 106960 105562
rect 106664 105508 106720 105510
rect 106744 105508 106800 105510
rect 106824 105508 106880 105510
rect 106904 105508 106960 105510
rect 105928 105018 105984 105020
rect 106008 105018 106064 105020
rect 106088 105018 106144 105020
rect 106168 105018 106224 105020
rect 105928 104966 105974 105018
rect 105974 104966 105984 105018
rect 106008 104966 106038 105018
rect 106038 104966 106050 105018
rect 106050 104966 106064 105018
rect 106088 104966 106102 105018
rect 106102 104966 106114 105018
rect 106114 104966 106144 105018
rect 106168 104966 106178 105018
rect 106178 104966 106224 105018
rect 105928 104964 105984 104966
rect 106008 104964 106064 104966
rect 106088 104964 106144 104966
rect 106168 104964 106224 104966
rect 106664 104474 106720 104476
rect 106744 104474 106800 104476
rect 106824 104474 106880 104476
rect 106904 104474 106960 104476
rect 106664 104422 106710 104474
rect 106710 104422 106720 104474
rect 106744 104422 106774 104474
rect 106774 104422 106786 104474
rect 106786 104422 106800 104474
rect 106824 104422 106838 104474
rect 106838 104422 106850 104474
rect 106850 104422 106880 104474
rect 106904 104422 106914 104474
rect 106914 104422 106960 104474
rect 106664 104420 106720 104422
rect 106744 104420 106800 104422
rect 106824 104420 106880 104422
rect 106904 104420 106960 104422
rect 105928 103930 105984 103932
rect 106008 103930 106064 103932
rect 106088 103930 106144 103932
rect 106168 103930 106224 103932
rect 105928 103878 105974 103930
rect 105974 103878 105984 103930
rect 106008 103878 106038 103930
rect 106038 103878 106050 103930
rect 106050 103878 106064 103930
rect 106088 103878 106102 103930
rect 106102 103878 106114 103930
rect 106114 103878 106144 103930
rect 106168 103878 106178 103930
rect 106178 103878 106224 103930
rect 105928 103876 105984 103878
rect 106008 103876 106064 103878
rect 106088 103876 106144 103878
rect 106168 103876 106224 103878
rect 106664 103386 106720 103388
rect 106744 103386 106800 103388
rect 106824 103386 106880 103388
rect 106904 103386 106960 103388
rect 106664 103334 106710 103386
rect 106710 103334 106720 103386
rect 106744 103334 106774 103386
rect 106774 103334 106786 103386
rect 106786 103334 106800 103386
rect 106824 103334 106838 103386
rect 106838 103334 106850 103386
rect 106850 103334 106880 103386
rect 106904 103334 106914 103386
rect 106914 103334 106960 103386
rect 106664 103332 106720 103334
rect 106744 103332 106800 103334
rect 106824 103332 106880 103334
rect 106904 103332 106960 103334
rect 105928 102842 105984 102844
rect 106008 102842 106064 102844
rect 106088 102842 106144 102844
rect 106168 102842 106224 102844
rect 105928 102790 105974 102842
rect 105974 102790 105984 102842
rect 106008 102790 106038 102842
rect 106038 102790 106050 102842
rect 106050 102790 106064 102842
rect 106088 102790 106102 102842
rect 106102 102790 106114 102842
rect 106114 102790 106144 102842
rect 106168 102790 106178 102842
rect 106178 102790 106224 102842
rect 105928 102788 105984 102790
rect 106008 102788 106064 102790
rect 106088 102788 106144 102790
rect 106168 102788 106224 102790
rect 106664 102298 106720 102300
rect 106744 102298 106800 102300
rect 106824 102298 106880 102300
rect 106904 102298 106960 102300
rect 106664 102246 106710 102298
rect 106710 102246 106720 102298
rect 106744 102246 106774 102298
rect 106774 102246 106786 102298
rect 106786 102246 106800 102298
rect 106824 102246 106838 102298
rect 106838 102246 106850 102298
rect 106850 102246 106880 102298
rect 106904 102246 106914 102298
rect 106914 102246 106960 102298
rect 106664 102244 106720 102246
rect 106744 102244 106800 102246
rect 106824 102244 106880 102246
rect 106904 102244 106960 102246
rect 105928 101754 105984 101756
rect 106008 101754 106064 101756
rect 106088 101754 106144 101756
rect 106168 101754 106224 101756
rect 105928 101702 105974 101754
rect 105974 101702 105984 101754
rect 106008 101702 106038 101754
rect 106038 101702 106050 101754
rect 106050 101702 106064 101754
rect 106088 101702 106102 101754
rect 106102 101702 106114 101754
rect 106114 101702 106144 101754
rect 106168 101702 106178 101754
rect 106178 101702 106224 101754
rect 105928 101700 105984 101702
rect 106008 101700 106064 101702
rect 106088 101700 106144 101702
rect 106168 101700 106224 101702
rect 106664 101210 106720 101212
rect 106744 101210 106800 101212
rect 106824 101210 106880 101212
rect 106904 101210 106960 101212
rect 106664 101158 106710 101210
rect 106710 101158 106720 101210
rect 106744 101158 106774 101210
rect 106774 101158 106786 101210
rect 106786 101158 106800 101210
rect 106824 101158 106838 101210
rect 106838 101158 106850 101210
rect 106850 101158 106880 101210
rect 106904 101158 106914 101210
rect 106914 101158 106960 101210
rect 106664 101156 106720 101158
rect 106744 101156 106800 101158
rect 106824 101156 106880 101158
rect 106904 101156 106960 101158
rect 105928 100666 105984 100668
rect 106008 100666 106064 100668
rect 106088 100666 106144 100668
rect 106168 100666 106224 100668
rect 105928 100614 105974 100666
rect 105974 100614 105984 100666
rect 106008 100614 106038 100666
rect 106038 100614 106050 100666
rect 106050 100614 106064 100666
rect 106088 100614 106102 100666
rect 106102 100614 106114 100666
rect 106114 100614 106144 100666
rect 106168 100614 106178 100666
rect 106178 100614 106224 100666
rect 105928 100612 105984 100614
rect 106008 100612 106064 100614
rect 106088 100612 106144 100614
rect 106168 100612 106224 100614
rect 106664 100122 106720 100124
rect 106744 100122 106800 100124
rect 106824 100122 106880 100124
rect 106904 100122 106960 100124
rect 106664 100070 106710 100122
rect 106710 100070 106720 100122
rect 106744 100070 106774 100122
rect 106774 100070 106786 100122
rect 106786 100070 106800 100122
rect 106824 100070 106838 100122
rect 106838 100070 106850 100122
rect 106850 100070 106880 100122
rect 106904 100070 106914 100122
rect 106914 100070 106960 100122
rect 106664 100068 106720 100070
rect 106744 100068 106800 100070
rect 106824 100068 106880 100070
rect 106904 100068 106960 100070
rect 105928 99578 105984 99580
rect 106008 99578 106064 99580
rect 106088 99578 106144 99580
rect 106168 99578 106224 99580
rect 105928 99526 105974 99578
rect 105974 99526 105984 99578
rect 106008 99526 106038 99578
rect 106038 99526 106050 99578
rect 106050 99526 106064 99578
rect 106088 99526 106102 99578
rect 106102 99526 106114 99578
rect 106114 99526 106144 99578
rect 106168 99526 106178 99578
rect 106178 99526 106224 99578
rect 105928 99524 105984 99526
rect 106008 99524 106064 99526
rect 106088 99524 106144 99526
rect 106168 99524 106224 99526
rect 106664 99034 106720 99036
rect 106744 99034 106800 99036
rect 106824 99034 106880 99036
rect 106904 99034 106960 99036
rect 106664 98982 106710 99034
rect 106710 98982 106720 99034
rect 106744 98982 106774 99034
rect 106774 98982 106786 99034
rect 106786 98982 106800 99034
rect 106824 98982 106838 99034
rect 106838 98982 106850 99034
rect 106850 98982 106880 99034
rect 106904 98982 106914 99034
rect 106914 98982 106960 99034
rect 106664 98980 106720 98982
rect 106744 98980 106800 98982
rect 106824 98980 106880 98982
rect 106904 98980 106960 98982
rect 105928 98490 105984 98492
rect 106008 98490 106064 98492
rect 106088 98490 106144 98492
rect 106168 98490 106224 98492
rect 105928 98438 105974 98490
rect 105974 98438 105984 98490
rect 106008 98438 106038 98490
rect 106038 98438 106050 98490
rect 106050 98438 106064 98490
rect 106088 98438 106102 98490
rect 106102 98438 106114 98490
rect 106114 98438 106144 98490
rect 106168 98438 106178 98490
rect 106178 98438 106224 98490
rect 105928 98436 105984 98438
rect 106008 98436 106064 98438
rect 106088 98436 106144 98438
rect 106168 98436 106224 98438
rect 106664 97946 106720 97948
rect 106744 97946 106800 97948
rect 106824 97946 106880 97948
rect 106904 97946 106960 97948
rect 106664 97894 106710 97946
rect 106710 97894 106720 97946
rect 106744 97894 106774 97946
rect 106774 97894 106786 97946
rect 106786 97894 106800 97946
rect 106824 97894 106838 97946
rect 106838 97894 106850 97946
rect 106850 97894 106880 97946
rect 106904 97894 106914 97946
rect 106914 97894 106960 97946
rect 106664 97892 106720 97894
rect 106744 97892 106800 97894
rect 106824 97892 106880 97894
rect 106904 97892 106960 97894
rect 105928 97402 105984 97404
rect 106008 97402 106064 97404
rect 106088 97402 106144 97404
rect 106168 97402 106224 97404
rect 105928 97350 105974 97402
rect 105974 97350 105984 97402
rect 106008 97350 106038 97402
rect 106038 97350 106050 97402
rect 106050 97350 106064 97402
rect 106088 97350 106102 97402
rect 106102 97350 106114 97402
rect 106114 97350 106144 97402
rect 106168 97350 106178 97402
rect 106178 97350 106224 97402
rect 105928 97348 105984 97350
rect 106008 97348 106064 97350
rect 106088 97348 106144 97350
rect 106168 97348 106224 97350
rect 106664 96858 106720 96860
rect 106744 96858 106800 96860
rect 106824 96858 106880 96860
rect 106904 96858 106960 96860
rect 106664 96806 106710 96858
rect 106710 96806 106720 96858
rect 106744 96806 106774 96858
rect 106774 96806 106786 96858
rect 106786 96806 106800 96858
rect 106824 96806 106838 96858
rect 106838 96806 106850 96858
rect 106850 96806 106880 96858
rect 106904 96806 106914 96858
rect 106914 96806 106960 96858
rect 106664 96804 106720 96806
rect 106744 96804 106800 96806
rect 106824 96804 106880 96806
rect 106904 96804 106960 96806
rect 105928 96314 105984 96316
rect 106008 96314 106064 96316
rect 106088 96314 106144 96316
rect 106168 96314 106224 96316
rect 105928 96262 105974 96314
rect 105974 96262 105984 96314
rect 106008 96262 106038 96314
rect 106038 96262 106050 96314
rect 106050 96262 106064 96314
rect 106088 96262 106102 96314
rect 106102 96262 106114 96314
rect 106114 96262 106144 96314
rect 106168 96262 106178 96314
rect 106178 96262 106224 96314
rect 105928 96260 105984 96262
rect 106008 96260 106064 96262
rect 106088 96260 106144 96262
rect 106168 96260 106224 96262
rect 106664 95770 106720 95772
rect 106744 95770 106800 95772
rect 106824 95770 106880 95772
rect 106904 95770 106960 95772
rect 106664 95718 106710 95770
rect 106710 95718 106720 95770
rect 106744 95718 106774 95770
rect 106774 95718 106786 95770
rect 106786 95718 106800 95770
rect 106824 95718 106838 95770
rect 106838 95718 106850 95770
rect 106850 95718 106880 95770
rect 106904 95718 106914 95770
rect 106914 95718 106960 95770
rect 106664 95716 106720 95718
rect 106744 95716 106800 95718
rect 106824 95716 106880 95718
rect 106904 95716 106960 95718
rect 105928 95226 105984 95228
rect 106008 95226 106064 95228
rect 106088 95226 106144 95228
rect 106168 95226 106224 95228
rect 105928 95174 105974 95226
rect 105974 95174 105984 95226
rect 106008 95174 106038 95226
rect 106038 95174 106050 95226
rect 106050 95174 106064 95226
rect 106088 95174 106102 95226
rect 106102 95174 106114 95226
rect 106114 95174 106144 95226
rect 106168 95174 106178 95226
rect 106178 95174 106224 95226
rect 105928 95172 105984 95174
rect 106008 95172 106064 95174
rect 106088 95172 106144 95174
rect 106168 95172 106224 95174
rect 106664 94682 106720 94684
rect 106744 94682 106800 94684
rect 106824 94682 106880 94684
rect 106904 94682 106960 94684
rect 106664 94630 106710 94682
rect 106710 94630 106720 94682
rect 106744 94630 106774 94682
rect 106774 94630 106786 94682
rect 106786 94630 106800 94682
rect 106824 94630 106838 94682
rect 106838 94630 106850 94682
rect 106850 94630 106880 94682
rect 106904 94630 106914 94682
rect 106914 94630 106960 94682
rect 106664 94628 106720 94630
rect 106744 94628 106800 94630
rect 106824 94628 106880 94630
rect 106904 94628 106960 94630
rect 105928 94138 105984 94140
rect 106008 94138 106064 94140
rect 106088 94138 106144 94140
rect 106168 94138 106224 94140
rect 105928 94086 105974 94138
rect 105974 94086 105984 94138
rect 106008 94086 106038 94138
rect 106038 94086 106050 94138
rect 106050 94086 106064 94138
rect 106088 94086 106102 94138
rect 106102 94086 106114 94138
rect 106114 94086 106144 94138
rect 106168 94086 106178 94138
rect 106178 94086 106224 94138
rect 105928 94084 105984 94086
rect 106008 94084 106064 94086
rect 106088 94084 106144 94086
rect 106168 94084 106224 94086
rect 106664 93594 106720 93596
rect 106744 93594 106800 93596
rect 106824 93594 106880 93596
rect 106904 93594 106960 93596
rect 106664 93542 106710 93594
rect 106710 93542 106720 93594
rect 106744 93542 106774 93594
rect 106774 93542 106786 93594
rect 106786 93542 106800 93594
rect 106824 93542 106838 93594
rect 106838 93542 106850 93594
rect 106850 93542 106880 93594
rect 106904 93542 106914 93594
rect 106914 93542 106960 93594
rect 106664 93540 106720 93542
rect 106744 93540 106800 93542
rect 106824 93540 106880 93542
rect 106904 93540 106960 93542
rect 105928 93050 105984 93052
rect 106008 93050 106064 93052
rect 106088 93050 106144 93052
rect 106168 93050 106224 93052
rect 105928 92998 105974 93050
rect 105974 92998 105984 93050
rect 106008 92998 106038 93050
rect 106038 92998 106050 93050
rect 106050 92998 106064 93050
rect 106088 92998 106102 93050
rect 106102 92998 106114 93050
rect 106114 92998 106144 93050
rect 106168 92998 106178 93050
rect 106178 92998 106224 93050
rect 105928 92996 105984 92998
rect 106008 92996 106064 92998
rect 106088 92996 106144 92998
rect 106168 92996 106224 92998
rect 106664 92506 106720 92508
rect 106744 92506 106800 92508
rect 106824 92506 106880 92508
rect 106904 92506 106960 92508
rect 106664 92454 106710 92506
rect 106710 92454 106720 92506
rect 106744 92454 106774 92506
rect 106774 92454 106786 92506
rect 106786 92454 106800 92506
rect 106824 92454 106838 92506
rect 106838 92454 106850 92506
rect 106850 92454 106880 92506
rect 106904 92454 106914 92506
rect 106914 92454 106960 92506
rect 106664 92452 106720 92454
rect 106744 92452 106800 92454
rect 106824 92452 106880 92454
rect 106904 92452 106960 92454
rect 105928 91962 105984 91964
rect 106008 91962 106064 91964
rect 106088 91962 106144 91964
rect 106168 91962 106224 91964
rect 105928 91910 105974 91962
rect 105974 91910 105984 91962
rect 106008 91910 106038 91962
rect 106038 91910 106050 91962
rect 106050 91910 106064 91962
rect 106088 91910 106102 91962
rect 106102 91910 106114 91962
rect 106114 91910 106144 91962
rect 106168 91910 106178 91962
rect 106178 91910 106224 91962
rect 105928 91908 105984 91910
rect 106008 91908 106064 91910
rect 106088 91908 106144 91910
rect 106168 91908 106224 91910
rect 106664 91418 106720 91420
rect 106744 91418 106800 91420
rect 106824 91418 106880 91420
rect 106904 91418 106960 91420
rect 106664 91366 106710 91418
rect 106710 91366 106720 91418
rect 106744 91366 106774 91418
rect 106774 91366 106786 91418
rect 106786 91366 106800 91418
rect 106824 91366 106838 91418
rect 106838 91366 106850 91418
rect 106850 91366 106880 91418
rect 106904 91366 106914 91418
rect 106914 91366 106960 91418
rect 106664 91364 106720 91366
rect 106744 91364 106800 91366
rect 106824 91364 106880 91366
rect 106904 91364 106960 91366
rect 103978 77424 104034 77480
rect 105928 90874 105984 90876
rect 106008 90874 106064 90876
rect 106088 90874 106144 90876
rect 106168 90874 106224 90876
rect 105928 90822 105974 90874
rect 105974 90822 105984 90874
rect 106008 90822 106038 90874
rect 106038 90822 106050 90874
rect 106050 90822 106064 90874
rect 106088 90822 106102 90874
rect 106102 90822 106114 90874
rect 106114 90822 106144 90874
rect 106168 90822 106178 90874
rect 106178 90822 106224 90874
rect 105928 90820 105984 90822
rect 106008 90820 106064 90822
rect 106088 90820 106144 90822
rect 106168 90820 106224 90822
rect 106664 90330 106720 90332
rect 106744 90330 106800 90332
rect 106824 90330 106880 90332
rect 106904 90330 106960 90332
rect 106664 90278 106710 90330
rect 106710 90278 106720 90330
rect 106744 90278 106774 90330
rect 106774 90278 106786 90330
rect 106786 90278 106800 90330
rect 106824 90278 106838 90330
rect 106838 90278 106850 90330
rect 106850 90278 106880 90330
rect 106904 90278 106914 90330
rect 106914 90278 106960 90330
rect 106664 90276 106720 90278
rect 106744 90276 106800 90278
rect 106824 90276 106880 90278
rect 106904 90276 106960 90278
rect 105928 89786 105984 89788
rect 106008 89786 106064 89788
rect 106088 89786 106144 89788
rect 106168 89786 106224 89788
rect 105928 89734 105974 89786
rect 105974 89734 105984 89786
rect 106008 89734 106038 89786
rect 106038 89734 106050 89786
rect 106050 89734 106064 89786
rect 106088 89734 106102 89786
rect 106102 89734 106114 89786
rect 106114 89734 106144 89786
rect 106168 89734 106178 89786
rect 106178 89734 106224 89786
rect 105928 89732 105984 89734
rect 106008 89732 106064 89734
rect 106088 89732 106144 89734
rect 106168 89732 106224 89734
rect 106664 89242 106720 89244
rect 106744 89242 106800 89244
rect 106824 89242 106880 89244
rect 106904 89242 106960 89244
rect 106664 89190 106710 89242
rect 106710 89190 106720 89242
rect 106744 89190 106774 89242
rect 106774 89190 106786 89242
rect 106786 89190 106800 89242
rect 106824 89190 106838 89242
rect 106838 89190 106850 89242
rect 106850 89190 106880 89242
rect 106904 89190 106914 89242
rect 106914 89190 106960 89242
rect 106664 89188 106720 89190
rect 106744 89188 106800 89190
rect 106824 89188 106880 89190
rect 106904 89188 106960 89190
rect 105928 88698 105984 88700
rect 106008 88698 106064 88700
rect 106088 88698 106144 88700
rect 106168 88698 106224 88700
rect 105928 88646 105974 88698
rect 105974 88646 105984 88698
rect 106008 88646 106038 88698
rect 106038 88646 106050 88698
rect 106050 88646 106064 88698
rect 106088 88646 106102 88698
rect 106102 88646 106114 88698
rect 106114 88646 106144 88698
rect 106168 88646 106178 88698
rect 106178 88646 106224 88698
rect 105928 88644 105984 88646
rect 106008 88644 106064 88646
rect 106088 88644 106144 88646
rect 106168 88644 106224 88646
rect 106664 88154 106720 88156
rect 106744 88154 106800 88156
rect 106824 88154 106880 88156
rect 106904 88154 106960 88156
rect 106664 88102 106710 88154
rect 106710 88102 106720 88154
rect 106744 88102 106774 88154
rect 106774 88102 106786 88154
rect 106786 88102 106800 88154
rect 106824 88102 106838 88154
rect 106838 88102 106850 88154
rect 106850 88102 106880 88154
rect 106904 88102 106914 88154
rect 106914 88102 106960 88154
rect 106664 88100 106720 88102
rect 106744 88100 106800 88102
rect 106824 88100 106880 88102
rect 106904 88100 106960 88102
rect 105928 87610 105984 87612
rect 106008 87610 106064 87612
rect 106088 87610 106144 87612
rect 106168 87610 106224 87612
rect 105928 87558 105974 87610
rect 105974 87558 105984 87610
rect 106008 87558 106038 87610
rect 106038 87558 106050 87610
rect 106050 87558 106064 87610
rect 106088 87558 106102 87610
rect 106102 87558 106114 87610
rect 106114 87558 106144 87610
rect 106168 87558 106178 87610
rect 106178 87558 106224 87610
rect 105928 87556 105984 87558
rect 106008 87556 106064 87558
rect 106088 87556 106144 87558
rect 106168 87556 106224 87558
rect 106664 87066 106720 87068
rect 106744 87066 106800 87068
rect 106824 87066 106880 87068
rect 106904 87066 106960 87068
rect 106664 87014 106710 87066
rect 106710 87014 106720 87066
rect 106744 87014 106774 87066
rect 106774 87014 106786 87066
rect 106786 87014 106800 87066
rect 106824 87014 106838 87066
rect 106838 87014 106850 87066
rect 106850 87014 106880 87066
rect 106904 87014 106914 87066
rect 106914 87014 106960 87066
rect 106664 87012 106720 87014
rect 106744 87012 106800 87014
rect 106824 87012 106880 87014
rect 106904 87012 106960 87014
rect 105928 86522 105984 86524
rect 106008 86522 106064 86524
rect 106088 86522 106144 86524
rect 106168 86522 106224 86524
rect 105928 86470 105974 86522
rect 105974 86470 105984 86522
rect 106008 86470 106038 86522
rect 106038 86470 106050 86522
rect 106050 86470 106064 86522
rect 106088 86470 106102 86522
rect 106102 86470 106114 86522
rect 106114 86470 106144 86522
rect 106168 86470 106178 86522
rect 106178 86470 106224 86522
rect 105928 86468 105984 86470
rect 106008 86468 106064 86470
rect 106088 86468 106144 86470
rect 106168 86468 106224 86470
rect 106664 85978 106720 85980
rect 106744 85978 106800 85980
rect 106824 85978 106880 85980
rect 106904 85978 106960 85980
rect 106664 85926 106710 85978
rect 106710 85926 106720 85978
rect 106744 85926 106774 85978
rect 106774 85926 106786 85978
rect 106786 85926 106800 85978
rect 106824 85926 106838 85978
rect 106838 85926 106850 85978
rect 106850 85926 106880 85978
rect 106904 85926 106914 85978
rect 106914 85926 106960 85978
rect 106664 85924 106720 85926
rect 106744 85924 106800 85926
rect 106824 85924 106880 85926
rect 106904 85924 106960 85926
rect 105928 85434 105984 85436
rect 106008 85434 106064 85436
rect 106088 85434 106144 85436
rect 106168 85434 106224 85436
rect 105928 85382 105974 85434
rect 105974 85382 105984 85434
rect 106008 85382 106038 85434
rect 106038 85382 106050 85434
rect 106050 85382 106064 85434
rect 106088 85382 106102 85434
rect 106102 85382 106114 85434
rect 106114 85382 106144 85434
rect 106168 85382 106178 85434
rect 106178 85382 106224 85434
rect 105928 85380 105984 85382
rect 106008 85380 106064 85382
rect 106088 85380 106144 85382
rect 106168 85380 106224 85382
rect 106664 84890 106720 84892
rect 106744 84890 106800 84892
rect 106824 84890 106880 84892
rect 106904 84890 106960 84892
rect 106664 84838 106710 84890
rect 106710 84838 106720 84890
rect 106744 84838 106774 84890
rect 106774 84838 106786 84890
rect 106786 84838 106800 84890
rect 106824 84838 106838 84890
rect 106838 84838 106850 84890
rect 106850 84838 106880 84890
rect 106904 84838 106914 84890
rect 106914 84838 106960 84890
rect 106664 84836 106720 84838
rect 106744 84836 106800 84838
rect 106824 84836 106880 84838
rect 106904 84836 106960 84838
rect 105928 84346 105984 84348
rect 106008 84346 106064 84348
rect 106088 84346 106144 84348
rect 106168 84346 106224 84348
rect 105928 84294 105974 84346
rect 105974 84294 105984 84346
rect 106008 84294 106038 84346
rect 106038 84294 106050 84346
rect 106050 84294 106064 84346
rect 106088 84294 106102 84346
rect 106102 84294 106114 84346
rect 106114 84294 106144 84346
rect 106168 84294 106178 84346
rect 106178 84294 106224 84346
rect 105928 84292 105984 84294
rect 106008 84292 106064 84294
rect 106088 84292 106144 84294
rect 106168 84292 106224 84294
rect 106664 83802 106720 83804
rect 106744 83802 106800 83804
rect 106824 83802 106880 83804
rect 106904 83802 106960 83804
rect 106664 83750 106710 83802
rect 106710 83750 106720 83802
rect 106744 83750 106774 83802
rect 106774 83750 106786 83802
rect 106786 83750 106800 83802
rect 106824 83750 106838 83802
rect 106838 83750 106850 83802
rect 106850 83750 106880 83802
rect 106904 83750 106914 83802
rect 106914 83750 106960 83802
rect 106664 83748 106720 83750
rect 106744 83748 106800 83750
rect 106824 83748 106880 83750
rect 106904 83748 106960 83750
rect 105928 83258 105984 83260
rect 106008 83258 106064 83260
rect 106088 83258 106144 83260
rect 106168 83258 106224 83260
rect 105928 83206 105974 83258
rect 105974 83206 105984 83258
rect 106008 83206 106038 83258
rect 106038 83206 106050 83258
rect 106050 83206 106064 83258
rect 106088 83206 106102 83258
rect 106102 83206 106114 83258
rect 106114 83206 106144 83258
rect 106168 83206 106178 83258
rect 106178 83206 106224 83258
rect 105928 83204 105984 83206
rect 106008 83204 106064 83206
rect 106088 83204 106144 83206
rect 106168 83204 106224 83206
rect 106664 82714 106720 82716
rect 106744 82714 106800 82716
rect 106824 82714 106880 82716
rect 106904 82714 106960 82716
rect 106664 82662 106710 82714
rect 106710 82662 106720 82714
rect 106744 82662 106774 82714
rect 106774 82662 106786 82714
rect 106786 82662 106800 82714
rect 106824 82662 106838 82714
rect 106838 82662 106850 82714
rect 106850 82662 106880 82714
rect 106904 82662 106914 82714
rect 106914 82662 106960 82714
rect 106664 82660 106720 82662
rect 106744 82660 106800 82662
rect 106824 82660 106880 82662
rect 106904 82660 106960 82662
rect 105928 82170 105984 82172
rect 106008 82170 106064 82172
rect 106088 82170 106144 82172
rect 106168 82170 106224 82172
rect 105928 82118 105974 82170
rect 105974 82118 105984 82170
rect 106008 82118 106038 82170
rect 106038 82118 106050 82170
rect 106050 82118 106064 82170
rect 106088 82118 106102 82170
rect 106102 82118 106114 82170
rect 106114 82118 106144 82170
rect 106168 82118 106178 82170
rect 106178 82118 106224 82170
rect 105928 82116 105984 82118
rect 106008 82116 106064 82118
rect 106088 82116 106144 82118
rect 106168 82116 106224 82118
rect 106664 81626 106720 81628
rect 106744 81626 106800 81628
rect 106824 81626 106880 81628
rect 106904 81626 106960 81628
rect 106664 81574 106710 81626
rect 106710 81574 106720 81626
rect 106744 81574 106774 81626
rect 106774 81574 106786 81626
rect 106786 81574 106800 81626
rect 106824 81574 106838 81626
rect 106838 81574 106850 81626
rect 106850 81574 106880 81626
rect 106904 81574 106914 81626
rect 106914 81574 106960 81626
rect 106664 81572 106720 81574
rect 106744 81572 106800 81574
rect 106824 81572 106880 81574
rect 106904 81572 106960 81574
rect 105928 81082 105984 81084
rect 106008 81082 106064 81084
rect 106088 81082 106144 81084
rect 106168 81082 106224 81084
rect 105928 81030 105974 81082
rect 105974 81030 105984 81082
rect 106008 81030 106038 81082
rect 106038 81030 106050 81082
rect 106050 81030 106064 81082
rect 106088 81030 106102 81082
rect 106102 81030 106114 81082
rect 106114 81030 106144 81082
rect 106168 81030 106178 81082
rect 106178 81030 106224 81082
rect 105928 81028 105984 81030
rect 106008 81028 106064 81030
rect 106088 81028 106144 81030
rect 106168 81028 106224 81030
rect 106664 80538 106720 80540
rect 106744 80538 106800 80540
rect 106824 80538 106880 80540
rect 106904 80538 106960 80540
rect 106664 80486 106710 80538
rect 106710 80486 106720 80538
rect 106744 80486 106774 80538
rect 106774 80486 106786 80538
rect 106786 80486 106800 80538
rect 106824 80486 106838 80538
rect 106838 80486 106850 80538
rect 106850 80486 106880 80538
rect 106904 80486 106914 80538
rect 106914 80486 106960 80538
rect 106664 80484 106720 80486
rect 106744 80484 106800 80486
rect 106824 80484 106880 80486
rect 106904 80484 106960 80486
rect 105928 79994 105984 79996
rect 106008 79994 106064 79996
rect 106088 79994 106144 79996
rect 106168 79994 106224 79996
rect 105928 79942 105974 79994
rect 105974 79942 105984 79994
rect 106008 79942 106038 79994
rect 106038 79942 106050 79994
rect 106050 79942 106064 79994
rect 106088 79942 106102 79994
rect 106102 79942 106114 79994
rect 106114 79942 106144 79994
rect 106168 79942 106178 79994
rect 106178 79942 106224 79994
rect 105928 79940 105984 79942
rect 106008 79940 106064 79942
rect 106088 79940 106144 79942
rect 106168 79940 106224 79942
rect 106664 79450 106720 79452
rect 106744 79450 106800 79452
rect 106824 79450 106880 79452
rect 106904 79450 106960 79452
rect 106664 79398 106710 79450
rect 106710 79398 106720 79450
rect 106744 79398 106774 79450
rect 106774 79398 106786 79450
rect 106786 79398 106800 79450
rect 106824 79398 106838 79450
rect 106838 79398 106850 79450
rect 106850 79398 106880 79450
rect 106904 79398 106914 79450
rect 106914 79398 106960 79450
rect 106664 79396 106720 79398
rect 106744 79396 106800 79398
rect 106824 79396 106880 79398
rect 106904 79396 106960 79398
rect 108486 78956 108488 78976
rect 108488 78956 108540 78976
rect 108540 78956 108542 78976
rect 108486 78920 108542 78956
rect 105928 78906 105984 78908
rect 106008 78906 106064 78908
rect 106088 78906 106144 78908
rect 106168 78906 106224 78908
rect 105928 78854 105974 78906
rect 105974 78854 105984 78906
rect 106008 78854 106038 78906
rect 106038 78854 106050 78906
rect 106050 78854 106064 78906
rect 106088 78854 106102 78906
rect 106102 78854 106114 78906
rect 106114 78854 106144 78906
rect 106168 78854 106178 78906
rect 106178 78854 106224 78906
rect 105928 78852 105984 78854
rect 106008 78852 106064 78854
rect 106088 78852 106144 78854
rect 106168 78852 106224 78854
rect 106664 78362 106720 78364
rect 106744 78362 106800 78364
rect 106824 78362 106880 78364
rect 106904 78362 106960 78364
rect 106664 78310 106710 78362
rect 106710 78310 106720 78362
rect 106744 78310 106774 78362
rect 106774 78310 106786 78362
rect 106786 78310 106800 78362
rect 106824 78310 106838 78362
rect 106838 78310 106850 78362
rect 106850 78310 106880 78362
rect 106904 78310 106914 78362
rect 106914 78310 106960 78362
rect 106664 78308 106720 78310
rect 106744 78308 106800 78310
rect 106824 78308 106880 78310
rect 106904 78308 106960 78310
rect 105928 77818 105984 77820
rect 106008 77818 106064 77820
rect 106088 77818 106144 77820
rect 106168 77818 106224 77820
rect 105928 77766 105974 77818
rect 105974 77766 105984 77818
rect 106008 77766 106038 77818
rect 106038 77766 106050 77818
rect 106050 77766 106064 77818
rect 106088 77766 106102 77818
rect 106102 77766 106114 77818
rect 106114 77766 106144 77818
rect 106168 77766 106178 77818
rect 106178 77766 106224 77818
rect 105928 77764 105984 77766
rect 106008 77764 106064 77766
rect 106088 77764 106144 77766
rect 106168 77764 106224 77766
rect 106664 77274 106720 77276
rect 106744 77274 106800 77276
rect 106824 77274 106880 77276
rect 106904 77274 106960 77276
rect 106664 77222 106710 77274
rect 106710 77222 106720 77274
rect 106744 77222 106774 77274
rect 106774 77222 106786 77274
rect 106786 77222 106800 77274
rect 106824 77222 106838 77274
rect 106838 77222 106850 77274
rect 106850 77222 106880 77274
rect 106904 77222 106914 77274
rect 106914 77222 106960 77274
rect 106664 77220 106720 77222
rect 106744 77220 106800 77222
rect 106824 77220 106880 77222
rect 106904 77220 106960 77222
rect 108486 78240 108542 78296
rect 108486 77560 108542 77616
rect 108486 76900 108542 76936
rect 108486 76880 108488 76900
rect 108488 76880 108540 76900
rect 108540 76880 108542 76900
rect 108486 76236 108488 76256
rect 108488 76236 108540 76256
rect 108540 76236 108542 76256
rect 108486 76200 108542 76236
rect 108486 75520 108542 75576
rect 108486 74840 108542 74896
rect 108486 74160 108542 74216
rect 108486 73516 108488 73536
rect 108488 73516 108540 73536
rect 108540 73516 108542 73536
rect 108486 73480 108542 73516
rect 108486 72800 108542 72856
rect 108486 67360 108542 67416
rect 102230 25032 102286 25088
rect 106664 66394 106720 66396
rect 106744 66394 106800 66396
rect 106824 66394 106880 66396
rect 106904 66394 106960 66396
rect 106664 66342 106710 66394
rect 106710 66342 106720 66394
rect 106744 66342 106774 66394
rect 106774 66342 106786 66394
rect 106786 66342 106800 66394
rect 106824 66342 106838 66394
rect 106838 66342 106850 66394
rect 106850 66342 106880 66394
rect 106904 66342 106914 66394
rect 106914 66342 106960 66394
rect 106664 66340 106720 66342
rect 106744 66340 106800 66342
rect 106824 66340 106880 66342
rect 106904 66340 106960 66342
rect 105928 65850 105984 65852
rect 106008 65850 106064 65852
rect 106088 65850 106144 65852
rect 106168 65850 106224 65852
rect 105928 65798 105974 65850
rect 105974 65798 105984 65850
rect 106008 65798 106038 65850
rect 106038 65798 106050 65850
rect 106050 65798 106064 65850
rect 106088 65798 106102 65850
rect 106102 65798 106114 65850
rect 106114 65798 106144 65850
rect 106168 65798 106178 65850
rect 106178 65798 106224 65850
rect 105928 65796 105984 65798
rect 106008 65796 106064 65798
rect 106088 65796 106144 65798
rect 106168 65796 106224 65798
rect 102598 25100 102600 25120
rect 102600 25100 102652 25120
rect 102652 25100 102654 25120
rect 102598 25064 102654 25100
rect 102322 22204 102378 22260
rect 106664 65306 106720 65308
rect 106744 65306 106800 65308
rect 106824 65306 106880 65308
rect 106904 65306 106960 65308
rect 106664 65254 106710 65306
rect 106710 65254 106720 65306
rect 106744 65254 106774 65306
rect 106774 65254 106786 65306
rect 106786 65254 106800 65306
rect 106824 65254 106838 65306
rect 106838 65254 106850 65306
rect 106850 65254 106880 65306
rect 106904 65254 106914 65306
rect 106914 65254 106960 65306
rect 106664 65252 106720 65254
rect 106744 65252 106800 65254
rect 106824 65252 106880 65254
rect 106904 65252 106960 65254
rect 105928 64762 105984 64764
rect 106008 64762 106064 64764
rect 106088 64762 106144 64764
rect 106168 64762 106224 64764
rect 105928 64710 105974 64762
rect 105974 64710 105984 64762
rect 106008 64710 106038 64762
rect 106038 64710 106050 64762
rect 106050 64710 106064 64762
rect 106088 64710 106102 64762
rect 106102 64710 106114 64762
rect 106114 64710 106144 64762
rect 106168 64710 106178 64762
rect 106178 64710 106224 64762
rect 105928 64708 105984 64710
rect 106008 64708 106064 64710
rect 106088 64708 106144 64710
rect 106168 64708 106224 64710
rect 106664 64218 106720 64220
rect 106744 64218 106800 64220
rect 106824 64218 106880 64220
rect 106904 64218 106960 64220
rect 106664 64166 106710 64218
rect 106710 64166 106720 64218
rect 106744 64166 106774 64218
rect 106774 64166 106786 64218
rect 106786 64166 106800 64218
rect 106824 64166 106838 64218
rect 106838 64166 106850 64218
rect 106850 64166 106880 64218
rect 106904 64166 106914 64218
rect 106914 64166 106960 64218
rect 106664 64164 106720 64166
rect 106744 64164 106800 64166
rect 106824 64164 106880 64166
rect 106904 64164 106960 64166
rect 105928 63674 105984 63676
rect 106008 63674 106064 63676
rect 106088 63674 106144 63676
rect 106168 63674 106224 63676
rect 105928 63622 105974 63674
rect 105974 63622 105984 63674
rect 106008 63622 106038 63674
rect 106038 63622 106050 63674
rect 106050 63622 106064 63674
rect 106088 63622 106102 63674
rect 106102 63622 106114 63674
rect 106114 63622 106144 63674
rect 106168 63622 106178 63674
rect 106178 63622 106224 63674
rect 105928 63620 105984 63622
rect 106008 63620 106064 63622
rect 106088 63620 106144 63622
rect 106168 63620 106224 63622
rect 106664 63130 106720 63132
rect 106744 63130 106800 63132
rect 106824 63130 106880 63132
rect 106904 63130 106960 63132
rect 106664 63078 106710 63130
rect 106710 63078 106720 63130
rect 106744 63078 106774 63130
rect 106774 63078 106786 63130
rect 106786 63078 106800 63130
rect 106824 63078 106838 63130
rect 106838 63078 106850 63130
rect 106850 63078 106880 63130
rect 106904 63078 106914 63130
rect 106914 63078 106960 63130
rect 106664 63076 106720 63078
rect 106744 63076 106800 63078
rect 106824 63076 106880 63078
rect 106904 63076 106960 63078
rect 105928 62586 105984 62588
rect 106008 62586 106064 62588
rect 106088 62586 106144 62588
rect 106168 62586 106224 62588
rect 105928 62534 105974 62586
rect 105974 62534 105984 62586
rect 106008 62534 106038 62586
rect 106038 62534 106050 62586
rect 106050 62534 106064 62586
rect 106088 62534 106102 62586
rect 106102 62534 106114 62586
rect 106114 62534 106144 62586
rect 106168 62534 106178 62586
rect 106178 62534 106224 62586
rect 105928 62532 105984 62534
rect 106008 62532 106064 62534
rect 106088 62532 106144 62534
rect 106168 62532 106224 62534
rect 106664 62042 106720 62044
rect 106744 62042 106800 62044
rect 106824 62042 106880 62044
rect 106904 62042 106960 62044
rect 106664 61990 106710 62042
rect 106710 61990 106720 62042
rect 106744 61990 106774 62042
rect 106774 61990 106786 62042
rect 106786 61990 106800 62042
rect 106824 61990 106838 62042
rect 106838 61990 106850 62042
rect 106850 61990 106880 62042
rect 106904 61990 106914 62042
rect 106914 61990 106960 62042
rect 106664 61988 106720 61990
rect 106744 61988 106800 61990
rect 106824 61988 106880 61990
rect 106904 61988 106960 61990
rect 105928 61498 105984 61500
rect 106008 61498 106064 61500
rect 106088 61498 106144 61500
rect 106168 61498 106224 61500
rect 105928 61446 105974 61498
rect 105974 61446 105984 61498
rect 106008 61446 106038 61498
rect 106038 61446 106050 61498
rect 106050 61446 106064 61498
rect 106088 61446 106102 61498
rect 106102 61446 106114 61498
rect 106114 61446 106144 61498
rect 106168 61446 106178 61498
rect 106178 61446 106224 61498
rect 105928 61444 105984 61446
rect 106008 61444 106064 61446
rect 106088 61444 106144 61446
rect 106168 61444 106224 61446
rect 106664 60954 106720 60956
rect 106744 60954 106800 60956
rect 106824 60954 106880 60956
rect 106904 60954 106960 60956
rect 106664 60902 106710 60954
rect 106710 60902 106720 60954
rect 106744 60902 106774 60954
rect 106774 60902 106786 60954
rect 106786 60902 106800 60954
rect 106824 60902 106838 60954
rect 106838 60902 106850 60954
rect 106850 60902 106880 60954
rect 106904 60902 106914 60954
rect 106914 60902 106960 60954
rect 106664 60900 106720 60902
rect 106744 60900 106800 60902
rect 106824 60900 106880 60902
rect 106904 60900 106960 60902
rect 105928 60410 105984 60412
rect 106008 60410 106064 60412
rect 106088 60410 106144 60412
rect 106168 60410 106224 60412
rect 105928 60358 105974 60410
rect 105974 60358 105984 60410
rect 106008 60358 106038 60410
rect 106038 60358 106050 60410
rect 106050 60358 106064 60410
rect 106088 60358 106102 60410
rect 106102 60358 106114 60410
rect 106114 60358 106144 60410
rect 106168 60358 106178 60410
rect 106178 60358 106224 60410
rect 105928 60356 105984 60358
rect 106008 60356 106064 60358
rect 106088 60356 106144 60358
rect 106168 60356 106224 60358
rect 106664 59866 106720 59868
rect 106744 59866 106800 59868
rect 106824 59866 106880 59868
rect 106904 59866 106960 59868
rect 106664 59814 106710 59866
rect 106710 59814 106720 59866
rect 106744 59814 106774 59866
rect 106774 59814 106786 59866
rect 106786 59814 106800 59866
rect 106824 59814 106838 59866
rect 106838 59814 106850 59866
rect 106850 59814 106880 59866
rect 106904 59814 106914 59866
rect 106914 59814 106960 59866
rect 106664 59812 106720 59814
rect 106744 59812 106800 59814
rect 106824 59812 106880 59814
rect 106904 59812 106960 59814
rect 104346 59744 104402 59800
rect 105928 59322 105984 59324
rect 106008 59322 106064 59324
rect 106088 59322 106144 59324
rect 106168 59322 106224 59324
rect 105928 59270 105974 59322
rect 105974 59270 105984 59322
rect 106008 59270 106038 59322
rect 106038 59270 106050 59322
rect 106050 59270 106064 59322
rect 106088 59270 106102 59322
rect 106102 59270 106114 59322
rect 106114 59270 106144 59322
rect 106168 59270 106178 59322
rect 106178 59270 106224 59322
rect 105928 59268 105984 59270
rect 106008 59268 106064 59270
rect 106088 59268 106144 59270
rect 106168 59268 106224 59270
rect 106664 58778 106720 58780
rect 106744 58778 106800 58780
rect 106824 58778 106880 58780
rect 106904 58778 106960 58780
rect 106664 58726 106710 58778
rect 106710 58726 106720 58778
rect 106744 58726 106774 58778
rect 106774 58726 106786 58778
rect 106786 58726 106800 58778
rect 106824 58726 106838 58778
rect 106838 58726 106850 58778
rect 106850 58726 106880 58778
rect 106904 58726 106914 58778
rect 106914 58726 106960 58778
rect 106664 58724 106720 58726
rect 106744 58724 106800 58726
rect 106824 58724 106880 58726
rect 106904 58724 106960 58726
rect 105928 58234 105984 58236
rect 106008 58234 106064 58236
rect 106088 58234 106144 58236
rect 106168 58234 106224 58236
rect 105928 58182 105974 58234
rect 105974 58182 105984 58234
rect 106008 58182 106038 58234
rect 106038 58182 106050 58234
rect 106050 58182 106064 58234
rect 106088 58182 106102 58234
rect 106102 58182 106114 58234
rect 106114 58182 106144 58234
rect 106168 58182 106178 58234
rect 106178 58182 106224 58234
rect 105928 58180 105984 58182
rect 106008 58180 106064 58182
rect 106088 58180 106144 58182
rect 106168 58180 106224 58182
rect 106664 57690 106720 57692
rect 106744 57690 106800 57692
rect 106824 57690 106880 57692
rect 106904 57690 106960 57692
rect 106664 57638 106710 57690
rect 106710 57638 106720 57690
rect 106744 57638 106774 57690
rect 106774 57638 106786 57690
rect 106786 57638 106800 57690
rect 106824 57638 106838 57690
rect 106838 57638 106850 57690
rect 106850 57638 106880 57690
rect 106904 57638 106914 57690
rect 106914 57638 106960 57690
rect 106664 57636 106720 57638
rect 106744 57636 106800 57638
rect 106824 57636 106880 57638
rect 106904 57636 106960 57638
rect 105928 57146 105984 57148
rect 106008 57146 106064 57148
rect 106088 57146 106144 57148
rect 106168 57146 106224 57148
rect 105928 57094 105974 57146
rect 105974 57094 105984 57146
rect 106008 57094 106038 57146
rect 106038 57094 106050 57146
rect 106050 57094 106064 57146
rect 106088 57094 106102 57146
rect 106102 57094 106114 57146
rect 106114 57094 106144 57146
rect 106168 57094 106178 57146
rect 106178 57094 106224 57146
rect 105928 57092 105984 57094
rect 106008 57092 106064 57094
rect 106088 57092 106144 57094
rect 106168 57092 106224 57094
rect 106664 56602 106720 56604
rect 106744 56602 106800 56604
rect 106824 56602 106880 56604
rect 106904 56602 106960 56604
rect 106664 56550 106710 56602
rect 106710 56550 106720 56602
rect 106744 56550 106774 56602
rect 106774 56550 106786 56602
rect 106786 56550 106800 56602
rect 106824 56550 106838 56602
rect 106838 56550 106850 56602
rect 106850 56550 106880 56602
rect 106904 56550 106914 56602
rect 106914 56550 106960 56602
rect 106664 56548 106720 56550
rect 106744 56548 106800 56550
rect 106824 56548 106880 56550
rect 106904 56548 106960 56550
rect 105928 56058 105984 56060
rect 106008 56058 106064 56060
rect 106088 56058 106144 56060
rect 106168 56058 106224 56060
rect 105928 56006 105974 56058
rect 105974 56006 105984 56058
rect 106008 56006 106038 56058
rect 106038 56006 106050 56058
rect 106050 56006 106064 56058
rect 106088 56006 106102 56058
rect 106102 56006 106114 56058
rect 106114 56006 106144 56058
rect 106168 56006 106178 56058
rect 106178 56006 106224 56058
rect 105928 56004 105984 56006
rect 106008 56004 106064 56006
rect 106088 56004 106144 56006
rect 106168 56004 106224 56006
rect 106664 55514 106720 55516
rect 106744 55514 106800 55516
rect 106824 55514 106880 55516
rect 106904 55514 106960 55516
rect 106664 55462 106710 55514
rect 106710 55462 106720 55514
rect 106744 55462 106774 55514
rect 106774 55462 106786 55514
rect 106786 55462 106800 55514
rect 106824 55462 106838 55514
rect 106838 55462 106850 55514
rect 106850 55462 106880 55514
rect 106904 55462 106914 55514
rect 106914 55462 106960 55514
rect 106664 55460 106720 55462
rect 106744 55460 106800 55462
rect 106824 55460 106880 55462
rect 106904 55460 106960 55462
rect 105928 54970 105984 54972
rect 106008 54970 106064 54972
rect 106088 54970 106144 54972
rect 106168 54970 106224 54972
rect 105928 54918 105974 54970
rect 105974 54918 105984 54970
rect 106008 54918 106038 54970
rect 106038 54918 106050 54970
rect 106050 54918 106064 54970
rect 106088 54918 106102 54970
rect 106102 54918 106114 54970
rect 106114 54918 106144 54970
rect 106168 54918 106178 54970
rect 106178 54918 106224 54970
rect 105928 54916 105984 54918
rect 106008 54916 106064 54918
rect 106088 54916 106144 54918
rect 106168 54916 106224 54918
rect 106664 54426 106720 54428
rect 106744 54426 106800 54428
rect 106824 54426 106880 54428
rect 106904 54426 106960 54428
rect 106664 54374 106710 54426
rect 106710 54374 106720 54426
rect 106744 54374 106774 54426
rect 106774 54374 106786 54426
rect 106786 54374 106800 54426
rect 106824 54374 106838 54426
rect 106838 54374 106850 54426
rect 106850 54374 106880 54426
rect 106904 54374 106914 54426
rect 106914 54374 106960 54426
rect 106664 54372 106720 54374
rect 106744 54372 106800 54374
rect 106824 54372 106880 54374
rect 106904 54372 106960 54374
rect 105928 53882 105984 53884
rect 106008 53882 106064 53884
rect 106088 53882 106144 53884
rect 106168 53882 106224 53884
rect 105928 53830 105974 53882
rect 105974 53830 105984 53882
rect 106008 53830 106038 53882
rect 106038 53830 106050 53882
rect 106050 53830 106064 53882
rect 106088 53830 106102 53882
rect 106102 53830 106114 53882
rect 106114 53830 106144 53882
rect 106168 53830 106178 53882
rect 106178 53830 106224 53882
rect 105928 53828 105984 53830
rect 106008 53828 106064 53830
rect 106088 53828 106144 53830
rect 106168 53828 106224 53830
rect 106664 53338 106720 53340
rect 106744 53338 106800 53340
rect 106824 53338 106880 53340
rect 106904 53338 106960 53340
rect 106664 53286 106710 53338
rect 106710 53286 106720 53338
rect 106744 53286 106774 53338
rect 106774 53286 106786 53338
rect 106786 53286 106800 53338
rect 106824 53286 106838 53338
rect 106838 53286 106850 53338
rect 106850 53286 106880 53338
rect 106904 53286 106914 53338
rect 106914 53286 106960 53338
rect 106664 53284 106720 53286
rect 106744 53284 106800 53286
rect 106824 53284 106880 53286
rect 106904 53284 106960 53286
rect 105928 52794 105984 52796
rect 106008 52794 106064 52796
rect 106088 52794 106144 52796
rect 106168 52794 106224 52796
rect 105928 52742 105974 52794
rect 105974 52742 105984 52794
rect 106008 52742 106038 52794
rect 106038 52742 106050 52794
rect 106050 52742 106064 52794
rect 106088 52742 106102 52794
rect 106102 52742 106114 52794
rect 106114 52742 106144 52794
rect 106168 52742 106178 52794
rect 106178 52742 106224 52794
rect 105928 52740 105984 52742
rect 106008 52740 106064 52742
rect 106088 52740 106144 52742
rect 106168 52740 106224 52742
rect 106664 52250 106720 52252
rect 106744 52250 106800 52252
rect 106824 52250 106880 52252
rect 106904 52250 106960 52252
rect 106664 52198 106710 52250
rect 106710 52198 106720 52250
rect 106744 52198 106774 52250
rect 106774 52198 106786 52250
rect 106786 52198 106800 52250
rect 106824 52198 106838 52250
rect 106838 52198 106850 52250
rect 106850 52198 106880 52250
rect 106904 52198 106914 52250
rect 106914 52198 106960 52250
rect 106664 52196 106720 52198
rect 106744 52196 106800 52198
rect 106824 52196 106880 52198
rect 106904 52196 106960 52198
rect 105928 51706 105984 51708
rect 106008 51706 106064 51708
rect 106088 51706 106144 51708
rect 106168 51706 106224 51708
rect 105928 51654 105974 51706
rect 105974 51654 105984 51706
rect 106008 51654 106038 51706
rect 106038 51654 106050 51706
rect 106050 51654 106064 51706
rect 106088 51654 106102 51706
rect 106102 51654 106114 51706
rect 106114 51654 106144 51706
rect 106168 51654 106178 51706
rect 106178 51654 106224 51706
rect 105928 51652 105984 51654
rect 106008 51652 106064 51654
rect 106088 51652 106144 51654
rect 106168 51652 106224 51654
rect 106664 51162 106720 51164
rect 106744 51162 106800 51164
rect 106824 51162 106880 51164
rect 106904 51162 106960 51164
rect 106664 51110 106710 51162
rect 106710 51110 106720 51162
rect 106744 51110 106774 51162
rect 106774 51110 106786 51162
rect 106786 51110 106800 51162
rect 106824 51110 106838 51162
rect 106838 51110 106850 51162
rect 106850 51110 106880 51162
rect 106904 51110 106914 51162
rect 106914 51110 106960 51162
rect 106664 51108 106720 51110
rect 106744 51108 106800 51110
rect 106824 51108 106880 51110
rect 106904 51108 106960 51110
rect 105928 50618 105984 50620
rect 106008 50618 106064 50620
rect 106088 50618 106144 50620
rect 106168 50618 106224 50620
rect 105928 50566 105974 50618
rect 105974 50566 105984 50618
rect 106008 50566 106038 50618
rect 106038 50566 106050 50618
rect 106050 50566 106064 50618
rect 106088 50566 106102 50618
rect 106102 50566 106114 50618
rect 106114 50566 106144 50618
rect 106168 50566 106178 50618
rect 106178 50566 106224 50618
rect 105928 50564 105984 50566
rect 106008 50564 106064 50566
rect 106088 50564 106144 50566
rect 106168 50564 106224 50566
rect 106664 50074 106720 50076
rect 106744 50074 106800 50076
rect 106824 50074 106880 50076
rect 106904 50074 106960 50076
rect 106664 50022 106710 50074
rect 106710 50022 106720 50074
rect 106744 50022 106774 50074
rect 106774 50022 106786 50074
rect 106786 50022 106800 50074
rect 106824 50022 106838 50074
rect 106838 50022 106850 50074
rect 106850 50022 106880 50074
rect 106904 50022 106914 50074
rect 106914 50022 106960 50074
rect 106664 50020 106720 50022
rect 106744 50020 106800 50022
rect 106824 50020 106880 50022
rect 106904 50020 106960 50022
rect 105928 49530 105984 49532
rect 106008 49530 106064 49532
rect 106088 49530 106144 49532
rect 106168 49530 106224 49532
rect 105928 49478 105974 49530
rect 105974 49478 105984 49530
rect 106008 49478 106038 49530
rect 106038 49478 106050 49530
rect 106050 49478 106064 49530
rect 106088 49478 106102 49530
rect 106102 49478 106114 49530
rect 106114 49478 106144 49530
rect 106168 49478 106178 49530
rect 106178 49478 106224 49530
rect 105928 49476 105984 49478
rect 106008 49476 106064 49478
rect 106088 49476 106144 49478
rect 106168 49476 106224 49478
rect 106664 48986 106720 48988
rect 106744 48986 106800 48988
rect 106824 48986 106880 48988
rect 106904 48986 106960 48988
rect 106664 48934 106710 48986
rect 106710 48934 106720 48986
rect 106744 48934 106774 48986
rect 106774 48934 106786 48986
rect 106786 48934 106800 48986
rect 106824 48934 106838 48986
rect 106838 48934 106850 48986
rect 106850 48934 106880 48986
rect 106904 48934 106914 48986
rect 106914 48934 106960 48986
rect 106664 48932 106720 48934
rect 106744 48932 106800 48934
rect 106824 48932 106880 48934
rect 106904 48932 106960 48934
rect 105928 48442 105984 48444
rect 106008 48442 106064 48444
rect 106088 48442 106144 48444
rect 106168 48442 106224 48444
rect 105928 48390 105974 48442
rect 105974 48390 105984 48442
rect 106008 48390 106038 48442
rect 106038 48390 106050 48442
rect 106050 48390 106064 48442
rect 106088 48390 106102 48442
rect 106102 48390 106114 48442
rect 106114 48390 106144 48442
rect 106168 48390 106178 48442
rect 106178 48390 106224 48442
rect 105928 48388 105984 48390
rect 106008 48388 106064 48390
rect 106088 48388 106144 48390
rect 106168 48388 106224 48390
rect 106664 47898 106720 47900
rect 106744 47898 106800 47900
rect 106824 47898 106880 47900
rect 106904 47898 106960 47900
rect 106664 47846 106710 47898
rect 106710 47846 106720 47898
rect 106744 47846 106774 47898
rect 106774 47846 106786 47898
rect 106786 47846 106800 47898
rect 106824 47846 106838 47898
rect 106838 47846 106850 47898
rect 106850 47846 106880 47898
rect 106904 47846 106914 47898
rect 106914 47846 106960 47898
rect 106664 47844 106720 47846
rect 106744 47844 106800 47846
rect 106824 47844 106880 47846
rect 106904 47844 106960 47846
rect 105928 47354 105984 47356
rect 106008 47354 106064 47356
rect 106088 47354 106144 47356
rect 106168 47354 106224 47356
rect 105928 47302 105974 47354
rect 105974 47302 105984 47354
rect 106008 47302 106038 47354
rect 106038 47302 106050 47354
rect 106050 47302 106064 47354
rect 106088 47302 106102 47354
rect 106102 47302 106114 47354
rect 106114 47302 106144 47354
rect 106168 47302 106178 47354
rect 106178 47302 106224 47354
rect 105928 47300 105984 47302
rect 106008 47300 106064 47302
rect 106088 47300 106144 47302
rect 106168 47300 106224 47302
rect 106664 46810 106720 46812
rect 106744 46810 106800 46812
rect 106824 46810 106880 46812
rect 106904 46810 106960 46812
rect 106664 46758 106710 46810
rect 106710 46758 106720 46810
rect 106744 46758 106774 46810
rect 106774 46758 106786 46810
rect 106786 46758 106800 46810
rect 106824 46758 106838 46810
rect 106838 46758 106850 46810
rect 106850 46758 106880 46810
rect 106904 46758 106914 46810
rect 106914 46758 106960 46810
rect 106664 46756 106720 46758
rect 106744 46756 106800 46758
rect 106824 46756 106880 46758
rect 106904 46756 106960 46758
rect 105928 46266 105984 46268
rect 106008 46266 106064 46268
rect 106088 46266 106144 46268
rect 106168 46266 106224 46268
rect 105928 46214 105974 46266
rect 105974 46214 105984 46266
rect 106008 46214 106038 46266
rect 106038 46214 106050 46266
rect 106050 46214 106064 46266
rect 106088 46214 106102 46266
rect 106102 46214 106114 46266
rect 106114 46214 106144 46266
rect 106168 46214 106178 46266
rect 106178 46214 106224 46266
rect 105928 46212 105984 46214
rect 106008 46212 106064 46214
rect 106088 46212 106144 46214
rect 106168 46212 106224 46214
rect 106664 45722 106720 45724
rect 106744 45722 106800 45724
rect 106824 45722 106880 45724
rect 106904 45722 106960 45724
rect 106664 45670 106710 45722
rect 106710 45670 106720 45722
rect 106744 45670 106774 45722
rect 106774 45670 106786 45722
rect 106786 45670 106800 45722
rect 106824 45670 106838 45722
rect 106838 45670 106850 45722
rect 106850 45670 106880 45722
rect 106904 45670 106914 45722
rect 106914 45670 106960 45722
rect 106664 45668 106720 45670
rect 106744 45668 106800 45670
rect 106824 45668 106880 45670
rect 106904 45668 106960 45670
rect 105928 45178 105984 45180
rect 106008 45178 106064 45180
rect 106088 45178 106144 45180
rect 106168 45178 106224 45180
rect 105928 45126 105974 45178
rect 105974 45126 105984 45178
rect 106008 45126 106038 45178
rect 106038 45126 106050 45178
rect 106050 45126 106064 45178
rect 106088 45126 106102 45178
rect 106102 45126 106114 45178
rect 106114 45126 106144 45178
rect 106168 45126 106178 45178
rect 106178 45126 106224 45178
rect 105928 45124 105984 45126
rect 106008 45124 106064 45126
rect 106088 45124 106144 45126
rect 106168 45124 106224 45126
rect 106664 44634 106720 44636
rect 106744 44634 106800 44636
rect 106824 44634 106880 44636
rect 106904 44634 106960 44636
rect 106664 44582 106710 44634
rect 106710 44582 106720 44634
rect 106744 44582 106774 44634
rect 106774 44582 106786 44634
rect 106786 44582 106800 44634
rect 106824 44582 106838 44634
rect 106838 44582 106850 44634
rect 106850 44582 106880 44634
rect 106904 44582 106914 44634
rect 106914 44582 106960 44634
rect 106664 44580 106720 44582
rect 106744 44580 106800 44582
rect 106824 44580 106880 44582
rect 106904 44580 106960 44582
rect 105928 44090 105984 44092
rect 106008 44090 106064 44092
rect 106088 44090 106144 44092
rect 106168 44090 106224 44092
rect 105928 44038 105974 44090
rect 105974 44038 105984 44090
rect 106008 44038 106038 44090
rect 106038 44038 106050 44090
rect 106050 44038 106064 44090
rect 106088 44038 106102 44090
rect 106102 44038 106114 44090
rect 106114 44038 106144 44090
rect 106168 44038 106178 44090
rect 106178 44038 106224 44090
rect 105928 44036 105984 44038
rect 106008 44036 106064 44038
rect 106088 44036 106144 44038
rect 106168 44036 106224 44038
rect 106664 43546 106720 43548
rect 106744 43546 106800 43548
rect 106824 43546 106880 43548
rect 106904 43546 106960 43548
rect 106664 43494 106710 43546
rect 106710 43494 106720 43546
rect 106744 43494 106774 43546
rect 106774 43494 106786 43546
rect 106786 43494 106800 43546
rect 106824 43494 106838 43546
rect 106838 43494 106850 43546
rect 106850 43494 106880 43546
rect 106904 43494 106914 43546
rect 106914 43494 106960 43546
rect 106664 43492 106720 43494
rect 106744 43492 106800 43494
rect 106824 43492 106880 43494
rect 106904 43492 106960 43494
rect 105928 43002 105984 43004
rect 106008 43002 106064 43004
rect 106088 43002 106144 43004
rect 106168 43002 106224 43004
rect 105928 42950 105974 43002
rect 105974 42950 105984 43002
rect 106008 42950 106038 43002
rect 106038 42950 106050 43002
rect 106050 42950 106064 43002
rect 106088 42950 106102 43002
rect 106102 42950 106114 43002
rect 106114 42950 106144 43002
rect 106168 42950 106178 43002
rect 106178 42950 106224 43002
rect 105928 42948 105984 42950
rect 106008 42948 106064 42950
rect 106088 42948 106144 42950
rect 106168 42948 106224 42950
rect 106664 42458 106720 42460
rect 106744 42458 106800 42460
rect 106824 42458 106880 42460
rect 106904 42458 106960 42460
rect 106664 42406 106710 42458
rect 106710 42406 106720 42458
rect 106744 42406 106774 42458
rect 106774 42406 106786 42458
rect 106786 42406 106800 42458
rect 106824 42406 106838 42458
rect 106838 42406 106850 42458
rect 106850 42406 106880 42458
rect 106904 42406 106914 42458
rect 106914 42406 106960 42458
rect 106664 42404 106720 42406
rect 106744 42404 106800 42406
rect 106824 42404 106880 42406
rect 106904 42404 106960 42406
rect 105928 41914 105984 41916
rect 106008 41914 106064 41916
rect 106088 41914 106144 41916
rect 106168 41914 106224 41916
rect 105928 41862 105974 41914
rect 105974 41862 105984 41914
rect 106008 41862 106038 41914
rect 106038 41862 106050 41914
rect 106050 41862 106064 41914
rect 106088 41862 106102 41914
rect 106102 41862 106114 41914
rect 106114 41862 106144 41914
rect 106168 41862 106178 41914
rect 106178 41862 106224 41914
rect 105928 41860 105984 41862
rect 106008 41860 106064 41862
rect 106088 41860 106144 41862
rect 106168 41860 106224 41862
rect 106664 41370 106720 41372
rect 106744 41370 106800 41372
rect 106824 41370 106880 41372
rect 106904 41370 106960 41372
rect 106664 41318 106710 41370
rect 106710 41318 106720 41370
rect 106744 41318 106774 41370
rect 106774 41318 106786 41370
rect 106786 41318 106800 41370
rect 106824 41318 106838 41370
rect 106838 41318 106850 41370
rect 106850 41318 106880 41370
rect 106904 41318 106914 41370
rect 106914 41318 106960 41370
rect 106664 41316 106720 41318
rect 106744 41316 106800 41318
rect 106824 41316 106880 41318
rect 106904 41316 106960 41318
rect 105928 40826 105984 40828
rect 106008 40826 106064 40828
rect 106088 40826 106144 40828
rect 106168 40826 106224 40828
rect 105928 40774 105974 40826
rect 105974 40774 105984 40826
rect 106008 40774 106038 40826
rect 106038 40774 106050 40826
rect 106050 40774 106064 40826
rect 106088 40774 106102 40826
rect 106102 40774 106114 40826
rect 106114 40774 106144 40826
rect 106168 40774 106178 40826
rect 106178 40774 106224 40826
rect 105928 40772 105984 40774
rect 106008 40772 106064 40774
rect 106088 40772 106144 40774
rect 106168 40772 106224 40774
rect 106664 40282 106720 40284
rect 106744 40282 106800 40284
rect 106824 40282 106880 40284
rect 106904 40282 106960 40284
rect 106664 40230 106710 40282
rect 106710 40230 106720 40282
rect 106744 40230 106774 40282
rect 106774 40230 106786 40282
rect 106786 40230 106800 40282
rect 106824 40230 106838 40282
rect 106838 40230 106850 40282
rect 106850 40230 106880 40282
rect 106904 40230 106914 40282
rect 106914 40230 106960 40282
rect 106664 40228 106720 40230
rect 106744 40228 106800 40230
rect 106824 40228 106880 40230
rect 106904 40228 106960 40230
rect 105928 39738 105984 39740
rect 106008 39738 106064 39740
rect 106088 39738 106144 39740
rect 106168 39738 106224 39740
rect 105928 39686 105974 39738
rect 105974 39686 105984 39738
rect 106008 39686 106038 39738
rect 106038 39686 106050 39738
rect 106050 39686 106064 39738
rect 106088 39686 106102 39738
rect 106102 39686 106114 39738
rect 106114 39686 106144 39738
rect 106168 39686 106178 39738
rect 106178 39686 106224 39738
rect 105928 39684 105984 39686
rect 106008 39684 106064 39686
rect 106088 39684 106144 39686
rect 106168 39684 106224 39686
rect 106664 39194 106720 39196
rect 106744 39194 106800 39196
rect 106824 39194 106880 39196
rect 106904 39194 106960 39196
rect 106664 39142 106710 39194
rect 106710 39142 106720 39194
rect 106744 39142 106774 39194
rect 106774 39142 106786 39194
rect 106786 39142 106800 39194
rect 106824 39142 106838 39194
rect 106838 39142 106850 39194
rect 106850 39142 106880 39194
rect 106904 39142 106914 39194
rect 106914 39142 106960 39194
rect 106664 39140 106720 39142
rect 106744 39140 106800 39142
rect 106824 39140 106880 39142
rect 106904 39140 106960 39142
rect 105928 38650 105984 38652
rect 106008 38650 106064 38652
rect 106088 38650 106144 38652
rect 106168 38650 106224 38652
rect 105928 38598 105974 38650
rect 105974 38598 105984 38650
rect 106008 38598 106038 38650
rect 106038 38598 106050 38650
rect 106050 38598 106064 38650
rect 106088 38598 106102 38650
rect 106102 38598 106114 38650
rect 106114 38598 106144 38650
rect 106168 38598 106178 38650
rect 106178 38598 106224 38650
rect 105928 38596 105984 38598
rect 106008 38596 106064 38598
rect 106088 38596 106144 38598
rect 106168 38596 106224 38598
rect 106664 38106 106720 38108
rect 106744 38106 106800 38108
rect 106824 38106 106880 38108
rect 106904 38106 106960 38108
rect 106664 38054 106710 38106
rect 106710 38054 106720 38106
rect 106744 38054 106774 38106
rect 106774 38054 106786 38106
rect 106786 38054 106800 38106
rect 106824 38054 106838 38106
rect 106838 38054 106850 38106
rect 106850 38054 106880 38106
rect 106904 38054 106914 38106
rect 106914 38054 106960 38106
rect 106664 38052 106720 38054
rect 106744 38052 106800 38054
rect 106824 38052 106880 38054
rect 106904 38052 106960 38054
rect 105928 37562 105984 37564
rect 106008 37562 106064 37564
rect 106088 37562 106144 37564
rect 106168 37562 106224 37564
rect 105928 37510 105974 37562
rect 105974 37510 105984 37562
rect 106008 37510 106038 37562
rect 106038 37510 106050 37562
rect 106050 37510 106064 37562
rect 106088 37510 106102 37562
rect 106102 37510 106114 37562
rect 106114 37510 106144 37562
rect 106168 37510 106178 37562
rect 106178 37510 106224 37562
rect 105928 37508 105984 37510
rect 106008 37508 106064 37510
rect 106088 37508 106144 37510
rect 106168 37508 106224 37510
rect 106664 37018 106720 37020
rect 106744 37018 106800 37020
rect 106824 37018 106880 37020
rect 106904 37018 106960 37020
rect 106664 36966 106710 37018
rect 106710 36966 106720 37018
rect 106744 36966 106774 37018
rect 106774 36966 106786 37018
rect 106786 36966 106800 37018
rect 106824 36966 106838 37018
rect 106838 36966 106850 37018
rect 106850 36966 106880 37018
rect 106904 36966 106914 37018
rect 106914 36966 106960 37018
rect 106664 36964 106720 36966
rect 106744 36964 106800 36966
rect 106824 36964 106880 36966
rect 106904 36964 106960 36966
rect 105928 36474 105984 36476
rect 106008 36474 106064 36476
rect 106088 36474 106144 36476
rect 106168 36474 106224 36476
rect 105928 36422 105974 36474
rect 105974 36422 105984 36474
rect 106008 36422 106038 36474
rect 106038 36422 106050 36474
rect 106050 36422 106064 36474
rect 106088 36422 106102 36474
rect 106102 36422 106114 36474
rect 106114 36422 106144 36474
rect 106168 36422 106178 36474
rect 106178 36422 106224 36474
rect 105928 36420 105984 36422
rect 106008 36420 106064 36422
rect 106088 36420 106144 36422
rect 106168 36420 106224 36422
rect 106664 35930 106720 35932
rect 106744 35930 106800 35932
rect 106824 35930 106880 35932
rect 106904 35930 106960 35932
rect 106664 35878 106710 35930
rect 106710 35878 106720 35930
rect 106744 35878 106774 35930
rect 106774 35878 106786 35930
rect 106786 35878 106800 35930
rect 106824 35878 106838 35930
rect 106838 35878 106850 35930
rect 106850 35878 106880 35930
rect 106904 35878 106914 35930
rect 106914 35878 106960 35930
rect 106664 35876 106720 35878
rect 106744 35876 106800 35878
rect 106824 35876 106880 35878
rect 106904 35876 106960 35878
rect 105928 35386 105984 35388
rect 106008 35386 106064 35388
rect 106088 35386 106144 35388
rect 106168 35386 106224 35388
rect 105928 35334 105974 35386
rect 105974 35334 105984 35386
rect 106008 35334 106038 35386
rect 106038 35334 106050 35386
rect 106050 35334 106064 35386
rect 106088 35334 106102 35386
rect 106102 35334 106114 35386
rect 106114 35334 106144 35386
rect 106168 35334 106178 35386
rect 106178 35334 106224 35386
rect 105928 35332 105984 35334
rect 106008 35332 106064 35334
rect 106088 35332 106144 35334
rect 106168 35332 106224 35334
rect 106664 34842 106720 34844
rect 106744 34842 106800 34844
rect 106824 34842 106880 34844
rect 106904 34842 106960 34844
rect 106664 34790 106710 34842
rect 106710 34790 106720 34842
rect 106744 34790 106774 34842
rect 106774 34790 106786 34842
rect 106786 34790 106800 34842
rect 106824 34790 106838 34842
rect 106838 34790 106850 34842
rect 106850 34790 106880 34842
rect 106904 34790 106914 34842
rect 106914 34790 106960 34842
rect 106664 34788 106720 34790
rect 106744 34788 106800 34790
rect 106824 34788 106880 34790
rect 106904 34788 106960 34790
rect 105928 34298 105984 34300
rect 106008 34298 106064 34300
rect 106088 34298 106144 34300
rect 106168 34298 106224 34300
rect 105928 34246 105974 34298
rect 105974 34246 105984 34298
rect 106008 34246 106038 34298
rect 106038 34246 106050 34298
rect 106050 34246 106064 34298
rect 106088 34246 106102 34298
rect 106102 34246 106114 34298
rect 106114 34246 106144 34298
rect 106168 34246 106178 34298
rect 106178 34246 106224 34298
rect 105928 34244 105984 34246
rect 106008 34244 106064 34246
rect 106088 34244 106144 34246
rect 106168 34244 106224 34246
rect 106664 33754 106720 33756
rect 106744 33754 106800 33756
rect 106824 33754 106880 33756
rect 106904 33754 106960 33756
rect 106664 33702 106710 33754
rect 106710 33702 106720 33754
rect 106744 33702 106774 33754
rect 106774 33702 106786 33754
rect 106786 33702 106800 33754
rect 106824 33702 106838 33754
rect 106838 33702 106850 33754
rect 106850 33702 106880 33754
rect 106904 33702 106914 33754
rect 106914 33702 106960 33754
rect 106664 33700 106720 33702
rect 106744 33700 106800 33702
rect 106824 33700 106880 33702
rect 106904 33700 106960 33702
rect 105928 33210 105984 33212
rect 106008 33210 106064 33212
rect 106088 33210 106144 33212
rect 106168 33210 106224 33212
rect 105928 33158 105974 33210
rect 105974 33158 105984 33210
rect 106008 33158 106038 33210
rect 106038 33158 106050 33210
rect 106050 33158 106064 33210
rect 106088 33158 106102 33210
rect 106102 33158 106114 33210
rect 106114 33158 106144 33210
rect 106168 33158 106178 33210
rect 106178 33158 106224 33210
rect 105928 33156 105984 33158
rect 106008 33156 106064 33158
rect 106088 33156 106144 33158
rect 106168 33156 106224 33158
rect 106664 32666 106720 32668
rect 106744 32666 106800 32668
rect 106824 32666 106880 32668
rect 106904 32666 106960 32668
rect 106664 32614 106710 32666
rect 106710 32614 106720 32666
rect 106744 32614 106774 32666
rect 106774 32614 106786 32666
rect 106786 32614 106800 32666
rect 106824 32614 106838 32666
rect 106838 32614 106850 32666
rect 106850 32614 106880 32666
rect 106904 32614 106914 32666
rect 106914 32614 106960 32666
rect 106664 32612 106720 32614
rect 106744 32612 106800 32614
rect 106824 32612 106880 32614
rect 106904 32612 106960 32614
rect 105928 32122 105984 32124
rect 106008 32122 106064 32124
rect 106088 32122 106144 32124
rect 106168 32122 106224 32124
rect 105928 32070 105974 32122
rect 105974 32070 105984 32122
rect 106008 32070 106038 32122
rect 106038 32070 106050 32122
rect 106050 32070 106064 32122
rect 106088 32070 106102 32122
rect 106102 32070 106114 32122
rect 106114 32070 106144 32122
rect 106168 32070 106178 32122
rect 106178 32070 106224 32122
rect 105928 32068 105984 32070
rect 106008 32068 106064 32070
rect 106088 32068 106144 32070
rect 106168 32068 106224 32070
rect 106664 31578 106720 31580
rect 106744 31578 106800 31580
rect 106824 31578 106880 31580
rect 106904 31578 106960 31580
rect 106664 31526 106710 31578
rect 106710 31526 106720 31578
rect 106744 31526 106774 31578
rect 106774 31526 106786 31578
rect 106786 31526 106800 31578
rect 106824 31526 106838 31578
rect 106838 31526 106850 31578
rect 106850 31526 106880 31578
rect 106904 31526 106914 31578
rect 106914 31526 106960 31578
rect 106664 31524 106720 31526
rect 106744 31524 106800 31526
rect 106824 31524 106880 31526
rect 106904 31524 106960 31526
rect 105928 31034 105984 31036
rect 106008 31034 106064 31036
rect 106088 31034 106144 31036
rect 106168 31034 106224 31036
rect 105928 30982 105974 31034
rect 105974 30982 105984 31034
rect 106008 30982 106038 31034
rect 106038 30982 106050 31034
rect 106050 30982 106064 31034
rect 106088 30982 106102 31034
rect 106102 30982 106114 31034
rect 106114 30982 106144 31034
rect 106168 30982 106178 31034
rect 106178 30982 106224 31034
rect 105928 30980 105984 30982
rect 106008 30980 106064 30982
rect 106088 30980 106144 30982
rect 106168 30980 106224 30982
rect 106664 30490 106720 30492
rect 106744 30490 106800 30492
rect 106824 30490 106880 30492
rect 106904 30490 106960 30492
rect 106664 30438 106710 30490
rect 106710 30438 106720 30490
rect 106744 30438 106774 30490
rect 106774 30438 106786 30490
rect 106786 30438 106800 30490
rect 106824 30438 106838 30490
rect 106838 30438 106850 30490
rect 106850 30438 106880 30490
rect 106904 30438 106914 30490
rect 106914 30438 106960 30490
rect 106664 30436 106720 30438
rect 106744 30436 106800 30438
rect 106824 30436 106880 30438
rect 106904 30436 106960 30438
rect 105928 29946 105984 29948
rect 106008 29946 106064 29948
rect 106088 29946 106144 29948
rect 106168 29946 106224 29948
rect 105928 29894 105974 29946
rect 105974 29894 105984 29946
rect 106008 29894 106038 29946
rect 106038 29894 106050 29946
rect 106050 29894 106064 29946
rect 106088 29894 106102 29946
rect 106102 29894 106114 29946
rect 106114 29894 106144 29946
rect 106168 29894 106178 29946
rect 106178 29894 106224 29946
rect 105928 29892 105984 29894
rect 106008 29892 106064 29894
rect 106088 29892 106144 29894
rect 106168 29892 106224 29894
rect 106664 29402 106720 29404
rect 106744 29402 106800 29404
rect 106824 29402 106880 29404
rect 106904 29402 106960 29404
rect 106664 29350 106710 29402
rect 106710 29350 106720 29402
rect 106744 29350 106774 29402
rect 106774 29350 106786 29402
rect 106786 29350 106800 29402
rect 106824 29350 106838 29402
rect 106838 29350 106850 29402
rect 106850 29350 106880 29402
rect 106904 29350 106914 29402
rect 106914 29350 106960 29402
rect 106664 29348 106720 29350
rect 106744 29348 106800 29350
rect 106824 29348 106880 29350
rect 106904 29348 106960 29350
rect 105928 28858 105984 28860
rect 106008 28858 106064 28860
rect 106088 28858 106144 28860
rect 106168 28858 106224 28860
rect 105928 28806 105974 28858
rect 105974 28806 105984 28858
rect 106008 28806 106038 28858
rect 106038 28806 106050 28858
rect 106050 28806 106064 28858
rect 106088 28806 106102 28858
rect 106102 28806 106114 28858
rect 106114 28806 106144 28858
rect 106168 28806 106178 28858
rect 106178 28806 106224 28858
rect 105928 28804 105984 28806
rect 106008 28804 106064 28806
rect 106088 28804 106144 28806
rect 106168 28804 106224 28806
rect 106664 28314 106720 28316
rect 106744 28314 106800 28316
rect 106824 28314 106880 28316
rect 106904 28314 106960 28316
rect 106664 28262 106710 28314
rect 106710 28262 106720 28314
rect 106744 28262 106774 28314
rect 106774 28262 106786 28314
rect 106786 28262 106800 28314
rect 106824 28262 106838 28314
rect 106838 28262 106850 28314
rect 106850 28262 106880 28314
rect 106904 28262 106914 28314
rect 106914 28262 106960 28314
rect 106664 28260 106720 28262
rect 106744 28260 106800 28262
rect 106824 28260 106880 28262
rect 106904 28260 106960 28262
rect 105928 27770 105984 27772
rect 106008 27770 106064 27772
rect 106088 27770 106144 27772
rect 106168 27770 106224 27772
rect 105928 27718 105974 27770
rect 105974 27718 105984 27770
rect 106008 27718 106038 27770
rect 106038 27718 106050 27770
rect 106050 27718 106064 27770
rect 106088 27718 106102 27770
rect 106102 27718 106114 27770
rect 106114 27718 106144 27770
rect 106168 27718 106178 27770
rect 106178 27718 106224 27770
rect 105928 27716 105984 27718
rect 106008 27716 106064 27718
rect 106088 27716 106144 27718
rect 106168 27716 106224 27718
rect 106664 27226 106720 27228
rect 106744 27226 106800 27228
rect 106824 27226 106880 27228
rect 106904 27226 106960 27228
rect 106664 27174 106710 27226
rect 106710 27174 106720 27226
rect 106744 27174 106774 27226
rect 106774 27174 106786 27226
rect 106786 27174 106800 27226
rect 106824 27174 106838 27226
rect 106838 27174 106850 27226
rect 106850 27174 106880 27226
rect 106904 27174 106914 27226
rect 106914 27174 106960 27226
rect 106664 27172 106720 27174
rect 106744 27172 106800 27174
rect 106824 27172 106880 27174
rect 106904 27172 106960 27174
rect 105928 26682 105984 26684
rect 106008 26682 106064 26684
rect 106088 26682 106144 26684
rect 106168 26682 106224 26684
rect 105928 26630 105974 26682
rect 105974 26630 105984 26682
rect 106008 26630 106038 26682
rect 106038 26630 106050 26682
rect 106050 26630 106064 26682
rect 106088 26630 106102 26682
rect 106102 26630 106114 26682
rect 106114 26630 106144 26682
rect 106168 26630 106178 26682
rect 106178 26630 106224 26682
rect 105928 26628 105984 26630
rect 106008 26628 106064 26630
rect 106088 26628 106144 26630
rect 106168 26628 106224 26630
rect 106664 26138 106720 26140
rect 106744 26138 106800 26140
rect 106824 26138 106880 26140
rect 106904 26138 106960 26140
rect 106664 26086 106710 26138
rect 106710 26086 106720 26138
rect 106744 26086 106774 26138
rect 106774 26086 106786 26138
rect 106786 26086 106800 26138
rect 106824 26086 106838 26138
rect 106838 26086 106850 26138
rect 106850 26086 106880 26138
rect 106904 26086 106914 26138
rect 106914 26086 106960 26138
rect 106664 26084 106720 26086
rect 106744 26084 106800 26086
rect 106824 26084 106880 26086
rect 106904 26084 106960 26086
rect 105928 25594 105984 25596
rect 106008 25594 106064 25596
rect 106088 25594 106144 25596
rect 106168 25594 106224 25596
rect 105928 25542 105974 25594
rect 105974 25542 105984 25594
rect 106008 25542 106038 25594
rect 106038 25542 106050 25594
rect 106050 25542 106064 25594
rect 106088 25542 106102 25594
rect 106102 25542 106114 25594
rect 106114 25542 106144 25594
rect 106168 25542 106178 25594
rect 106178 25542 106224 25594
rect 105928 25540 105984 25542
rect 106008 25540 106064 25542
rect 106088 25540 106144 25542
rect 106168 25540 106224 25542
rect 106664 25050 106720 25052
rect 106744 25050 106800 25052
rect 106824 25050 106880 25052
rect 106904 25050 106960 25052
rect 106664 24998 106710 25050
rect 106710 24998 106720 25050
rect 106744 24998 106774 25050
rect 106774 24998 106786 25050
rect 106786 24998 106800 25050
rect 106824 24998 106838 25050
rect 106838 24998 106850 25050
rect 106850 24998 106880 25050
rect 106904 24998 106914 25050
rect 106914 24998 106960 25050
rect 106664 24996 106720 24998
rect 106744 24996 106800 24998
rect 106824 24996 106880 24998
rect 106904 24996 106960 24998
rect 105928 24506 105984 24508
rect 106008 24506 106064 24508
rect 106088 24506 106144 24508
rect 106168 24506 106224 24508
rect 105928 24454 105974 24506
rect 105974 24454 105984 24506
rect 106008 24454 106038 24506
rect 106038 24454 106050 24506
rect 106050 24454 106064 24506
rect 106088 24454 106102 24506
rect 106102 24454 106114 24506
rect 106114 24454 106144 24506
rect 106168 24454 106178 24506
rect 106178 24454 106224 24506
rect 105928 24452 105984 24454
rect 106008 24452 106064 24454
rect 106088 24452 106144 24454
rect 106168 24452 106224 24454
rect 106664 23962 106720 23964
rect 106744 23962 106800 23964
rect 106824 23962 106880 23964
rect 106904 23962 106960 23964
rect 106664 23910 106710 23962
rect 106710 23910 106720 23962
rect 106744 23910 106774 23962
rect 106774 23910 106786 23962
rect 106786 23910 106800 23962
rect 106824 23910 106838 23962
rect 106838 23910 106850 23962
rect 106850 23910 106880 23962
rect 106904 23910 106914 23962
rect 106914 23910 106960 23962
rect 106664 23908 106720 23910
rect 106744 23908 106800 23910
rect 106824 23908 106880 23910
rect 106904 23908 106960 23910
rect 105928 23418 105984 23420
rect 106008 23418 106064 23420
rect 106088 23418 106144 23420
rect 106168 23418 106224 23420
rect 105928 23366 105974 23418
rect 105974 23366 105984 23418
rect 106008 23366 106038 23418
rect 106038 23366 106050 23418
rect 106050 23366 106064 23418
rect 106088 23366 106102 23418
rect 106102 23366 106114 23418
rect 106114 23366 106144 23418
rect 106168 23366 106178 23418
rect 106178 23366 106224 23418
rect 105928 23364 105984 23366
rect 106008 23364 106064 23366
rect 106088 23364 106144 23366
rect 106168 23364 106224 23366
rect 106664 22874 106720 22876
rect 106744 22874 106800 22876
rect 106824 22874 106880 22876
rect 106904 22874 106960 22876
rect 106664 22822 106710 22874
rect 106710 22822 106720 22874
rect 106744 22822 106774 22874
rect 106774 22822 106786 22874
rect 106786 22822 106800 22874
rect 106824 22822 106838 22874
rect 106838 22822 106850 22874
rect 106850 22822 106880 22874
rect 106904 22822 106914 22874
rect 106914 22822 106960 22874
rect 106664 22820 106720 22822
rect 106744 22820 106800 22822
rect 106824 22820 106880 22822
rect 106904 22820 106960 22822
rect 105928 22330 105984 22332
rect 106008 22330 106064 22332
rect 106088 22330 106144 22332
rect 106168 22330 106224 22332
rect 105928 22278 105974 22330
rect 105974 22278 105984 22330
rect 106008 22278 106038 22330
rect 106038 22278 106050 22330
rect 106050 22278 106064 22330
rect 106088 22278 106102 22330
rect 106102 22278 106114 22330
rect 106114 22278 106144 22330
rect 106168 22278 106178 22330
rect 106178 22278 106224 22330
rect 105928 22276 105984 22278
rect 106008 22276 106064 22278
rect 106088 22276 106144 22278
rect 106168 22276 106224 22278
rect 106664 21786 106720 21788
rect 106744 21786 106800 21788
rect 106824 21786 106880 21788
rect 106904 21786 106960 21788
rect 106664 21734 106710 21786
rect 106710 21734 106720 21786
rect 106744 21734 106774 21786
rect 106774 21734 106786 21786
rect 106786 21734 106800 21786
rect 106824 21734 106838 21786
rect 106838 21734 106850 21786
rect 106850 21734 106880 21786
rect 106904 21734 106914 21786
rect 106914 21734 106960 21786
rect 106664 21732 106720 21734
rect 106744 21732 106800 21734
rect 106824 21732 106880 21734
rect 106904 21732 106960 21734
rect 105928 21242 105984 21244
rect 106008 21242 106064 21244
rect 106088 21242 106144 21244
rect 106168 21242 106224 21244
rect 105928 21190 105974 21242
rect 105974 21190 105984 21242
rect 106008 21190 106038 21242
rect 106038 21190 106050 21242
rect 106050 21190 106064 21242
rect 106088 21190 106102 21242
rect 106102 21190 106114 21242
rect 106114 21190 106144 21242
rect 106168 21190 106178 21242
rect 106178 21190 106224 21242
rect 105928 21188 105984 21190
rect 106008 21188 106064 21190
rect 106088 21188 106144 21190
rect 106168 21188 106224 21190
rect 106664 20698 106720 20700
rect 106744 20698 106800 20700
rect 106824 20698 106880 20700
rect 106904 20698 106960 20700
rect 106664 20646 106710 20698
rect 106710 20646 106720 20698
rect 106744 20646 106774 20698
rect 106774 20646 106786 20698
rect 106786 20646 106800 20698
rect 106824 20646 106838 20698
rect 106838 20646 106850 20698
rect 106850 20646 106880 20698
rect 106904 20646 106914 20698
rect 106914 20646 106960 20698
rect 106664 20644 106720 20646
rect 106744 20644 106800 20646
rect 106824 20644 106880 20646
rect 106904 20644 106960 20646
rect 105928 20154 105984 20156
rect 106008 20154 106064 20156
rect 106088 20154 106144 20156
rect 106168 20154 106224 20156
rect 105928 20102 105974 20154
rect 105974 20102 105984 20154
rect 106008 20102 106038 20154
rect 106038 20102 106050 20154
rect 106050 20102 106064 20154
rect 106088 20102 106102 20154
rect 106102 20102 106114 20154
rect 106114 20102 106144 20154
rect 106168 20102 106178 20154
rect 106178 20102 106224 20154
rect 105928 20100 105984 20102
rect 106008 20100 106064 20102
rect 106088 20100 106144 20102
rect 106168 20100 106224 20102
rect 106664 19610 106720 19612
rect 106744 19610 106800 19612
rect 106824 19610 106880 19612
rect 106904 19610 106960 19612
rect 106664 19558 106710 19610
rect 106710 19558 106720 19610
rect 106744 19558 106774 19610
rect 106774 19558 106786 19610
rect 106786 19558 106800 19610
rect 106824 19558 106838 19610
rect 106838 19558 106850 19610
rect 106850 19558 106880 19610
rect 106904 19558 106914 19610
rect 106914 19558 106960 19610
rect 106664 19556 106720 19558
rect 106744 19556 106800 19558
rect 106824 19556 106880 19558
rect 106904 19556 106960 19558
rect 105928 19066 105984 19068
rect 106008 19066 106064 19068
rect 106088 19066 106144 19068
rect 106168 19066 106224 19068
rect 105928 19014 105974 19066
rect 105974 19014 105984 19066
rect 106008 19014 106038 19066
rect 106038 19014 106050 19066
rect 106050 19014 106064 19066
rect 106088 19014 106102 19066
rect 106102 19014 106114 19066
rect 106114 19014 106144 19066
rect 106168 19014 106178 19066
rect 106178 19014 106224 19066
rect 105928 19012 105984 19014
rect 106008 19012 106064 19014
rect 106088 19012 106144 19014
rect 106168 19012 106224 19014
rect 106664 18522 106720 18524
rect 106744 18522 106800 18524
rect 106824 18522 106880 18524
rect 106904 18522 106960 18524
rect 106664 18470 106710 18522
rect 106710 18470 106720 18522
rect 106744 18470 106774 18522
rect 106774 18470 106786 18522
rect 106786 18470 106800 18522
rect 106824 18470 106838 18522
rect 106838 18470 106850 18522
rect 106850 18470 106880 18522
rect 106904 18470 106914 18522
rect 106914 18470 106960 18522
rect 106664 18468 106720 18470
rect 106744 18468 106800 18470
rect 106824 18468 106880 18470
rect 106904 18468 106960 18470
rect 105928 17978 105984 17980
rect 106008 17978 106064 17980
rect 106088 17978 106144 17980
rect 106168 17978 106224 17980
rect 105928 17926 105974 17978
rect 105974 17926 105984 17978
rect 106008 17926 106038 17978
rect 106038 17926 106050 17978
rect 106050 17926 106064 17978
rect 106088 17926 106102 17978
rect 106102 17926 106114 17978
rect 106114 17926 106144 17978
rect 106168 17926 106178 17978
rect 106178 17926 106224 17978
rect 105928 17924 105984 17926
rect 106008 17924 106064 17926
rect 106088 17924 106144 17926
rect 106168 17924 106224 17926
rect 106664 17434 106720 17436
rect 106744 17434 106800 17436
rect 106824 17434 106880 17436
rect 106904 17434 106960 17436
rect 106664 17382 106710 17434
rect 106710 17382 106720 17434
rect 106744 17382 106774 17434
rect 106774 17382 106786 17434
rect 106786 17382 106800 17434
rect 106824 17382 106838 17434
rect 106838 17382 106850 17434
rect 106850 17382 106880 17434
rect 106904 17382 106914 17434
rect 106914 17382 106960 17434
rect 106664 17380 106720 17382
rect 106744 17380 106800 17382
rect 106824 17380 106880 17382
rect 106904 17380 106960 17382
rect 105928 16890 105984 16892
rect 106008 16890 106064 16892
rect 106088 16890 106144 16892
rect 106168 16890 106224 16892
rect 105928 16838 105974 16890
rect 105974 16838 105984 16890
rect 106008 16838 106038 16890
rect 106038 16838 106050 16890
rect 106050 16838 106064 16890
rect 106088 16838 106102 16890
rect 106102 16838 106114 16890
rect 106114 16838 106144 16890
rect 106168 16838 106178 16890
rect 106178 16838 106224 16890
rect 105928 16836 105984 16838
rect 106008 16836 106064 16838
rect 106088 16836 106144 16838
rect 106168 16836 106224 16838
rect 106664 16346 106720 16348
rect 106744 16346 106800 16348
rect 106824 16346 106880 16348
rect 106904 16346 106960 16348
rect 106664 16294 106710 16346
rect 106710 16294 106720 16346
rect 106744 16294 106774 16346
rect 106774 16294 106786 16346
rect 106786 16294 106800 16346
rect 106824 16294 106838 16346
rect 106838 16294 106850 16346
rect 106850 16294 106880 16346
rect 106904 16294 106914 16346
rect 106914 16294 106960 16346
rect 106664 16292 106720 16294
rect 106744 16292 106800 16294
rect 106824 16292 106880 16294
rect 106904 16292 106960 16294
rect 105928 15802 105984 15804
rect 106008 15802 106064 15804
rect 106088 15802 106144 15804
rect 106168 15802 106224 15804
rect 105928 15750 105974 15802
rect 105974 15750 105984 15802
rect 106008 15750 106038 15802
rect 106038 15750 106050 15802
rect 106050 15750 106064 15802
rect 106088 15750 106102 15802
rect 106102 15750 106114 15802
rect 106114 15750 106144 15802
rect 106168 15750 106178 15802
rect 106178 15750 106224 15802
rect 105928 15748 105984 15750
rect 106008 15748 106064 15750
rect 106088 15748 106144 15750
rect 106168 15748 106224 15750
rect 106664 15258 106720 15260
rect 106744 15258 106800 15260
rect 106824 15258 106880 15260
rect 106904 15258 106960 15260
rect 106664 15206 106710 15258
rect 106710 15206 106720 15258
rect 106744 15206 106774 15258
rect 106774 15206 106786 15258
rect 106786 15206 106800 15258
rect 106824 15206 106838 15258
rect 106838 15206 106850 15258
rect 106850 15206 106880 15258
rect 106904 15206 106914 15258
rect 106914 15206 106960 15258
rect 106664 15204 106720 15206
rect 106744 15204 106800 15206
rect 106824 15204 106880 15206
rect 106904 15204 106960 15206
rect 105928 14714 105984 14716
rect 106008 14714 106064 14716
rect 106088 14714 106144 14716
rect 106168 14714 106224 14716
rect 105928 14662 105974 14714
rect 105974 14662 105984 14714
rect 106008 14662 106038 14714
rect 106038 14662 106050 14714
rect 106050 14662 106064 14714
rect 106088 14662 106102 14714
rect 106102 14662 106114 14714
rect 106114 14662 106144 14714
rect 106168 14662 106178 14714
rect 106178 14662 106224 14714
rect 105928 14660 105984 14662
rect 106008 14660 106064 14662
rect 106088 14660 106144 14662
rect 106168 14660 106224 14662
rect 106664 14170 106720 14172
rect 106744 14170 106800 14172
rect 106824 14170 106880 14172
rect 106904 14170 106960 14172
rect 106664 14118 106710 14170
rect 106710 14118 106720 14170
rect 106744 14118 106774 14170
rect 106774 14118 106786 14170
rect 106786 14118 106800 14170
rect 106824 14118 106838 14170
rect 106838 14118 106850 14170
rect 106850 14118 106880 14170
rect 106904 14118 106914 14170
rect 106914 14118 106960 14170
rect 106664 14116 106720 14118
rect 106744 14116 106800 14118
rect 106824 14116 106880 14118
rect 106904 14116 106960 14118
rect 105928 13626 105984 13628
rect 106008 13626 106064 13628
rect 106088 13626 106144 13628
rect 106168 13626 106224 13628
rect 105928 13574 105974 13626
rect 105974 13574 105984 13626
rect 106008 13574 106038 13626
rect 106038 13574 106050 13626
rect 106050 13574 106064 13626
rect 106088 13574 106102 13626
rect 106102 13574 106114 13626
rect 106114 13574 106144 13626
rect 106168 13574 106178 13626
rect 106178 13574 106224 13626
rect 105928 13572 105984 13574
rect 106008 13572 106064 13574
rect 106088 13572 106144 13574
rect 106168 13572 106224 13574
rect 106664 13082 106720 13084
rect 106744 13082 106800 13084
rect 106824 13082 106880 13084
rect 106904 13082 106960 13084
rect 106664 13030 106710 13082
rect 106710 13030 106720 13082
rect 106744 13030 106774 13082
rect 106774 13030 106786 13082
rect 106786 13030 106800 13082
rect 106824 13030 106838 13082
rect 106838 13030 106850 13082
rect 106850 13030 106880 13082
rect 106904 13030 106914 13082
rect 106914 13030 106960 13082
rect 106664 13028 106720 13030
rect 106744 13028 106800 13030
rect 106824 13028 106880 13030
rect 106904 13028 106960 13030
rect 105928 12538 105984 12540
rect 106008 12538 106064 12540
rect 106088 12538 106144 12540
rect 106168 12538 106224 12540
rect 105928 12486 105974 12538
rect 105974 12486 105984 12538
rect 106008 12486 106038 12538
rect 106038 12486 106050 12538
rect 106050 12486 106064 12538
rect 106088 12486 106102 12538
rect 106102 12486 106114 12538
rect 106114 12486 106144 12538
rect 106168 12486 106178 12538
rect 106178 12486 106224 12538
rect 105928 12484 105984 12486
rect 106008 12484 106064 12486
rect 106088 12484 106144 12486
rect 106168 12484 106224 12486
rect 106664 11994 106720 11996
rect 106744 11994 106800 11996
rect 106824 11994 106880 11996
rect 106904 11994 106960 11996
rect 106664 11942 106710 11994
rect 106710 11942 106720 11994
rect 106744 11942 106774 11994
rect 106774 11942 106786 11994
rect 106786 11942 106800 11994
rect 106824 11942 106838 11994
rect 106838 11942 106850 11994
rect 106850 11942 106880 11994
rect 106904 11942 106914 11994
rect 106914 11942 106960 11994
rect 106664 11940 106720 11942
rect 106744 11940 106800 11942
rect 106824 11940 106880 11942
rect 106904 11940 106960 11942
rect 105928 11450 105984 11452
rect 106008 11450 106064 11452
rect 106088 11450 106144 11452
rect 106168 11450 106224 11452
rect 105928 11398 105974 11450
rect 105974 11398 105984 11450
rect 106008 11398 106038 11450
rect 106038 11398 106050 11450
rect 106050 11398 106064 11450
rect 106088 11398 106102 11450
rect 106102 11398 106114 11450
rect 106114 11398 106144 11450
rect 106168 11398 106178 11450
rect 106178 11398 106224 11450
rect 105928 11396 105984 11398
rect 106008 11396 106064 11398
rect 106088 11396 106144 11398
rect 106168 11396 106224 11398
rect 106664 10906 106720 10908
rect 106744 10906 106800 10908
rect 106824 10906 106880 10908
rect 106904 10906 106960 10908
rect 106664 10854 106710 10906
rect 106710 10854 106720 10906
rect 106744 10854 106774 10906
rect 106774 10854 106786 10906
rect 106786 10854 106800 10906
rect 106824 10854 106838 10906
rect 106838 10854 106850 10906
rect 106850 10854 106880 10906
rect 106904 10854 106914 10906
rect 106914 10854 106960 10906
rect 106664 10852 106720 10854
rect 106744 10852 106800 10854
rect 106824 10852 106880 10854
rect 106904 10852 106960 10854
rect 105928 10362 105984 10364
rect 106008 10362 106064 10364
rect 106088 10362 106144 10364
rect 106168 10362 106224 10364
rect 105928 10310 105974 10362
rect 105974 10310 105984 10362
rect 106008 10310 106038 10362
rect 106038 10310 106050 10362
rect 106050 10310 106064 10362
rect 106088 10310 106102 10362
rect 106102 10310 106114 10362
rect 106114 10310 106144 10362
rect 106168 10310 106178 10362
rect 106178 10310 106224 10362
rect 105928 10308 105984 10310
rect 106008 10308 106064 10310
rect 106088 10308 106144 10310
rect 106168 10308 106224 10310
rect 106664 9818 106720 9820
rect 106744 9818 106800 9820
rect 106824 9818 106880 9820
rect 106904 9818 106960 9820
rect 106664 9766 106710 9818
rect 106710 9766 106720 9818
rect 106744 9766 106774 9818
rect 106774 9766 106786 9818
rect 106786 9766 106800 9818
rect 106824 9766 106838 9818
rect 106838 9766 106850 9818
rect 106850 9766 106880 9818
rect 106904 9766 106914 9818
rect 106914 9766 106960 9818
rect 106664 9764 106720 9766
rect 106744 9764 106800 9766
rect 106824 9764 106880 9766
rect 106904 9764 106960 9766
rect 105928 9274 105984 9276
rect 106008 9274 106064 9276
rect 106088 9274 106144 9276
rect 106168 9274 106224 9276
rect 105928 9222 105974 9274
rect 105974 9222 105984 9274
rect 106008 9222 106038 9274
rect 106038 9222 106050 9274
rect 106050 9222 106064 9274
rect 106088 9222 106102 9274
rect 106102 9222 106114 9274
rect 106114 9222 106144 9274
rect 106168 9222 106178 9274
rect 106178 9222 106224 9274
rect 105928 9220 105984 9222
rect 106008 9220 106064 9222
rect 106088 9220 106144 9222
rect 106168 9220 106224 9222
rect 106664 8730 106720 8732
rect 106744 8730 106800 8732
rect 106824 8730 106880 8732
rect 106904 8730 106960 8732
rect 106664 8678 106710 8730
rect 106710 8678 106720 8730
rect 106744 8678 106774 8730
rect 106774 8678 106786 8730
rect 106786 8678 106800 8730
rect 106824 8678 106838 8730
rect 106838 8678 106850 8730
rect 106850 8678 106880 8730
rect 106904 8678 106914 8730
rect 106914 8678 106960 8730
rect 106664 8676 106720 8678
rect 106744 8676 106800 8678
rect 106824 8676 106880 8678
rect 106904 8676 106960 8678
rect 105928 8186 105984 8188
rect 106008 8186 106064 8188
rect 106088 8186 106144 8188
rect 106168 8186 106224 8188
rect 105928 8134 105974 8186
rect 105974 8134 105984 8186
rect 106008 8134 106038 8186
rect 106038 8134 106050 8186
rect 106050 8134 106064 8186
rect 106088 8134 106102 8186
rect 106102 8134 106114 8186
rect 106114 8134 106144 8186
rect 106168 8134 106178 8186
rect 106178 8134 106224 8186
rect 105928 8132 105984 8134
rect 106008 8132 106064 8134
rect 106088 8132 106144 8134
rect 106168 8132 106224 8134
rect 97040 7642 97096 7644
rect 97120 7642 97176 7644
rect 97200 7642 97256 7644
rect 97280 7642 97336 7644
rect 97040 7590 97086 7642
rect 97086 7590 97096 7642
rect 97120 7590 97150 7642
rect 97150 7590 97162 7642
rect 97162 7590 97176 7642
rect 97200 7590 97214 7642
rect 97214 7590 97226 7642
rect 97226 7590 97256 7642
rect 97280 7590 97290 7642
rect 97290 7590 97336 7642
rect 97040 7588 97096 7590
rect 97120 7588 97176 7590
rect 97200 7588 97256 7590
rect 97280 7588 97336 7590
rect 106664 7642 106720 7644
rect 106744 7642 106800 7644
rect 106824 7642 106880 7644
rect 106904 7642 106960 7644
rect 106664 7590 106710 7642
rect 106710 7590 106720 7642
rect 106744 7590 106774 7642
rect 106774 7590 106786 7642
rect 106786 7590 106800 7642
rect 106824 7590 106838 7642
rect 106838 7590 106850 7642
rect 106850 7590 106880 7642
rect 106904 7590 106914 7642
rect 106914 7590 106960 7642
rect 106664 7588 106720 7590
rect 106744 7588 106800 7590
rect 106824 7588 106880 7590
rect 106904 7588 106960 7590
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 96380 7098 96436 7100
rect 96460 7098 96516 7100
rect 96540 7098 96596 7100
rect 96620 7098 96676 7100
rect 96380 7046 96426 7098
rect 96426 7046 96436 7098
rect 96460 7046 96490 7098
rect 96490 7046 96502 7098
rect 96502 7046 96516 7098
rect 96540 7046 96554 7098
rect 96554 7046 96566 7098
rect 96566 7046 96596 7098
rect 96620 7046 96630 7098
rect 96630 7046 96676 7098
rect 96380 7044 96436 7046
rect 96460 7044 96516 7046
rect 96540 7044 96596 7046
rect 96620 7044 96676 7046
rect 105928 7098 105984 7100
rect 106008 7098 106064 7100
rect 106088 7098 106144 7100
rect 106168 7098 106224 7100
rect 105928 7046 105974 7098
rect 105974 7046 105984 7098
rect 106008 7046 106038 7098
rect 106038 7046 106050 7098
rect 106050 7046 106064 7098
rect 106088 7046 106102 7098
rect 106102 7046 106114 7098
rect 106114 7046 106144 7098
rect 106168 7046 106178 7098
rect 106178 7046 106224 7098
rect 105928 7044 105984 7046
rect 106008 7044 106064 7046
rect 106088 7044 106144 7046
rect 106168 7044 106224 7046
rect 66320 6554 66376 6556
rect 66400 6554 66456 6556
rect 66480 6554 66536 6556
rect 66560 6554 66616 6556
rect 66320 6502 66366 6554
rect 66366 6502 66376 6554
rect 66400 6502 66430 6554
rect 66430 6502 66442 6554
rect 66442 6502 66456 6554
rect 66480 6502 66494 6554
rect 66494 6502 66506 6554
rect 66506 6502 66536 6554
rect 66560 6502 66570 6554
rect 66570 6502 66616 6554
rect 66320 6500 66376 6502
rect 66400 6500 66456 6502
rect 66480 6500 66536 6502
rect 66560 6500 66616 6502
rect 97040 6554 97096 6556
rect 97120 6554 97176 6556
rect 97200 6554 97256 6556
rect 97280 6554 97336 6556
rect 97040 6502 97086 6554
rect 97086 6502 97096 6554
rect 97120 6502 97150 6554
rect 97150 6502 97162 6554
rect 97162 6502 97176 6554
rect 97200 6502 97214 6554
rect 97214 6502 97226 6554
rect 97226 6502 97256 6554
rect 97280 6502 97290 6554
rect 97290 6502 97336 6554
rect 97040 6500 97096 6502
rect 97120 6500 97176 6502
rect 97200 6500 97256 6502
rect 97280 6500 97336 6502
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 96380 6010 96436 6012
rect 96460 6010 96516 6012
rect 96540 6010 96596 6012
rect 96620 6010 96676 6012
rect 96380 5958 96426 6010
rect 96426 5958 96436 6010
rect 96460 5958 96490 6010
rect 96490 5958 96502 6010
rect 96502 5958 96516 6010
rect 96540 5958 96554 6010
rect 96554 5958 96566 6010
rect 96566 5958 96596 6010
rect 96620 5958 96630 6010
rect 96630 5958 96676 6010
rect 96380 5956 96436 5958
rect 96460 5956 96516 5958
rect 96540 5956 96596 5958
rect 96620 5956 96676 5958
rect 66320 5466 66376 5468
rect 66400 5466 66456 5468
rect 66480 5466 66536 5468
rect 66560 5466 66616 5468
rect 66320 5414 66366 5466
rect 66366 5414 66376 5466
rect 66400 5414 66430 5466
rect 66430 5414 66442 5466
rect 66442 5414 66456 5466
rect 66480 5414 66494 5466
rect 66494 5414 66506 5466
rect 66506 5414 66536 5466
rect 66560 5414 66570 5466
rect 66570 5414 66616 5466
rect 66320 5412 66376 5414
rect 66400 5412 66456 5414
rect 66480 5412 66536 5414
rect 66560 5412 66616 5414
rect 97040 5466 97096 5468
rect 97120 5466 97176 5468
rect 97200 5466 97256 5468
rect 97280 5466 97336 5468
rect 97040 5414 97086 5466
rect 97086 5414 97096 5466
rect 97120 5414 97150 5466
rect 97150 5414 97162 5466
rect 97162 5414 97176 5466
rect 97200 5414 97214 5466
rect 97214 5414 97226 5466
rect 97226 5414 97256 5466
rect 97280 5414 97290 5466
rect 97290 5414 97336 5466
rect 97040 5412 97096 5414
rect 97120 5412 97176 5414
rect 97200 5412 97256 5414
rect 97280 5412 97336 5414
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 96380 4922 96436 4924
rect 96460 4922 96516 4924
rect 96540 4922 96596 4924
rect 96620 4922 96676 4924
rect 96380 4870 96426 4922
rect 96426 4870 96436 4922
rect 96460 4870 96490 4922
rect 96490 4870 96502 4922
rect 96502 4870 96516 4922
rect 96540 4870 96554 4922
rect 96554 4870 96566 4922
rect 96566 4870 96596 4922
rect 96620 4870 96630 4922
rect 96630 4870 96676 4922
rect 96380 4868 96436 4870
rect 96460 4868 96516 4870
rect 96540 4868 96596 4870
rect 96620 4868 96676 4870
rect 66320 4378 66376 4380
rect 66400 4378 66456 4380
rect 66480 4378 66536 4380
rect 66560 4378 66616 4380
rect 66320 4326 66366 4378
rect 66366 4326 66376 4378
rect 66400 4326 66430 4378
rect 66430 4326 66442 4378
rect 66442 4326 66456 4378
rect 66480 4326 66494 4378
rect 66494 4326 66506 4378
rect 66506 4326 66536 4378
rect 66560 4326 66570 4378
rect 66570 4326 66616 4378
rect 66320 4324 66376 4326
rect 66400 4324 66456 4326
rect 66480 4324 66536 4326
rect 66560 4324 66616 4326
rect 97040 4378 97096 4380
rect 97120 4378 97176 4380
rect 97200 4378 97256 4380
rect 97280 4378 97336 4380
rect 97040 4326 97086 4378
rect 97086 4326 97096 4378
rect 97120 4326 97150 4378
rect 97150 4326 97162 4378
rect 97162 4326 97176 4378
rect 97200 4326 97214 4378
rect 97214 4326 97226 4378
rect 97226 4326 97256 4378
rect 97280 4326 97290 4378
rect 97290 4326 97336 4378
rect 97040 4324 97096 4326
rect 97120 4324 97176 4326
rect 97200 4324 97256 4326
rect 97280 4324 97336 4326
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 96380 3834 96436 3836
rect 96460 3834 96516 3836
rect 96540 3834 96596 3836
rect 96620 3834 96676 3836
rect 96380 3782 96426 3834
rect 96426 3782 96436 3834
rect 96460 3782 96490 3834
rect 96490 3782 96502 3834
rect 96502 3782 96516 3834
rect 96540 3782 96554 3834
rect 96554 3782 96566 3834
rect 96566 3782 96596 3834
rect 96620 3782 96630 3834
rect 96630 3782 96676 3834
rect 96380 3780 96436 3782
rect 96460 3780 96516 3782
rect 96540 3780 96596 3782
rect 96620 3780 96676 3782
rect 66320 3290 66376 3292
rect 66400 3290 66456 3292
rect 66480 3290 66536 3292
rect 66560 3290 66616 3292
rect 66320 3238 66366 3290
rect 66366 3238 66376 3290
rect 66400 3238 66430 3290
rect 66430 3238 66442 3290
rect 66442 3238 66456 3290
rect 66480 3238 66494 3290
rect 66494 3238 66506 3290
rect 66506 3238 66536 3290
rect 66560 3238 66570 3290
rect 66570 3238 66616 3290
rect 66320 3236 66376 3238
rect 66400 3236 66456 3238
rect 66480 3236 66536 3238
rect 66560 3236 66616 3238
rect 97040 3290 97096 3292
rect 97120 3290 97176 3292
rect 97200 3290 97256 3292
rect 97280 3290 97336 3292
rect 97040 3238 97086 3290
rect 97086 3238 97096 3290
rect 97120 3238 97150 3290
rect 97150 3238 97162 3290
rect 97162 3238 97176 3290
rect 97200 3238 97214 3290
rect 97214 3238 97226 3290
rect 97226 3238 97256 3290
rect 97280 3238 97290 3290
rect 97290 3238 97336 3290
rect 97040 3236 97096 3238
rect 97120 3236 97176 3238
rect 97200 3236 97256 3238
rect 97280 3236 97336 3238
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 96380 2746 96436 2748
rect 96460 2746 96516 2748
rect 96540 2746 96596 2748
rect 96620 2746 96676 2748
rect 96380 2694 96426 2746
rect 96426 2694 96436 2746
rect 96460 2694 96490 2746
rect 96490 2694 96502 2746
rect 96502 2694 96516 2746
rect 96540 2694 96554 2746
rect 96554 2694 96566 2746
rect 96566 2694 96596 2746
rect 96620 2694 96630 2746
rect 96630 2694 96676 2746
rect 96380 2692 96436 2694
rect 96460 2692 96516 2694
rect 96540 2692 96596 2694
rect 96620 2692 96676 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 66320 2202 66376 2204
rect 66400 2202 66456 2204
rect 66480 2202 66536 2204
rect 66560 2202 66616 2204
rect 66320 2150 66366 2202
rect 66366 2150 66376 2202
rect 66400 2150 66430 2202
rect 66430 2150 66442 2202
rect 66442 2150 66456 2202
rect 66480 2150 66494 2202
rect 66494 2150 66506 2202
rect 66506 2150 66536 2202
rect 66560 2150 66570 2202
rect 66570 2150 66616 2202
rect 66320 2148 66376 2150
rect 66400 2148 66456 2150
rect 66480 2148 66536 2150
rect 66560 2148 66616 2150
rect 97040 2202 97096 2204
rect 97120 2202 97176 2204
rect 97200 2202 97256 2204
rect 97280 2202 97336 2204
rect 97040 2150 97086 2202
rect 97086 2150 97096 2202
rect 97120 2150 97150 2202
rect 97150 2150 97162 2202
rect 97162 2150 97176 2202
rect 97200 2150 97214 2202
rect 97214 2150 97226 2202
rect 97226 2150 97256 2202
rect 97280 2150 97290 2202
rect 97290 2150 97336 2202
rect 97040 2148 97096 2150
rect 97120 2148 97176 2150
rect 97200 2148 97256 2150
rect 97280 2148 97336 2150
<< metal3 >>
rect 4210 147456 4526 147457
rect 4210 147392 4216 147456
rect 4280 147392 4296 147456
rect 4360 147392 4376 147456
rect 4440 147392 4456 147456
rect 4520 147392 4526 147456
rect 4210 147391 4526 147392
rect 34930 147456 35246 147457
rect 34930 147392 34936 147456
rect 35000 147392 35016 147456
rect 35080 147392 35096 147456
rect 35160 147392 35176 147456
rect 35240 147392 35246 147456
rect 34930 147391 35246 147392
rect 65650 147456 65966 147457
rect 65650 147392 65656 147456
rect 65720 147392 65736 147456
rect 65800 147392 65816 147456
rect 65880 147392 65896 147456
rect 65960 147392 65966 147456
rect 65650 147391 65966 147392
rect 96370 147456 96686 147457
rect 96370 147392 96376 147456
rect 96440 147392 96456 147456
rect 96520 147392 96536 147456
rect 96600 147392 96616 147456
rect 96680 147392 96686 147456
rect 96370 147391 96686 147392
rect 4870 146912 5186 146913
rect 4870 146848 4876 146912
rect 4940 146848 4956 146912
rect 5020 146848 5036 146912
rect 5100 146848 5116 146912
rect 5180 146848 5186 146912
rect 4870 146847 5186 146848
rect 35590 146912 35906 146913
rect 35590 146848 35596 146912
rect 35660 146848 35676 146912
rect 35740 146848 35756 146912
rect 35820 146848 35836 146912
rect 35900 146848 35906 146912
rect 35590 146847 35906 146848
rect 66310 146912 66626 146913
rect 66310 146848 66316 146912
rect 66380 146848 66396 146912
rect 66460 146848 66476 146912
rect 66540 146848 66556 146912
rect 66620 146848 66626 146912
rect 66310 146847 66626 146848
rect 97030 146912 97346 146913
rect 97030 146848 97036 146912
rect 97100 146848 97116 146912
rect 97180 146848 97196 146912
rect 97260 146848 97276 146912
rect 97340 146848 97346 146912
rect 97030 146847 97346 146848
rect 4210 146368 4526 146369
rect 4210 146304 4216 146368
rect 4280 146304 4296 146368
rect 4360 146304 4376 146368
rect 4440 146304 4456 146368
rect 4520 146304 4526 146368
rect 4210 146303 4526 146304
rect 34930 146368 35246 146369
rect 34930 146304 34936 146368
rect 35000 146304 35016 146368
rect 35080 146304 35096 146368
rect 35160 146304 35176 146368
rect 35240 146304 35246 146368
rect 34930 146303 35246 146304
rect 65650 146368 65966 146369
rect 65650 146304 65656 146368
rect 65720 146304 65736 146368
rect 65800 146304 65816 146368
rect 65880 146304 65896 146368
rect 65960 146304 65966 146368
rect 65650 146303 65966 146304
rect 96370 146368 96686 146369
rect 96370 146304 96376 146368
rect 96440 146304 96456 146368
rect 96520 146304 96536 146368
rect 96600 146304 96616 146368
rect 96680 146304 96686 146368
rect 96370 146303 96686 146304
rect 4870 145824 5186 145825
rect 4870 145760 4876 145824
rect 4940 145760 4956 145824
rect 5020 145760 5036 145824
rect 5100 145760 5116 145824
rect 5180 145760 5186 145824
rect 4870 145759 5186 145760
rect 35590 145824 35906 145825
rect 35590 145760 35596 145824
rect 35660 145760 35676 145824
rect 35740 145760 35756 145824
rect 35820 145760 35836 145824
rect 35900 145760 35906 145824
rect 35590 145759 35906 145760
rect 66310 145824 66626 145825
rect 66310 145760 66316 145824
rect 66380 145760 66396 145824
rect 66460 145760 66476 145824
rect 66540 145760 66556 145824
rect 66620 145760 66626 145824
rect 66310 145759 66626 145760
rect 97030 145824 97346 145825
rect 97030 145760 97036 145824
rect 97100 145760 97116 145824
rect 97180 145760 97196 145824
rect 97260 145760 97276 145824
rect 97340 145760 97346 145824
rect 97030 145759 97346 145760
rect 4210 145280 4526 145281
rect 4210 145216 4216 145280
rect 4280 145216 4296 145280
rect 4360 145216 4376 145280
rect 4440 145216 4456 145280
rect 4520 145216 4526 145280
rect 4210 145215 4526 145216
rect 34930 145280 35246 145281
rect 34930 145216 34936 145280
rect 35000 145216 35016 145280
rect 35080 145216 35096 145280
rect 35160 145216 35176 145280
rect 35240 145216 35246 145280
rect 34930 145215 35246 145216
rect 65650 145280 65966 145281
rect 65650 145216 65656 145280
rect 65720 145216 65736 145280
rect 65800 145216 65816 145280
rect 65880 145216 65896 145280
rect 65960 145216 65966 145280
rect 65650 145215 65966 145216
rect 96370 145280 96686 145281
rect 96370 145216 96376 145280
rect 96440 145216 96456 145280
rect 96520 145216 96536 145280
rect 96600 145216 96616 145280
rect 96680 145216 96686 145280
rect 96370 145215 96686 145216
rect 4870 144736 5186 144737
rect 4870 144672 4876 144736
rect 4940 144672 4956 144736
rect 5020 144672 5036 144736
rect 5100 144672 5116 144736
rect 5180 144672 5186 144736
rect 4870 144671 5186 144672
rect 35590 144736 35906 144737
rect 35590 144672 35596 144736
rect 35660 144672 35676 144736
rect 35740 144672 35756 144736
rect 35820 144672 35836 144736
rect 35900 144672 35906 144736
rect 35590 144671 35906 144672
rect 66310 144736 66626 144737
rect 66310 144672 66316 144736
rect 66380 144672 66396 144736
rect 66460 144672 66476 144736
rect 66540 144672 66556 144736
rect 66620 144672 66626 144736
rect 66310 144671 66626 144672
rect 97030 144736 97346 144737
rect 97030 144672 97036 144736
rect 97100 144672 97116 144736
rect 97180 144672 97196 144736
rect 97260 144672 97276 144736
rect 97340 144672 97346 144736
rect 97030 144671 97346 144672
rect 4210 144192 4526 144193
rect 4210 144128 4216 144192
rect 4280 144128 4296 144192
rect 4360 144128 4376 144192
rect 4440 144128 4456 144192
rect 4520 144128 4526 144192
rect 4210 144127 4526 144128
rect 34930 144192 35246 144193
rect 34930 144128 34936 144192
rect 35000 144128 35016 144192
rect 35080 144128 35096 144192
rect 35160 144128 35176 144192
rect 35240 144128 35246 144192
rect 34930 144127 35246 144128
rect 65650 144192 65966 144193
rect 65650 144128 65656 144192
rect 65720 144128 65736 144192
rect 65800 144128 65816 144192
rect 65880 144128 65896 144192
rect 65960 144128 65966 144192
rect 65650 144127 65966 144128
rect 96370 144192 96686 144193
rect 96370 144128 96376 144192
rect 96440 144128 96456 144192
rect 96520 144128 96536 144192
rect 96600 144128 96616 144192
rect 96680 144128 96686 144192
rect 96370 144127 96686 144128
rect 4870 143648 5186 143649
rect 4870 143584 4876 143648
rect 4940 143584 4956 143648
rect 5020 143584 5036 143648
rect 5100 143584 5116 143648
rect 5180 143584 5186 143648
rect 4870 143583 5186 143584
rect 35590 143648 35906 143649
rect 35590 143584 35596 143648
rect 35660 143584 35676 143648
rect 35740 143584 35756 143648
rect 35820 143584 35836 143648
rect 35900 143584 35906 143648
rect 35590 143583 35906 143584
rect 66310 143648 66626 143649
rect 66310 143584 66316 143648
rect 66380 143584 66396 143648
rect 66460 143584 66476 143648
rect 66540 143584 66556 143648
rect 66620 143584 66626 143648
rect 66310 143583 66626 143584
rect 97030 143648 97346 143649
rect 97030 143584 97036 143648
rect 97100 143584 97116 143648
rect 97180 143584 97196 143648
rect 97260 143584 97276 143648
rect 97340 143584 97346 143648
rect 97030 143583 97346 143584
rect 4210 143104 4526 143105
rect 4210 143040 4216 143104
rect 4280 143040 4296 143104
rect 4360 143040 4376 143104
rect 4440 143040 4456 143104
rect 4520 143040 4526 143104
rect 4210 143039 4526 143040
rect 34930 143104 35246 143105
rect 34930 143040 34936 143104
rect 35000 143040 35016 143104
rect 35080 143040 35096 143104
rect 35160 143040 35176 143104
rect 35240 143040 35246 143104
rect 34930 143039 35246 143040
rect 65650 143104 65966 143105
rect 65650 143040 65656 143104
rect 65720 143040 65736 143104
rect 65800 143040 65816 143104
rect 65880 143040 65896 143104
rect 65960 143040 65966 143104
rect 65650 143039 65966 143040
rect 96370 143104 96686 143105
rect 96370 143040 96376 143104
rect 96440 143040 96456 143104
rect 96520 143040 96536 143104
rect 96600 143040 96616 143104
rect 96680 143040 96686 143104
rect 96370 143039 96686 143040
rect 4870 142560 5186 142561
rect 4870 142496 4876 142560
rect 4940 142496 4956 142560
rect 5020 142496 5036 142560
rect 5100 142496 5116 142560
rect 5180 142496 5186 142560
rect 4870 142495 5186 142496
rect 35590 142560 35906 142561
rect 35590 142496 35596 142560
rect 35660 142496 35676 142560
rect 35740 142496 35756 142560
rect 35820 142496 35836 142560
rect 35900 142496 35906 142560
rect 35590 142495 35906 142496
rect 66310 142560 66626 142561
rect 66310 142496 66316 142560
rect 66380 142496 66396 142560
rect 66460 142496 66476 142560
rect 66540 142496 66556 142560
rect 66620 142496 66626 142560
rect 66310 142495 66626 142496
rect 97030 142560 97346 142561
rect 97030 142496 97036 142560
rect 97100 142496 97116 142560
rect 97180 142496 97196 142560
rect 97260 142496 97276 142560
rect 97340 142496 97346 142560
rect 97030 142495 97346 142496
rect 4210 142016 4526 142017
rect 4210 141952 4216 142016
rect 4280 141952 4296 142016
rect 4360 141952 4376 142016
rect 4440 141952 4456 142016
rect 4520 141952 4526 142016
rect 4210 141951 4526 141952
rect 34930 142016 35246 142017
rect 34930 141952 34936 142016
rect 35000 141952 35016 142016
rect 35080 141952 35096 142016
rect 35160 141952 35176 142016
rect 35240 141952 35246 142016
rect 34930 141951 35246 141952
rect 65650 142016 65966 142017
rect 65650 141952 65656 142016
rect 65720 141952 65736 142016
rect 65800 141952 65816 142016
rect 65880 141952 65896 142016
rect 65960 141952 65966 142016
rect 65650 141951 65966 141952
rect 96370 142016 96686 142017
rect 96370 141952 96376 142016
rect 96440 141952 96456 142016
rect 96520 141952 96536 142016
rect 96600 141952 96616 142016
rect 96680 141952 96686 142016
rect 96370 141951 96686 141952
rect 4870 141472 5186 141473
rect 4870 141408 4876 141472
rect 4940 141408 4956 141472
rect 5020 141408 5036 141472
rect 5100 141408 5116 141472
rect 5180 141408 5186 141472
rect 4870 141407 5186 141408
rect 35590 141472 35906 141473
rect 35590 141408 35596 141472
rect 35660 141408 35676 141472
rect 35740 141408 35756 141472
rect 35820 141408 35836 141472
rect 35900 141408 35906 141472
rect 35590 141407 35906 141408
rect 66310 141472 66626 141473
rect 66310 141408 66316 141472
rect 66380 141408 66396 141472
rect 66460 141408 66476 141472
rect 66540 141408 66556 141472
rect 66620 141408 66626 141472
rect 66310 141407 66626 141408
rect 97030 141472 97346 141473
rect 97030 141408 97036 141472
rect 97100 141408 97116 141472
rect 97180 141408 97196 141472
rect 97260 141408 97276 141472
rect 97340 141408 97346 141472
rect 97030 141407 97346 141408
rect 4210 140928 4526 140929
rect 4210 140864 4216 140928
rect 4280 140864 4296 140928
rect 4360 140864 4376 140928
rect 4440 140864 4456 140928
rect 4520 140864 4526 140928
rect 4210 140863 4526 140864
rect 34930 140928 35246 140929
rect 34930 140864 34936 140928
rect 35000 140864 35016 140928
rect 35080 140864 35096 140928
rect 35160 140864 35176 140928
rect 35240 140864 35246 140928
rect 34930 140863 35246 140864
rect 65650 140928 65966 140929
rect 65650 140864 65656 140928
rect 65720 140864 65736 140928
rect 65800 140864 65816 140928
rect 65880 140864 65896 140928
rect 65960 140864 65966 140928
rect 65650 140863 65966 140864
rect 96370 140928 96686 140929
rect 96370 140864 96376 140928
rect 96440 140864 96456 140928
rect 96520 140864 96536 140928
rect 96600 140864 96616 140928
rect 96680 140864 96686 140928
rect 96370 140863 96686 140864
rect 4870 140384 5186 140385
rect 4870 140320 4876 140384
rect 4940 140320 4956 140384
rect 5020 140320 5036 140384
rect 5100 140320 5116 140384
rect 5180 140320 5186 140384
rect 4870 140319 5186 140320
rect 35590 140384 35906 140385
rect 35590 140320 35596 140384
rect 35660 140320 35676 140384
rect 35740 140320 35756 140384
rect 35820 140320 35836 140384
rect 35900 140320 35906 140384
rect 35590 140319 35906 140320
rect 66310 140384 66626 140385
rect 66310 140320 66316 140384
rect 66380 140320 66396 140384
rect 66460 140320 66476 140384
rect 66540 140320 66556 140384
rect 66620 140320 66626 140384
rect 66310 140319 66626 140320
rect 97030 140384 97346 140385
rect 97030 140320 97036 140384
rect 97100 140320 97116 140384
rect 97180 140320 97196 140384
rect 97260 140320 97276 140384
rect 97340 140320 97346 140384
rect 97030 140319 97346 140320
rect 4210 139840 4526 139841
rect 4210 139776 4216 139840
rect 4280 139776 4296 139840
rect 4360 139776 4376 139840
rect 4440 139776 4456 139840
rect 4520 139776 4526 139840
rect 4210 139775 4526 139776
rect 34930 139840 35246 139841
rect 34930 139776 34936 139840
rect 35000 139776 35016 139840
rect 35080 139776 35096 139840
rect 35160 139776 35176 139840
rect 35240 139776 35246 139840
rect 34930 139775 35246 139776
rect 65650 139840 65966 139841
rect 65650 139776 65656 139840
rect 65720 139776 65736 139840
rect 65800 139776 65816 139840
rect 65880 139776 65896 139840
rect 65960 139776 65966 139840
rect 65650 139775 65966 139776
rect 96370 139840 96686 139841
rect 96370 139776 96376 139840
rect 96440 139776 96456 139840
rect 96520 139776 96536 139840
rect 96600 139776 96616 139840
rect 96680 139776 96686 139840
rect 96370 139775 96686 139776
rect 4870 139296 5186 139297
rect 4870 139232 4876 139296
rect 4940 139232 4956 139296
rect 5020 139232 5036 139296
rect 5100 139232 5116 139296
rect 5180 139232 5186 139296
rect 4870 139231 5186 139232
rect 35590 139296 35906 139297
rect 35590 139232 35596 139296
rect 35660 139232 35676 139296
rect 35740 139232 35756 139296
rect 35820 139232 35836 139296
rect 35900 139232 35906 139296
rect 35590 139231 35906 139232
rect 66310 139296 66626 139297
rect 66310 139232 66316 139296
rect 66380 139232 66396 139296
rect 66460 139232 66476 139296
rect 66540 139232 66556 139296
rect 66620 139232 66626 139296
rect 66310 139231 66626 139232
rect 97030 139296 97346 139297
rect 97030 139232 97036 139296
rect 97100 139232 97116 139296
rect 97180 139232 97196 139296
rect 97260 139232 97276 139296
rect 97340 139232 97346 139296
rect 97030 139231 97346 139232
rect 4210 138752 4526 138753
rect 4210 138688 4216 138752
rect 4280 138688 4296 138752
rect 4360 138688 4376 138752
rect 4440 138688 4456 138752
rect 4520 138688 4526 138752
rect 4210 138687 4526 138688
rect 34930 138752 35246 138753
rect 34930 138688 34936 138752
rect 35000 138688 35016 138752
rect 35080 138688 35096 138752
rect 35160 138688 35176 138752
rect 35240 138688 35246 138752
rect 34930 138687 35246 138688
rect 65650 138752 65966 138753
rect 65650 138688 65656 138752
rect 65720 138688 65736 138752
rect 65800 138688 65816 138752
rect 65880 138688 65896 138752
rect 65960 138688 65966 138752
rect 65650 138687 65966 138688
rect 96370 138752 96686 138753
rect 96370 138688 96376 138752
rect 96440 138688 96456 138752
rect 96520 138688 96536 138752
rect 96600 138688 96616 138752
rect 96680 138688 96686 138752
rect 96370 138687 96686 138688
rect 4870 138208 5186 138209
rect 4870 138144 4876 138208
rect 4940 138144 4956 138208
rect 5020 138144 5036 138208
rect 5100 138144 5116 138208
rect 5180 138144 5186 138208
rect 4870 138143 5186 138144
rect 35590 138208 35906 138209
rect 35590 138144 35596 138208
rect 35660 138144 35676 138208
rect 35740 138144 35756 138208
rect 35820 138144 35836 138208
rect 35900 138144 35906 138208
rect 35590 138143 35906 138144
rect 66310 138208 66626 138209
rect 66310 138144 66316 138208
rect 66380 138144 66396 138208
rect 66460 138144 66476 138208
rect 66540 138144 66556 138208
rect 66620 138144 66626 138208
rect 66310 138143 66626 138144
rect 97030 138208 97346 138209
rect 97030 138144 97036 138208
rect 97100 138144 97116 138208
rect 97180 138144 97196 138208
rect 97260 138144 97276 138208
rect 97340 138144 97346 138208
rect 97030 138143 97346 138144
rect 4210 137664 4526 137665
rect 4210 137600 4216 137664
rect 4280 137600 4296 137664
rect 4360 137600 4376 137664
rect 4440 137600 4456 137664
rect 4520 137600 4526 137664
rect 4210 137599 4526 137600
rect 34930 137664 35246 137665
rect 34930 137600 34936 137664
rect 35000 137600 35016 137664
rect 35080 137600 35096 137664
rect 35160 137600 35176 137664
rect 35240 137600 35246 137664
rect 34930 137599 35246 137600
rect 65650 137664 65966 137665
rect 65650 137600 65656 137664
rect 65720 137600 65736 137664
rect 65800 137600 65816 137664
rect 65880 137600 65896 137664
rect 65960 137600 65966 137664
rect 65650 137599 65966 137600
rect 96370 137664 96686 137665
rect 96370 137600 96376 137664
rect 96440 137600 96456 137664
rect 96520 137600 96536 137664
rect 96600 137600 96616 137664
rect 96680 137600 96686 137664
rect 96370 137599 96686 137600
rect 4870 137120 5186 137121
rect 4870 137056 4876 137120
rect 4940 137056 4956 137120
rect 5020 137056 5036 137120
rect 5100 137056 5116 137120
rect 5180 137056 5186 137120
rect 4870 137055 5186 137056
rect 35590 137120 35906 137121
rect 35590 137056 35596 137120
rect 35660 137056 35676 137120
rect 35740 137056 35756 137120
rect 35820 137056 35836 137120
rect 35900 137056 35906 137120
rect 35590 137055 35906 137056
rect 66310 137120 66626 137121
rect 66310 137056 66316 137120
rect 66380 137056 66396 137120
rect 66460 137056 66476 137120
rect 66540 137056 66556 137120
rect 66620 137056 66626 137120
rect 66310 137055 66626 137056
rect 97030 137120 97346 137121
rect 97030 137056 97036 137120
rect 97100 137056 97116 137120
rect 97180 137056 97196 137120
rect 97260 137056 97276 137120
rect 97340 137056 97346 137120
rect 97030 137055 97346 137056
rect 4210 136576 4526 136577
rect 4210 136512 4216 136576
rect 4280 136512 4296 136576
rect 4360 136512 4376 136576
rect 4440 136512 4456 136576
rect 4520 136512 4526 136576
rect 4210 136511 4526 136512
rect 34930 136576 35246 136577
rect 34930 136512 34936 136576
rect 35000 136512 35016 136576
rect 35080 136512 35096 136576
rect 35160 136512 35176 136576
rect 35240 136512 35246 136576
rect 34930 136511 35246 136512
rect 65650 136576 65966 136577
rect 65650 136512 65656 136576
rect 65720 136512 65736 136576
rect 65800 136512 65816 136576
rect 65880 136512 65896 136576
rect 65960 136512 65966 136576
rect 65650 136511 65966 136512
rect 96370 136576 96686 136577
rect 96370 136512 96376 136576
rect 96440 136512 96456 136576
rect 96520 136512 96536 136576
rect 96600 136512 96616 136576
rect 96680 136512 96686 136576
rect 96370 136511 96686 136512
rect 105918 136576 106234 136577
rect 105918 136512 105924 136576
rect 105988 136512 106004 136576
rect 106068 136512 106084 136576
rect 106148 136512 106164 136576
rect 106228 136512 106234 136576
rect 105918 136511 106234 136512
rect 4870 136032 5186 136033
rect 4870 135968 4876 136032
rect 4940 135968 4956 136032
rect 5020 135968 5036 136032
rect 5100 135968 5116 136032
rect 5180 135968 5186 136032
rect 4870 135967 5186 135968
rect 35590 136032 35906 136033
rect 35590 135968 35596 136032
rect 35660 135968 35676 136032
rect 35740 135968 35756 136032
rect 35820 135968 35836 136032
rect 35900 135968 35906 136032
rect 35590 135967 35906 135968
rect 66310 136032 66626 136033
rect 66310 135968 66316 136032
rect 66380 135968 66396 136032
rect 66460 135968 66476 136032
rect 66540 135968 66556 136032
rect 66620 135968 66626 136032
rect 66310 135967 66626 135968
rect 97030 136032 97346 136033
rect 97030 135968 97036 136032
rect 97100 135968 97116 136032
rect 97180 135968 97196 136032
rect 97260 135968 97276 136032
rect 97340 135968 97346 136032
rect 97030 135967 97346 135968
rect 106654 136032 106970 136033
rect 106654 135968 106660 136032
rect 106724 135968 106740 136032
rect 106804 135968 106820 136032
rect 106884 135968 106900 136032
rect 106964 135968 106970 136032
rect 106654 135967 106970 135968
rect 4210 135488 4526 135489
rect 4210 135424 4216 135488
rect 4280 135424 4296 135488
rect 4360 135424 4376 135488
rect 4440 135424 4456 135488
rect 4520 135424 4526 135488
rect 4210 135423 4526 135424
rect 105918 135488 106234 135489
rect 105918 135424 105924 135488
rect 105988 135424 106004 135488
rect 106068 135424 106084 135488
rect 106148 135424 106164 135488
rect 106228 135424 106234 135488
rect 105918 135423 106234 135424
rect 58566 135220 58572 135284
rect 58636 135282 58642 135284
rect 60641 135282 60707 135285
rect 58636 135280 60707 135282
rect 58636 135224 60646 135280
rect 60702 135224 60707 135280
rect 58636 135222 60707 135224
rect 58636 135220 58642 135222
rect 60641 135219 60707 135222
rect 61142 135220 61148 135284
rect 61212 135282 61218 135284
rect 63125 135282 63191 135285
rect 61212 135280 63191 135282
rect 61212 135224 63130 135280
rect 63186 135224 63191 135280
rect 61212 135222 63191 135224
rect 61212 135220 61218 135222
rect 63125 135219 63191 135222
rect 66110 135220 66116 135284
rect 66180 135282 66186 135284
rect 67541 135282 67607 135285
rect 66180 135280 67607 135282
rect 66180 135224 67546 135280
rect 67602 135224 67607 135280
rect 66180 135222 67607 135224
rect 66180 135220 66186 135222
rect 67541 135219 67607 135222
rect 68502 135220 68508 135284
rect 68572 135282 68578 135284
rect 69749 135282 69815 135285
rect 68572 135280 69815 135282
rect 68572 135224 69754 135280
rect 69810 135224 69815 135280
rect 68572 135222 69815 135224
rect 68572 135220 68578 135222
rect 69749 135219 69815 135222
rect 71078 135220 71084 135284
rect 71148 135282 71154 135284
rect 72141 135282 72207 135285
rect 71148 135280 72207 135282
rect 71148 135224 72146 135280
rect 72202 135224 72207 135280
rect 71148 135222 72207 135224
rect 71148 135220 71154 135222
rect 72141 135219 72207 135222
rect 63534 135084 63540 135148
rect 63604 135146 63610 135148
rect 64413 135146 64479 135149
rect 63604 135144 64479 135146
rect 63604 135088 64418 135144
rect 64474 135088 64479 135144
rect 63604 135086 64479 135088
rect 63604 135084 63610 135086
rect 64413 135083 64479 135086
rect 4870 134944 5186 134945
rect 4870 134880 4876 134944
rect 4940 134880 4956 134944
rect 5020 134880 5036 134944
rect 5100 134880 5116 134944
rect 5180 134880 5186 134944
rect 4870 134879 5186 134880
rect 106654 134944 106970 134945
rect 106654 134880 106660 134944
rect 106724 134880 106740 134944
rect 106804 134880 106820 134944
rect 106884 134880 106900 134944
rect 106964 134880 106970 134944
rect 106654 134879 106970 134880
rect 95969 134468 96035 134469
rect 95918 134466 95924 134468
rect 95878 134406 95924 134466
rect 95988 134464 96035 134468
rect 96030 134408 96035 134464
rect 95918 134404 95924 134406
rect 95988 134404 96035 134408
rect 95969 134403 96035 134404
rect 4210 134400 4526 134401
rect 4210 134336 4216 134400
rect 4280 134336 4296 134400
rect 4360 134336 4376 134400
rect 4440 134336 4456 134400
rect 4520 134336 4526 134400
rect 4210 134335 4526 134336
rect 105918 134400 106234 134401
rect 105918 134336 105924 134400
rect 105988 134336 106004 134400
rect 106068 134336 106084 134400
rect 106148 134336 106164 134400
rect 106228 134336 106234 134400
rect 105918 134335 106234 134336
rect 38193 134194 38259 134197
rect 38565 134194 38571 134196
rect 38193 134192 38571 134194
rect 38193 134136 38198 134192
rect 38254 134136 38571 134192
rect 38193 134134 38571 134136
rect 38193 134131 38259 134134
rect 38565 134132 38571 134134
rect 38635 134132 38641 134196
rect 40677 134194 40743 134197
rect 41061 134194 41067 134196
rect 40677 134192 41067 134194
rect 40677 134136 40682 134192
rect 40738 134136 41067 134192
rect 40677 134134 41067 134136
rect 40677 134131 40743 134134
rect 41061 134132 41067 134134
rect 41131 134132 41137 134196
rect 51045 134132 51051 134196
rect 51115 134194 51121 134196
rect 52361 134194 52427 134197
rect 51115 134192 52427 134194
rect 51115 134136 52366 134192
rect 52422 134136 52427 134192
rect 51115 134134 52427 134136
rect 51115 134132 51121 134134
rect 52361 134131 52427 134134
rect 56037 134132 56043 134196
rect 56107 134194 56113 134196
rect 58157 134194 58223 134197
rect 56107 134192 58223 134194
rect 56107 134136 58162 134192
rect 58218 134136 58223 134192
rect 56107 134134 58223 134136
rect 56107 134132 56113 134134
rect 58157 134131 58223 134134
rect 73509 134132 73515 134196
rect 73579 134194 73585 134196
rect 74165 134194 74231 134197
rect 73579 134192 74231 134194
rect 73579 134136 74170 134192
rect 74226 134136 74231 134192
rect 73579 134134 74231 134136
rect 73579 134132 73585 134134
rect 74165 134131 74231 134134
rect 53541 133996 53547 134060
rect 53611 134058 53617 134060
rect 55765 134058 55831 134061
rect 53611 134056 55831 134058
rect 53611 134000 55770 134056
rect 55826 134000 55831 134056
rect 53611 133998 55831 134000
rect 53611 133996 53617 133998
rect 55765 133995 55831 133998
rect 36077 133924 36143 133925
rect 36069 133922 36075 133924
rect 35986 133862 36075 133922
rect 36069 133860 36075 133862
rect 36139 133860 36145 133924
rect 42977 133922 43043 133925
rect 46013 133924 46079 133925
rect 48497 133924 48563 133925
rect 86125 133924 86191 133925
rect 87321 133924 87387 133925
rect 43557 133922 43563 133924
rect 42977 133920 43563 133922
rect 42977 133864 42982 133920
rect 43038 133864 43563 133920
rect 42977 133862 43563 133864
rect 36077 133859 36143 133860
rect 42977 133859 43043 133862
rect 43557 133860 43563 133862
rect 43627 133860 43633 133924
rect 46013 133920 46059 133924
rect 46123 133922 46129 133924
rect 46013 133864 46018 133920
rect 46013 133860 46059 133864
rect 46123 133862 46170 133922
rect 48497 133920 48544 133924
rect 48608 133922 48614 133924
rect 48497 133864 48502 133920
rect 46123 133860 46129 133862
rect 48497 133860 48544 133864
rect 48608 133862 48654 133922
rect 86125 133920 86142 133924
rect 86206 133922 86212 133924
rect 87304 133922 87310 133924
rect 86125 133864 86130 133920
rect 48608 133860 48614 133862
rect 86125 133860 86142 133864
rect 86206 133862 86282 133922
rect 87230 133862 87310 133922
rect 87374 133920 87387 133924
rect 87382 133864 87387 133920
rect 86206 133860 86212 133862
rect 87304 133860 87310 133862
rect 87374 133860 87387 133864
rect 46013 133859 46079 133860
rect 48497 133859 48563 133860
rect 86125 133859 86191 133860
rect 87321 133859 87387 133860
rect 4870 133856 5186 133857
rect 4870 133792 4876 133856
rect 4940 133792 4956 133856
rect 5020 133792 5036 133856
rect 5100 133792 5116 133856
rect 5180 133792 5186 133856
rect 4870 133791 5186 133792
rect 106654 133856 106970 133857
rect 106654 133792 106660 133856
rect 106724 133792 106740 133856
rect 106804 133792 106820 133856
rect 106884 133792 106900 133856
rect 106964 133792 106970 133856
rect 106654 133791 106970 133792
rect 4210 133312 4526 133313
rect 4210 133248 4216 133312
rect 4280 133248 4296 133312
rect 4360 133248 4376 133312
rect 4440 133248 4456 133312
rect 4520 133248 4526 133312
rect 4210 133247 4526 133248
rect 105918 133312 106234 133313
rect 105918 133248 105924 133312
rect 105988 133248 106004 133312
rect 106068 133248 106084 133312
rect 106148 133248 106164 133312
rect 106228 133248 106234 133312
rect 105918 133247 106234 133248
rect 4870 132768 5186 132769
rect 4870 132704 4876 132768
rect 4940 132704 4956 132768
rect 5020 132704 5036 132768
rect 5100 132704 5116 132768
rect 5180 132704 5186 132768
rect 4870 132703 5186 132704
rect 106654 132768 106970 132769
rect 106654 132704 106660 132768
rect 106724 132704 106740 132768
rect 106804 132704 106820 132768
rect 106884 132704 106900 132768
rect 106964 132704 106970 132768
rect 106654 132703 106970 132704
rect 4210 132224 4526 132225
rect 4210 132160 4216 132224
rect 4280 132160 4296 132224
rect 4360 132160 4376 132224
rect 4440 132160 4456 132224
rect 4520 132160 4526 132224
rect 4210 132159 4526 132160
rect 105918 132224 106234 132225
rect 105918 132160 105924 132224
rect 105988 132160 106004 132224
rect 106068 132160 106084 132224
rect 106148 132160 106164 132224
rect 106228 132160 106234 132224
rect 105918 132159 106234 132160
rect 4870 131680 5186 131681
rect 4870 131616 4876 131680
rect 4940 131616 4956 131680
rect 5020 131616 5036 131680
rect 5100 131616 5116 131680
rect 5180 131616 5186 131680
rect 4870 131615 5186 131616
rect 106654 131680 106970 131681
rect 106654 131616 106660 131680
rect 106724 131616 106740 131680
rect 106804 131616 106820 131680
rect 106884 131616 106900 131680
rect 106964 131616 106970 131680
rect 106654 131615 106970 131616
rect 4210 131136 4526 131137
rect 4210 131072 4216 131136
rect 4280 131072 4296 131136
rect 4360 131072 4376 131136
rect 4440 131072 4456 131136
rect 4520 131072 4526 131136
rect 4210 131071 4526 131072
rect 105918 131136 106234 131137
rect 105918 131072 105924 131136
rect 105988 131072 106004 131136
rect 106068 131072 106084 131136
rect 106148 131072 106164 131136
rect 106228 131072 106234 131136
rect 105918 131071 106234 131072
rect 4870 130592 5186 130593
rect 4870 130528 4876 130592
rect 4940 130528 4956 130592
rect 5020 130528 5036 130592
rect 5100 130528 5116 130592
rect 5180 130528 5186 130592
rect 4870 130527 5186 130528
rect 106654 130592 106970 130593
rect 106654 130528 106660 130592
rect 106724 130528 106740 130592
rect 106804 130528 106820 130592
rect 106884 130528 106900 130592
rect 106964 130528 106970 130592
rect 106654 130527 106970 130528
rect 4210 130048 4526 130049
rect 4210 129984 4216 130048
rect 4280 129984 4296 130048
rect 4360 129984 4376 130048
rect 4440 129984 4456 130048
rect 4520 129984 4526 130048
rect 4210 129983 4526 129984
rect 105918 130048 106234 130049
rect 105918 129984 105924 130048
rect 105988 129984 106004 130048
rect 106068 129984 106084 130048
rect 106148 129984 106164 130048
rect 106228 129984 106234 130048
rect 105918 129983 106234 129984
rect 104341 129842 104407 129845
rect 102550 129840 104407 129842
rect 102550 129784 104346 129840
rect 104402 129784 104407 129840
rect 102550 129782 104407 129784
rect 102550 129768 102610 129782
rect 104341 129779 104407 129782
rect 101948 129708 102610 129768
rect 4870 129504 5186 129505
rect 4870 129440 4876 129504
rect 4940 129440 4956 129504
rect 5020 129440 5036 129504
rect 5100 129440 5116 129504
rect 5180 129440 5186 129504
rect 4870 129439 5186 129440
rect 106654 129504 106970 129505
rect 106654 129440 106660 129504
rect 106724 129440 106740 129504
rect 106804 129440 106820 129504
rect 106884 129440 106900 129504
rect 106964 129440 106970 129504
rect 106654 129439 106970 129440
rect 4210 128960 4526 128961
rect 4210 128896 4216 128960
rect 4280 128896 4296 128960
rect 4360 128896 4376 128960
rect 4440 128896 4456 128960
rect 4520 128896 4526 128960
rect 4210 128895 4526 128896
rect 105918 128960 106234 128961
rect 105918 128896 105924 128960
rect 105988 128896 106004 128960
rect 106068 128896 106084 128960
rect 106148 128896 106164 128960
rect 106228 128896 106234 128960
rect 105918 128895 106234 128896
rect 4870 128416 5186 128417
rect 4870 128352 4876 128416
rect 4940 128352 4956 128416
rect 5020 128352 5036 128416
rect 5100 128352 5116 128416
rect 5180 128352 5186 128416
rect 4870 128351 5186 128352
rect 106654 128416 106970 128417
rect 106654 128352 106660 128416
rect 106724 128352 106740 128416
rect 106804 128352 106820 128416
rect 106884 128352 106900 128416
rect 106964 128352 106970 128416
rect 106654 128351 106970 128352
rect 4210 127872 4526 127873
rect 4210 127808 4216 127872
rect 4280 127808 4296 127872
rect 4360 127808 4376 127872
rect 4440 127808 4456 127872
rect 4520 127808 4526 127872
rect 4210 127807 4526 127808
rect 105918 127872 106234 127873
rect 105918 127808 105924 127872
rect 105988 127808 106004 127872
rect 106068 127808 106084 127872
rect 106148 127808 106164 127872
rect 106228 127808 106234 127872
rect 105918 127807 106234 127808
rect 4870 127328 5186 127329
rect 4870 127264 4876 127328
rect 4940 127264 4956 127328
rect 5020 127264 5036 127328
rect 5100 127264 5116 127328
rect 5180 127264 5186 127328
rect 4870 127263 5186 127264
rect 106654 127328 106970 127329
rect 106654 127264 106660 127328
rect 106724 127264 106740 127328
rect 106804 127264 106820 127328
rect 106884 127264 106900 127328
rect 106964 127264 106970 127328
rect 106654 127263 106970 127264
rect 4210 126784 4526 126785
rect 4210 126720 4216 126784
rect 4280 126720 4296 126784
rect 4360 126720 4376 126784
rect 4440 126720 4456 126784
rect 4520 126720 4526 126784
rect 4210 126719 4526 126720
rect 105918 126784 106234 126785
rect 105918 126720 105924 126784
rect 105988 126720 106004 126784
rect 106068 126720 106084 126784
rect 106148 126720 106164 126784
rect 106228 126720 106234 126784
rect 105918 126719 106234 126720
rect 4870 126240 5186 126241
rect 4870 126176 4876 126240
rect 4940 126176 4956 126240
rect 5020 126176 5036 126240
rect 5100 126176 5116 126240
rect 5180 126176 5186 126240
rect 4870 126175 5186 126176
rect 106654 126240 106970 126241
rect 106654 126176 106660 126240
rect 106724 126176 106740 126240
rect 106804 126176 106820 126240
rect 106884 126176 106900 126240
rect 106964 126176 106970 126240
rect 106654 126175 106970 126176
rect 4210 125696 4526 125697
rect 4210 125632 4216 125696
rect 4280 125632 4296 125696
rect 4360 125632 4376 125696
rect 4440 125632 4456 125696
rect 4520 125632 4526 125696
rect 4210 125631 4526 125632
rect 105918 125696 106234 125697
rect 105918 125632 105924 125696
rect 105988 125632 106004 125696
rect 106068 125632 106084 125696
rect 106148 125632 106164 125696
rect 106228 125632 106234 125696
rect 105918 125631 106234 125632
rect 4870 125152 5186 125153
rect 4870 125088 4876 125152
rect 4940 125088 4956 125152
rect 5020 125088 5036 125152
rect 5100 125088 5116 125152
rect 5180 125088 5186 125152
rect 4870 125087 5186 125088
rect 106654 125152 106970 125153
rect 106654 125088 106660 125152
rect 106724 125088 106740 125152
rect 106804 125088 106820 125152
rect 106884 125088 106900 125152
rect 106964 125088 106970 125152
rect 106654 125087 106970 125088
rect 4210 124608 4526 124609
rect 4210 124544 4216 124608
rect 4280 124544 4296 124608
rect 4360 124544 4376 124608
rect 4440 124544 4456 124608
rect 4520 124544 4526 124608
rect 4210 124543 4526 124544
rect 105918 124608 106234 124609
rect 105918 124544 105924 124608
rect 105988 124544 106004 124608
rect 106068 124544 106084 124608
rect 106148 124544 106164 124608
rect 106228 124544 106234 124608
rect 105918 124543 106234 124544
rect 4870 124064 5186 124065
rect 4870 124000 4876 124064
rect 4940 124000 4956 124064
rect 5020 124000 5036 124064
rect 5100 124000 5116 124064
rect 5180 124000 5186 124064
rect 4870 123999 5186 124000
rect 106654 124064 106970 124065
rect 106654 124000 106660 124064
rect 106724 124000 106740 124064
rect 106804 124000 106820 124064
rect 106884 124000 106900 124064
rect 106964 124000 106970 124064
rect 106654 123999 106970 124000
rect 4210 123520 4526 123521
rect 4210 123456 4216 123520
rect 4280 123456 4296 123520
rect 4360 123456 4376 123520
rect 4440 123456 4456 123520
rect 4520 123456 4526 123520
rect 4210 123455 4526 123456
rect 105918 123520 106234 123521
rect 105918 123456 105924 123520
rect 105988 123456 106004 123520
rect 106068 123456 106084 123520
rect 106148 123456 106164 123520
rect 106228 123456 106234 123520
rect 105918 123455 106234 123456
rect 4870 122976 5186 122977
rect 4870 122912 4876 122976
rect 4940 122912 4956 122976
rect 5020 122912 5036 122976
rect 5100 122912 5116 122976
rect 5180 122912 5186 122976
rect 4870 122911 5186 122912
rect 106654 122976 106970 122977
rect 106654 122912 106660 122976
rect 106724 122912 106740 122976
rect 106804 122912 106820 122976
rect 106884 122912 106900 122976
rect 106964 122912 106970 122976
rect 106654 122911 106970 122912
rect 4210 122432 4526 122433
rect 4210 122368 4216 122432
rect 4280 122368 4296 122432
rect 4360 122368 4376 122432
rect 4440 122368 4456 122432
rect 4520 122368 4526 122432
rect 4210 122367 4526 122368
rect 105918 122432 106234 122433
rect 105918 122368 105924 122432
rect 105988 122368 106004 122432
rect 106068 122368 106084 122432
rect 106148 122368 106164 122432
rect 106228 122368 106234 122432
rect 105918 122367 106234 122368
rect 4870 121888 5186 121889
rect 4870 121824 4876 121888
rect 4940 121824 4956 121888
rect 5020 121824 5036 121888
rect 5100 121824 5116 121888
rect 5180 121824 5186 121888
rect 4870 121823 5186 121824
rect 106654 121888 106970 121889
rect 106654 121824 106660 121888
rect 106724 121824 106740 121888
rect 106804 121824 106820 121888
rect 106884 121824 106900 121888
rect 106964 121824 106970 121888
rect 106654 121823 106970 121824
rect 4210 121344 4526 121345
rect 4210 121280 4216 121344
rect 4280 121280 4296 121344
rect 4360 121280 4376 121344
rect 4440 121280 4456 121344
rect 4520 121280 4526 121344
rect 4210 121279 4526 121280
rect 105918 121344 106234 121345
rect 105918 121280 105924 121344
rect 105988 121280 106004 121344
rect 106068 121280 106084 121344
rect 106148 121280 106164 121344
rect 106228 121280 106234 121344
rect 105918 121279 106234 121280
rect 4870 120800 5186 120801
rect 4870 120736 4876 120800
rect 4940 120736 4956 120800
rect 5020 120736 5036 120800
rect 5100 120736 5116 120800
rect 5180 120736 5186 120800
rect 4870 120735 5186 120736
rect 106654 120800 106970 120801
rect 106654 120736 106660 120800
rect 106724 120736 106740 120800
rect 106804 120736 106820 120800
rect 106884 120736 106900 120800
rect 106964 120736 106970 120800
rect 106654 120735 106970 120736
rect 4210 120256 4526 120257
rect 4210 120192 4216 120256
rect 4280 120192 4296 120256
rect 4360 120192 4376 120256
rect 4440 120192 4456 120256
rect 4520 120192 4526 120256
rect 4210 120191 4526 120192
rect 105918 120256 106234 120257
rect 105918 120192 105924 120256
rect 105988 120192 106004 120256
rect 106068 120192 106084 120256
rect 106148 120192 106164 120256
rect 106228 120192 106234 120256
rect 105918 120191 106234 120192
rect 4870 119712 5186 119713
rect 4870 119648 4876 119712
rect 4940 119648 4956 119712
rect 5020 119648 5036 119712
rect 5100 119648 5116 119712
rect 5180 119648 5186 119712
rect 4870 119647 5186 119648
rect 106654 119712 106970 119713
rect 106654 119648 106660 119712
rect 106724 119648 106740 119712
rect 106804 119648 106820 119712
rect 106884 119648 106900 119712
rect 106964 119648 106970 119712
rect 106654 119647 106970 119648
rect 4210 119168 4526 119169
rect 4210 119104 4216 119168
rect 4280 119104 4296 119168
rect 4360 119104 4376 119168
rect 4440 119104 4456 119168
rect 4520 119104 4526 119168
rect 4210 119103 4526 119104
rect 105918 119168 106234 119169
rect 105918 119104 105924 119168
rect 105988 119104 106004 119168
rect 106068 119104 106084 119168
rect 106148 119104 106164 119168
rect 106228 119104 106234 119168
rect 105918 119103 106234 119104
rect 4870 118624 5186 118625
rect 4870 118560 4876 118624
rect 4940 118560 4956 118624
rect 5020 118560 5036 118624
rect 5100 118560 5116 118624
rect 5180 118560 5186 118624
rect 4870 118559 5186 118560
rect 106654 118624 106970 118625
rect 106654 118560 106660 118624
rect 106724 118560 106740 118624
rect 106804 118560 106820 118624
rect 106884 118560 106900 118624
rect 106964 118560 106970 118624
rect 106654 118559 106970 118560
rect 4210 118080 4526 118081
rect 4210 118016 4216 118080
rect 4280 118016 4296 118080
rect 4360 118016 4376 118080
rect 4440 118016 4456 118080
rect 4520 118016 4526 118080
rect 4210 118015 4526 118016
rect 105918 118080 106234 118081
rect 105918 118016 105924 118080
rect 105988 118016 106004 118080
rect 106068 118016 106084 118080
rect 106148 118016 106164 118080
rect 106228 118016 106234 118080
rect 105918 118015 106234 118016
rect 4870 117536 5186 117537
rect 4870 117472 4876 117536
rect 4940 117472 4956 117536
rect 5020 117472 5036 117536
rect 5100 117472 5116 117536
rect 5180 117472 5186 117536
rect 4870 117471 5186 117472
rect 106654 117536 106970 117537
rect 106654 117472 106660 117536
rect 106724 117472 106740 117536
rect 106804 117472 106820 117536
rect 106884 117472 106900 117536
rect 106964 117472 106970 117536
rect 106654 117471 106970 117472
rect 4210 116992 4526 116993
rect 4210 116928 4216 116992
rect 4280 116928 4296 116992
rect 4360 116928 4376 116992
rect 4440 116928 4456 116992
rect 4520 116928 4526 116992
rect 4210 116927 4526 116928
rect 105918 116992 106234 116993
rect 105918 116928 105924 116992
rect 105988 116928 106004 116992
rect 106068 116928 106084 116992
rect 106148 116928 106164 116992
rect 106228 116928 106234 116992
rect 105918 116927 106234 116928
rect 4870 116448 5186 116449
rect 4870 116384 4876 116448
rect 4940 116384 4956 116448
rect 5020 116384 5036 116448
rect 5100 116384 5116 116448
rect 5180 116384 5186 116448
rect 4870 116383 5186 116384
rect 106654 116448 106970 116449
rect 106654 116384 106660 116448
rect 106724 116384 106740 116448
rect 106804 116384 106820 116448
rect 106884 116384 106900 116448
rect 106964 116384 106970 116448
rect 106654 116383 106970 116384
rect 4210 115904 4526 115905
rect 4210 115840 4216 115904
rect 4280 115840 4296 115904
rect 4360 115840 4376 115904
rect 4440 115840 4456 115904
rect 4520 115840 4526 115904
rect 4210 115839 4526 115840
rect 105918 115904 106234 115905
rect 105918 115840 105924 115904
rect 105988 115840 106004 115904
rect 106068 115840 106084 115904
rect 106148 115840 106164 115904
rect 106228 115840 106234 115904
rect 105918 115839 106234 115840
rect 4870 115360 5186 115361
rect 4870 115296 4876 115360
rect 4940 115296 4956 115360
rect 5020 115296 5036 115360
rect 5100 115296 5116 115360
rect 5180 115296 5186 115360
rect 4870 115295 5186 115296
rect 106654 115360 106970 115361
rect 106654 115296 106660 115360
rect 106724 115296 106740 115360
rect 106804 115296 106820 115360
rect 106884 115296 106900 115360
rect 106964 115296 106970 115360
rect 106654 115295 106970 115296
rect 4210 114816 4526 114817
rect 4210 114752 4216 114816
rect 4280 114752 4296 114816
rect 4360 114752 4376 114816
rect 4440 114752 4456 114816
rect 4520 114752 4526 114816
rect 4210 114751 4526 114752
rect 105918 114816 106234 114817
rect 105918 114752 105924 114816
rect 105988 114752 106004 114816
rect 106068 114752 106084 114816
rect 106148 114752 106164 114816
rect 106228 114752 106234 114816
rect 105918 114751 106234 114752
rect 4870 114272 5186 114273
rect 4870 114208 4876 114272
rect 4940 114208 4956 114272
rect 5020 114208 5036 114272
rect 5100 114208 5116 114272
rect 5180 114208 5186 114272
rect 4870 114207 5186 114208
rect 106654 114272 106970 114273
rect 106654 114208 106660 114272
rect 106724 114208 106740 114272
rect 106804 114208 106820 114272
rect 106884 114208 106900 114272
rect 106964 114208 106970 114272
rect 106654 114207 106970 114208
rect 4210 113728 4526 113729
rect 4210 113664 4216 113728
rect 4280 113664 4296 113728
rect 4360 113664 4376 113728
rect 4440 113664 4456 113728
rect 4520 113664 4526 113728
rect 4210 113663 4526 113664
rect 105918 113728 106234 113729
rect 105918 113664 105924 113728
rect 105988 113664 106004 113728
rect 106068 113664 106084 113728
rect 106148 113664 106164 113728
rect 106228 113664 106234 113728
rect 105918 113663 106234 113664
rect 4870 113184 5186 113185
rect 4870 113120 4876 113184
rect 4940 113120 4956 113184
rect 5020 113120 5036 113184
rect 5100 113120 5116 113184
rect 5180 113120 5186 113184
rect 4870 113119 5186 113120
rect 106654 113184 106970 113185
rect 106654 113120 106660 113184
rect 106724 113120 106740 113184
rect 106804 113120 106820 113184
rect 106884 113120 106900 113184
rect 106964 113120 106970 113184
rect 106654 113119 106970 113120
rect 4210 112640 4526 112641
rect 4210 112576 4216 112640
rect 4280 112576 4296 112640
rect 4360 112576 4376 112640
rect 4440 112576 4456 112640
rect 4520 112576 4526 112640
rect 4210 112575 4526 112576
rect 105918 112640 106234 112641
rect 105918 112576 105924 112640
rect 105988 112576 106004 112640
rect 106068 112576 106084 112640
rect 106148 112576 106164 112640
rect 106228 112576 106234 112640
rect 105918 112575 106234 112576
rect 4870 112096 5186 112097
rect 4870 112032 4876 112096
rect 4940 112032 4956 112096
rect 5020 112032 5036 112096
rect 5100 112032 5116 112096
rect 5180 112032 5186 112096
rect 4870 112031 5186 112032
rect 106654 112096 106970 112097
rect 106654 112032 106660 112096
rect 106724 112032 106740 112096
rect 106804 112032 106820 112096
rect 106884 112032 106900 112096
rect 106964 112032 106970 112096
rect 106654 112031 106970 112032
rect 4210 111552 4526 111553
rect 4210 111488 4216 111552
rect 4280 111488 4296 111552
rect 4360 111488 4376 111552
rect 4440 111488 4456 111552
rect 4520 111488 4526 111552
rect 4210 111487 4526 111488
rect 105918 111552 106234 111553
rect 105918 111488 105924 111552
rect 105988 111488 106004 111552
rect 106068 111488 106084 111552
rect 106148 111488 106164 111552
rect 106228 111488 106234 111552
rect 105918 111487 106234 111488
rect 8385 111210 8451 111213
rect 9446 111210 10028 111254
rect 8385 111208 10028 111210
rect 8385 111152 8390 111208
rect 8446 111194 10028 111208
rect 8446 111152 9506 111194
rect 8385 111150 9506 111152
rect 8385 111147 8451 111150
rect 4870 111008 5186 111009
rect 0 110938 800 110968
rect 4870 110944 4876 111008
rect 4940 110944 4956 111008
rect 5020 110944 5036 111008
rect 5100 110944 5116 111008
rect 5180 110944 5186 111008
rect 4870 110943 5186 110944
rect 106654 111008 106970 111009
rect 106654 110944 106660 111008
rect 106724 110944 106740 111008
rect 106804 110944 106820 111008
rect 106884 110944 106900 111008
rect 106964 110944 106970 111008
rect 106654 110943 106970 110944
rect 1301 110938 1367 110941
rect 0 110936 1367 110938
rect 0 110880 1306 110936
rect 1362 110880 1367 110936
rect 0 110878 1367 110880
rect 0 110848 800 110878
rect 1301 110875 1367 110878
rect 4210 110464 4526 110465
rect 4210 110400 4216 110464
rect 4280 110400 4296 110464
rect 4360 110400 4376 110464
rect 4440 110400 4456 110464
rect 4520 110400 4526 110464
rect 4210 110399 4526 110400
rect 105918 110464 106234 110465
rect 105918 110400 105924 110464
rect 105988 110400 106004 110464
rect 106068 110400 106084 110464
rect 106148 110400 106164 110464
rect 106228 110400 106234 110464
rect 105918 110399 106234 110400
rect 4870 109920 5186 109921
rect 4870 109856 4876 109920
rect 4940 109856 4956 109920
rect 5020 109856 5036 109920
rect 5100 109856 5116 109920
rect 5180 109856 5186 109920
rect 4870 109855 5186 109856
rect 106654 109920 106970 109921
rect 106654 109856 106660 109920
rect 106724 109856 106740 109920
rect 106804 109856 106820 109920
rect 106884 109856 106900 109920
rect 106964 109856 106970 109920
rect 106654 109855 106970 109856
rect 0 109578 800 109608
rect 1301 109578 1367 109581
rect 0 109576 1367 109578
rect 0 109520 1306 109576
rect 1362 109520 1367 109576
rect 0 109518 1367 109520
rect 0 109488 800 109518
rect 1301 109515 1367 109518
rect 8385 109578 8451 109581
rect 8385 109576 9506 109578
rect 8385 109520 8390 109576
rect 8446 109554 9506 109576
rect 8446 109520 10028 109554
rect 8385 109518 10028 109520
rect 8385 109515 8451 109518
rect 9446 109494 10028 109518
rect 4210 109376 4526 109377
rect 4210 109312 4216 109376
rect 4280 109312 4296 109376
rect 4360 109312 4376 109376
rect 4440 109312 4456 109376
rect 4520 109312 4526 109376
rect 4210 109311 4526 109312
rect 105918 109376 106234 109377
rect 105918 109312 105924 109376
rect 105988 109312 106004 109376
rect 106068 109312 106084 109376
rect 106148 109312 106164 109376
rect 106228 109312 106234 109376
rect 105918 109311 106234 109312
rect 4870 108832 5186 108833
rect 4870 108768 4876 108832
rect 4940 108768 4956 108832
rect 5020 108768 5036 108832
rect 5100 108768 5116 108832
rect 5180 108768 5186 108832
rect 4870 108767 5186 108768
rect 106654 108832 106970 108833
rect 106654 108768 106660 108832
rect 106724 108768 106740 108832
rect 106804 108768 106820 108832
rect 106884 108768 106900 108832
rect 106964 108768 106970 108832
rect 106654 108767 106970 108768
rect 8385 108490 8451 108493
rect 8385 108488 9506 108490
rect 8385 108432 8390 108488
rect 8446 108432 9506 108488
rect 8385 108430 9506 108432
rect 8385 108427 8451 108430
rect 9446 108426 9506 108430
rect 9446 108366 10028 108426
rect 4210 108288 4526 108289
rect 0 108218 800 108248
rect 4210 108224 4216 108288
rect 4280 108224 4296 108288
rect 4360 108224 4376 108288
rect 4440 108224 4456 108288
rect 4520 108224 4526 108288
rect 4210 108223 4526 108224
rect 105918 108288 106234 108289
rect 105918 108224 105924 108288
rect 105988 108224 106004 108288
rect 106068 108224 106084 108288
rect 106148 108224 106164 108288
rect 106228 108224 106234 108288
rect 105918 108223 106234 108224
rect 1301 108218 1367 108221
rect 0 108216 1367 108218
rect 0 108160 1306 108216
rect 1362 108160 1367 108216
rect 0 108158 1367 108160
rect 0 108128 800 108158
rect 1301 108155 1367 108158
rect 4870 107744 5186 107745
rect 4870 107680 4876 107744
rect 4940 107680 4956 107744
rect 5020 107680 5036 107744
rect 5100 107680 5116 107744
rect 5180 107680 5186 107744
rect 4870 107679 5186 107680
rect 106654 107744 106970 107745
rect 106654 107680 106660 107744
rect 106724 107680 106740 107744
rect 106804 107680 106820 107744
rect 106884 107680 106900 107744
rect 106964 107680 106970 107744
rect 106654 107679 106970 107680
rect 4210 107200 4526 107201
rect 4210 107136 4216 107200
rect 4280 107136 4296 107200
rect 4360 107136 4376 107200
rect 4440 107136 4456 107200
rect 4520 107136 4526 107200
rect 4210 107135 4526 107136
rect 105918 107200 106234 107201
rect 105918 107136 105924 107200
rect 105988 107136 106004 107200
rect 106068 107136 106084 107200
rect 106148 107136 106164 107200
rect 106228 107136 106234 107200
rect 105918 107135 106234 107136
rect 0 106858 800 106888
rect 1209 106858 1275 106861
rect 0 106856 1275 106858
rect 0 106800 1214 106856
rect 1270 106800 1275 106856
rect 0 106798 1275 106800
rect 0 106768 800 106798
rect 1209 106795 1275 106798
rect 8385 106722 8451 106725
rect 9446 106722 10028 106726
rect 8385 106720 10028 106722
rect 8385 106664 8390 106720
rect 8446 106666 10028 106720
rect 8446 106664 9506 106666
rect 8385 106662 9506 106664
rect 8385 106659 8451 106662
rect 4870 106656 5186 106657
rect 4870 106592 4876 106656
rect 4940 106592 4956 106656
rect 5020 106592 5036 106656
rect 5100 106592 5116 106656
rect 5180 106592 5186 106656
rect 4870 106591 5186 106592
rect 106654 106656 106970 106657
rect 106654 106592 106660 106656
rect 106724 106592 106740 106656
rect 106804 106592 106820 106656
rect 106884 106592 106900 106656
rect 106964 106592 106970 106656
rect 106654 106591 106970 106592
rect 4210 106112 4526 106113
rect 4210 106048 4216 106112
rect 4280 106048 4296 106112
rect 4360 106048 4376 106112
rect 4440 106048 4456 106112
rect 4520 106048 4526 106112
rect 4210 106047 4526 106048
rect 105918 106112 106234 106113
rect 105918 106048 105924 106112
rect 105988 106048 106004 106112
rect 106068 106048 106084 106112
rect 106148 106048 106164 106112
rect 106228 106048 106234 106112
rect 105918 106047 106234 106048
rect 8385 105634 8451 105637
rect 9446 105634 10028 105643
rect 8385 105632 10028 105634
rect 8385 105576 8390 105632
rect 8446 105583 10028 105632
rect 8446 105576 9506 105583
rect 8385 105574 9506 105576
rect 8385 105571 8451 105574
rect 4870 105568 5186 105569
rect 0 105498 800 105528
rect 4870 105504 4876 105568
rect 4940 105504 4956 105568
rect 5020 105504 5036 105568
rect 5100 105504 5116 105568
rect 5180 105504 5186 105568
rect 4870 105503 5186 105504
rect 106654 105568 106970 105569
rect 106654 105504 106660 105568
rect 106724 105504 106740 105568
rect 106804 105504 106820 105568
rect 106884 105504 106900 105568
rect 106964 105504 106970 105568
rect 106654 105503 106970 105504
rect 1301 105498 1367 105501
rect 0 105496 1367 105498
rect 0 105440 1306 105496
rect 1362 105440 1367 105496
rect 0 105438 1367 105440
rect 0 105408 800 105438
rect 1301 105435 1367 105438
rect 4210 105024 4526 105025
rect 4210 104960 4216 105024
rect 4280 104960 4296 105024
rect 4360 104960 4376 105024
rect 4440 104960 4456 105024
rect 4520 104960 4526 105024
rect 4210 104959 4526 104960
rect 105918 105024 106234 105025
rect 105918 104960 105924 105024
rect 105988 104960 106004 105024
rect 106068 104960 106084 105024
rect 106148 104960 106164 105024
rect 106228 104960 106234 105024
rect 105918 104959 106234 104960
rect 4870 104480 5186 104481
rect 4870 104416 4876 104480
rect 4940 104416 4956 104480
rect 5020 104416 5036 104480
rect 5100 104416 5116 104480
rect 5180 104416 5186 104480
rect 4870 104415 5186 104416
rect 106654 104480 106970 104481
rect 106654 104416 106660 104480
rect 106724 104416 106740 104480
rect 106804 104416 106820 104480
rect 106884 104416 106900 104480
rect 106964 104416 106970 104480
rect 106654 104415 106970 104416
rect 0 104138 800 104168
rect 1301 104138 1367 104141
rect 0 104136 1367 104138
rect 0 104080 1306 104136
rect 1362 104080 1367 104136
rect 0 104078 1367 104080
rect 0 104048 800 104078
rect 1301 104075 1367 104078
rect 8385 104002 8451 104005
rect 8385 104000 9506 104002
rect 8385 103944 8390 104000
rect 8446 103963 9506 104000
rect 8446 103944 10028 103963
rect 8385 103942 10028 103944
rect 8385 103939 8451 103942
rect 4210 103936 4526 103937
rect 4210 103872 4216 103936
rect 4280 103872 4296 103936
rect 4360 103872 4376 103936
rect 4440 103872 4456 103936
rect 4520 103872 4526 103936
rect 9446 103903 10028 103942
rect 105918 103936 106234 103937
rect 4210 103871 4526 103872
rect 105918 103872 105924 103936
rect 105988 103872 106004 103936
rect 106068 103872 106084 103936
rect 106148 103872 106164 103936
rect 106228 103872 106234 103936
rect 105918 103871 106234 103872
rect 4870 103392 5186 103393
rect 4870 103328 4876 103392
rect 4940 103328 4956 103392
rect 5020 103328 5036 103392
rect 5100 103328 5116 103392
rect 5180 103328 5186 103392
rect 4870 103327 5186 103328
rect 106654 103392 106970 103393
rect 106654 103328 106660 103392
rect 106724 103328 106740 103392
rect 106804 103328 106820 103392
rect 106884 103328 106900 103392
rect 106964 103328 106970 103392
rect 106654 103327 106970 103328
rect 4210 102848 4526 102849
rect 4210 102784 4216 102848
rect 4280 102784 4296 102848
rect 4360 102784 4376 102848
rect 4440 102784 4456 102848
rect 4520 102784 4526 102848
rect 4210 102783 4526 102784
rect 105918 102848 106234 102849
rect 105918 102784 105924 102848
rect 105988 102784 106004 102848
rect 106068 102784 106084 102848
rect 106148 102784 106164 102848
rect 106228 102784 106234 102848
rect 105918 102783 106234 102784
rect 4870 102304 5186 102305
rect 4870 102240 4876 102304
rect 4940 102240 4956 102304
rect 5020 102240 5036 102304
rect 5100 102240 5116 102304
rect 5180 102240 5186 102304
rect 4870 102239 5186 102240
rect 106654 102304 106970 102305
rect 106654 102240 106660 102304
rect 106724 102240 106740 102304
rect 106804 102240 106820 102304
rect 106884 102240 106900 102304
rect 106964 102240 106970 102304
rect 106654 102239 106970 102240
rect 4210 101760 4526 101761
rect 4210 101696 4216 101760
rect 4280 101696 4296 101760
rect 4360 101696 4376 101760
rect 4440 101696 4456 101760
rect 4520 101696 4526 101760
rect 4210 101695 4526 101696
rect 105918 101760 106234 101761
rect 105918 101696 105924 101760
rect 105988 101696 106004 101760
rect 106068 101696 106084 101760
rect 106148 101696 106164 101760
rect 106228 101696 106234 101760
rect 105918 101695 106234 101696
rect 4870 101216 5186 101217
rect 4870 101152 4876 101216
rect 4940 101152 4956 101216
rect 5020 101152 5036 101216
rect 5100 101152 5116 101216
rect 5180 101152 5186 101216
rect 4870 101151 5186 101152
rect 106654 101216 106970 101217
rect 106654 101152 106660 101216
rect 106724 101152 106740 101216
rect 106804 101152 106820 101216
rect 106884 101152 106900 101216
rect 106964 101152 106970 101216
rect 106654 101151 106970 101152
rect 4210 100672 4526 100673
rect 4210 100608 4216 100672
rect 4280 100608 4296 100672
rect 4360 100608 4376 100672
rect 4440 100608 4456 100672
rect 4520 100608 4526 100672
rect 4210 100607 4526 100608
rect 105918 100672 106234 100673
rect 105918 100608 105924 100672
rect 105988 100608 106004 100672
rect 106068 100608 106084 100672
rect 106148 100608 106164 100672
rect 106228 100608 106234 100672
rect 105918 100607 106234 100608
rect 4870 100128 5186 100129
rect 4870 100064 4876 100128
rect 4940 100064 4956 100128
rect 5020 100064 5036 100128
rect 5100 100064 5116 100128
rect 5180 100064 5186 100128
rect 4870 100063 5186 100064
rect 106654 100128 106970 100129
rect 106654 100064 106660 100128
rect 106724 100064 106740 100128
rect 106804 100064 106820 100128
rect 106884 100064 106900 100128
rect 106964 100064 106970 100128
rect 106654 100063 106970 100064
rect 4210 99584 4526 99585
rect 4210 99520 4216 99584
rect 4280 99520 4296 99584
rect 4360 99520 4376 99584
rect 4440 99520 4456 99584
rect 4520 99520 4526 99584
rect 4210 99519 4526 99520
rect 105918 99584 106234 99585
rect 105918 99520 105924 99584
rect 105988 99520 106004 99584
rect 106068 99520 106084 99584
rect 106148 99520 106164 99584
rect 106228 99520 106234 99584
rect 105918 99519 106234 99520
rect 4870 99040 5186 99041
rect 4870 98976 4876 99040
rect 4940 98976 4956 99040
rect 5020 98976 5036 99040
rect 5100 98976 5116 99040
rect 5180 98976 5186 99040
rect 4870 98975 5186 98976
rect 106654 99040 106970 99041
rect 106654 98976 106660 99040
rect 106724 98976 106740 99040
rect 106804 98976 106820 99040
rect 106884 98976 106900 99040
rect 106964 98976 106970 99040
rect 106654 98975 106970 98976
rect 4210 98496 4526 98497
rect 4210 98432 4216 98496
rect 4280 98432 4296 98496
rect 4360 98432 4376 98496
rect 4440 98432 4456 98496
rect 4520 98432 4526 98496
rect 4210 98431 4526 98432
rect 105918 98496 106234 98497
rect 105918 98432 105924 98496
rect 105988 98432 106004 98496
rect 106068 98432 106084 98496
rect 106148 98432 106164 98496
rect 106228 98432 106234 98496
rect 105918 98431 106234 98432
rect 4870 97952 5186 97953
rect 4870 97888 4876 97952
rect 4940 97888 4956 97952
rect 5020 97888 5036 97952
rect 5100 97888 5116 97952
rect 5180 97888 5186 97952
rect 4870 97887 5186 97888
rect 106654 97952 106970 97953
rect 106654 97888 106660 97952
rect 106724 97888 106740 97952
rect 106804 97888 106820 97952
rect 106884 97888 106900 97952
rect 106964 97888 106970 97952
rect 106654 97887 106970 97888
rect 4210 97408 4526 97409
rect 4210 97344 4216 97408
rect 4280 97344 4296 97408
rect 4360 97344 4376 97408
rect 4440 97344 4456 97408
rect 4520 97344 4526 97408
rect 4210 97343 4526 97344
rect 105918 97408 106234 97409
rect 105918 97344 105924 97408
rect 105988 97344 106004 97408
rect 106068 97344 106084 97408
rect 106148 97344 106164 97408
rect 106228 97344 106234 97408
rect 105918 97343 106234 97344
rect 4870 96864 5186 96865
rect 4870 96800 4876 96864
rect 4940 96800 4956 96864
rect 5020 96800 5036 96864
rect 5100 96800 5116 96864
rect 5180 96800 5186 96864
rect 4870 96799 5186 96800
rect 106654 96864 106970 96865
rect 106654 96800 106660 96864
rect 106724 96800 106740 96864
rect 106804 96800 106820 96864
rect 106884 96800 106900 96864
rect 106964 96800 106970 96864
rect 106654 96799 106970 96800
rect 4210 96320 4526 96321
rect 4210 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4526 96320
rect 4210 96255 4526 96256
rect 105918 96320 106234 96321
rect 105918 96256 105924 96320
rect 105988 96256 106004 96320
rect 106068 96256 106084 96320
rect 106148 96256 106164 96320
rect 106228 96256 106234 96320
rect 105918 96255 106234 96256
rect 4870 95776 5186 95777
rect 4870 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5186 95776
rect 4870 95711 5186 95712
rect 106654 95776 106970 95777
rect 106654 95712 106660 95776
rect 106724 95712 106740 95776
rect 106804 95712 106820 95776
rect 106884 95712 106900 95776
rect 106964 95712 106970 95776
rect 106654 95711 106970 95712
rect 4210 95232 4526 95233
rect 4210 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4526 95232
rect 4210 95167 4526 95168
rect 105918 95232 106234 95233
rect 105918 95168 105924 95232
rect 105988 95168 106004 95232
rect 106068 95168 106084 95232
rect 106148 95168 106164 95232
rect 106228 95168 106234 95232
rect 105918 95167 106234 95168
rect 101948 95030 102242 95090
rect 102182 95026 102242 95030
rect 102685 95026 102751 95029
rect 102182 95024 102751 95026
rect 102182 94968 102690 95024
rect 102746 94968 102751 95024
rect 102182 94966 102751 94968
rect 102685 94963 102751 94966
rect 4870 94688 5186 94689
rect 4870 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5186 94688
rect 4870 94623 5186 94624
rect 106654 94688 106970 94689
rect 106654 94624 106660 94688
rect 106724 94624 106740 94688
rect 106804 94624 106820 94688
rect 106884 94624 106900 94688
rect 106964 94624 106970 94688
rect 106654 94623 106970 94624
rect 4210 94144 4526 94145
rect 4210 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4526 94144
rect 4210 94079 4526 94080
rect 105918 94144 106234 94145
rect 105918 94080 105924 94144
rect 105988 94080 106004 94144
rect 106068 94080 106084 94144
rect 106148 94080 106164 94144
rect 106228 94080 106234 94144
rect 105918 94079 106234 94080
rect 4870 93600 5186 93601
rect 4870 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5186 93600
rect 4870 93535 5186 93536
rect 106654 93600 106970 93601
rect 106654 93536 106660 93600
rect 106724 93536 106740 93600
rect 106804 93536 106820 93600
rect 106884 93536 106900 93600
rect 106964 93536 106970 93600
rect 106654 93535 106970 93536
rect 102869 93394 102935 93397
rect 102550 93392 102935 93394
rect 102550 93390 102874 93392
rect 101948 93336 102874 93390
rect 102930 93336 102935 93392
rect 101948 93334 102935 93336
rect 101948 93330 102610 93334
rect 102869 93331 102935 93334
rect 4210 93056 4526 93057
rect 4210 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4526 93056
rect 4210 92991 4526 92992
rect 105918 93056 106234 93057
rect 105918 92992 105924 93056
rect 105988 92992 106004 93056
rect 106068 92992 106084 93056
rect 106148 92992 106164 93056
rect 106228 92992 106234 93056
rect 105918 92991 106234 92992
rect 4870 92512 5186 92513
rect 4870 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5186 92512
rect 4870 92447 5186 92448
rect 106654 92512 106970 92513
rect 106654 92448 106660 92512
rect 106724 92448 106740 92512
rect 106804 92448 106820 92512
rect 106884 92448 106900 92512
rect 106964 92448 106970 92512
rect 106654 92447 106970 92448
rect 102961 92306 103027 92309
rect 102550 92304 103027 92306
rect 102550 92262 102966 92304
rect 101948 92248 102966 92262
rect 103022 92248 103027 92304
rect 101948 92246 103027 92248
rect 101948 92202 102610 92246
rect 102961 92243 103027 92246
rect 4210 91968 4526 91969
rect 4210 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4526 91968
rect 4210 91903 4526 91904
rect 105918 91968 106234 91969
rect 105918 91904 105924 91968
rect 105988 91904 106004 91968
rect 106068 91904 106084 91968
rect 106148 91904 106164 91968
rect 106228 91904 106234 91968
rect 105918 91903 106234 91904
rect 4870 91424 5186 91425
rect 4870 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5186 91424
rect 4870 91359 5186 91360
rect 106654 91424 106970 91425
rect 106654 91360 106660 91424
rect 106724 91360 106740 91424
rect 106804 91360 106820 91424
rect 106884 91360 106900 91424
rect 106964 91360 106970 91424
rect 106654 91359 106970 91360
rect 4210 90880 4526 90881
rect 4210 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4526 90880
rect 4210 90815 4526 90816
rect 105918 90880 106234 90881
rect 105918 90816 105924 90880
rect 105988 90816 106004 90880
rect 106068 90816 106084 90880
rect 106148 90816 106164 90880
rect 106228 90816 106234 90880
rect 105918 90815 106234 90816
rect 4870 90336 5186 90337
rect 4870 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5186 90336
rect 4870 90271 5186 90272
rect 106654 90336 106970 90337
rect 106654 90272 106660 90336
rect 106724 90272 106740 90336
rect 106804 90272 106820 90336
rect 106884 90272 106900 90336
rect 106964 90272 106970 90336
rect 106654 90271 106970 90272
rect 4210 89792 4526 89793
rect 4210 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4526 89792
rect 4210 89727 4526 89728
rect 105918 89792 106234 89793
rect 105918 89728 105924 89792
rect 105988 89728 106004 89792
rect 106068 89728 106084 89792
rect 106148 89728 106164 89792
rect 106228 89728 106234 89792
rect 105918 89727 106234 89728
rect 4870 89248 5186 89249
rect 4870 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5186 89248
rect 4870 89183 5186 89184
rect 106654 89248 106970 89249
rect 106654 89184 106660 89248
rect 106724 89184 106740 89248
rect 106804 89184 106820 89248
rect 106884 89184 106900 89248
rect 106964 89184 106970 89248
rect 106654 89183 106970 89184
rect 4210 88704 4526 88705
rect 4210 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4526 88704
rect 4210 88639 4526 88640
rect 105918 88704 106234 88705
rect 105918 88640 105924 88704
rect 105988 88640 106004 88704
rect 106068 88640 106084 88704
rect 106148 88640 106164 88704
rect 106228 88640 106234 88704
rect 105918 88639 106234 88640
rect 0 88498 800 88528
rect 1301 88498 1367 88501
rect 0 88496 1367 88498
rect 0 88440 1306 88496
rect 1362 88440 1367 88496
rect 0 88438 1367 88440
rect 0 88408 800 88438
rect 1301 88435 1367 88438
rect 4870 88160 5186 88161
rect 4870 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5186 88160
rect 4870 88095 5186 88096
rect 106654 88160 106970 88161
rect 106654 88096 106660 88160
rect 106724 88096 106740 88160
rect 106804 88096 106820 88160
rect 106884 88096 106900 88160
rect 106964 88096 106970 88160
rect 106654 88095 106970 88096
rect 0 87818 800 87848
rect 1209 87818 1275 87821
rect 0 87816 1275 87818
rect 0 87760 1214 87816
rect 1270 87760 1275 87816
rect 0 87758 1275 87760
rect 0 87728 800 87758
rect 1209 87755 1275 87758
rect 4210 87616 4526 87617
rect 4210 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4526 87616
rect 4210 87551 4526 87552
rect 105918 87616 106234 87617
rect 105918 87552 105924 87616
rect 105988 87552 106004 87616
rect 106068 87552 106084 87616
rect 106148 87552 106164 87616
rect 106228 87552 106234 87616
rect 105918 87551 106234 87552
rect 0 87138 800 87168
rect 1209 87138 1275 87141
rect 0 87136 1275 87138
rect 0 87080 1214 87136
rect 1270 87080 1275 87136
rect 0 87078 1275 87080
rect 0 87048 800 87078
rect 1209 87075 1275 87078
rect 4870 87072 5186 87073
rect 4870 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5186 87072
rect 4870 87007 5186 87008
rect 106654 87072 106970 87073
rect 106654 87008 106660 87072
rect 106724 87008 106740 87072
rect 106804 87008 106820 87072
rect 106884 87008 106900 87072
rect 106964 87008 106970 87072
rect 106654 87007 106970 87008
rect 4210 86528 4526 86529
rect 0 86458 800 86488
rect 4210 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4526 86528
rect 4210 86463 4526 86464
rect 105918 86528 106234 86529
rect 105918 86464 105924 86528
rect 105988 86464 106004 86528
rect 106068 86464 106084 86528
rect 106148 86464 106164 86528
rect 106228 86464 106234 86528
rect 105918 86463 106234 86464
rect 1301 86458 1367 86461
rect 0 86456 1367 86458
rect 0 86400 1306 86456
rect 1362 86400 1367 86456
rect 0 86398 1367 86400
rect 0 86368 800 86398
rect 1301 86395 1367 86398
rect 4870 85984 5186 85985
rect 4870 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5186 85984
rect 4870 85919 5186 85920
rect 106654 85984 106970 85985
rect 106654 85920 106660 85984
rect 106724 85920 106740 85984
rect 106804 85920 106820 85984
rect 106884 85920 106900 85984
rect 106964 85920 106970 85984
rect 106654 85919 106970 85920
rect 0 85778 800 85808
rect 1301 85778 1367 85781
rect 0 85776 1367 85778
rect 0 85720 1306 85776
rect 1362 85720 1367 85776
rect 0 85718 1367 85720
rect 0 85688 800 85718
rect 1301 85715 1367 85718
rect 5993 85506 6059 85509
rect 5993 85504 9506 85506
rect 5993 85448 5998 85504
rect 6054 85483 9506 85504
rect 6054 85448 10028 85483
rect 5993 85446 10028 85448
rect 5993 85443 6059 85446
rect 4210 85440 4526 85441
rect 4210 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4526 85440
rect 9446 85423 10028 85446
rect 105918 85440 106234 85441
rect 4210 85375 4526 85376
rect 105918 85376 105924 85440
rect 105988 85376 106004 85440
rect 106068 85376 106084 85440
rect 106148 85376 106164 85440
rect 106228 85376 106234 85440
rect 105918 85375 106234 85376
rect 0 85098 800 85128
rect 1209 85098 1275 85101
rect 0 85096 1275 85098
rect 0 85040 1214 85096
rect 1270 85040 1275 85096
rect 0 85038 1275 85040
rect 0 85008 800 85038
rect 1209 85035 1275 85038
rect 4870 84896 5186 84897
rect 4870 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5186 84896
rect 4870 84831 5186 84832
rect 106654 84896 106970 84897
rect 106654 84832 106660 84896
rect 106724 84832 106740 84896
rect 106804 84832 106820 84896
rect 106884 84832 106900 84896
rect 106964 84832 106970 84896
rect 106654 84831 106970 84832
rect 0 84418 800 84448
rect 1301 84418 1367 84421
rect 0 84416 1367 84418
rect 0 84360 1306 84416
rect 1362 84360 1367 84416
rect 0 84358 1367 84360
rect 0 84328 800 84358
rect 1301 84355 1367 84358
rect 4210 84352 4526 84353
rect 4210 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4526 84352
rect 4210 84287 4526 84288
rect 105918 84352 106234 84353
rect 105918 84288 105924 84352
rect 105988 84288 106004 84352
rect 106068 84288 106084 84352
rect 106148 84288 106164 84352
rect 106228 84288 106234 84352
rect 105918 84287 106234 84288
rect 4870 83808 5186 83809
rect 0 83738 800 83768
rect 4870 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5186 83808
rect 4870 83743 5186 83744
rect 106654 83808 106970 83809
rect 106654 83744 106660 83808
rect 106724 83744 106740 83808
rect 106804 83744 106820 83808
rect 106884 83744 106900 83808
rect 106964 83744 106970 83808
rect 106654 83743 106970 83744
rect 1301 83738 1367 83741
rect 0 83736 1367 83738
rect 0 83680 1306 83736
rect 1362 83680 1367 83736
rect 0 83678 1367 83680
rect 0 83648 800 83678
rect 1301 83675 1367 83678
rect 4210 83264 4526 83265
rect 4210 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4526 83264
rect 4210 83199 4526 83200
rect 105918 83264 106234 83265
rect 105918 83200 105924 83264
rect 105988 83200 106004 83264
rect 106068 83200 106084 83264
rect 106148 83200 106164 83264
rect 106228 83200 106234 83264
rect 105918 83199 106234 83200
rect 0 83058 800 83088
rect 1301 83058 1367 83061
rect 0 83056 1367 83058
rect 0 83000 1306 83056
rect 1362 83000 1367 83056
rect 0 82998 1367 83000
rect 0 82968 800 82998
rect 1301 82995 1367 82998
rect 4870 82720 5186 82721
rect 4870 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5186 82720
rect 4870 82655 5186 82656
rect 106654 82720 106970 82721
rect 106654 82656 106660 82720
rect 106724 82656 106740 82720
rect 106804 82656 106820 82720
rect 106884 82656 106900 82720
rect 106964 82656 106970 82720
rect 106654 82655 106970 82656
rect 0 82378 800 82408
rect 1209 82378 1275 82381
rect 0 82376 1275 82378
rect 0 82320 1214 82376
rect 1270 82320 1275 82376
rect 0 82318 1275 82320
rect 0 82288 800 82318
rect 1209 82315 1275 82318
rect 4210 82176 4526 82177
rect 4210 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4526 82176
rect 4210 82111 4526 82112
rect 105918 82176 106234 82177
rect 105918 82112 105924 82176
rect 105988 82112 106004 82176
rect 106068 82112 106084 82176
rect 106148 82112 106164 82176
rect 106228 82112 106234 82176
rect 105918 82111 106234 82112
rect 0 81698 800 81728
rect 1209 81698 1275 81701
rect 0 81696 1275 81698
rect 0 81640 1214 81696
rect 1270 81640 1275 81696
rect 0 81638 1275 81640
rect 0 81608 800 81638
rect 1209 81635 1275 81638
rect 4870 81632 5186 81633
rect 4870 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5186 81632
rect 4870 81567 5186 81568
rect 106654 81632 106970 81633
rect 106654 81568 106660 81632
rect 106724 81568 106740 81632
rect 106804 81568 106820 81632
rect 106884 81568 106900 81632
rect 106964 81568 106970 81632
rect 106654 81567 106970 81568
rect 4210 81088 4526 81089
rect 0 81018 800 81048
rect 4210 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4526 81088
rect 4210 81023 4526 81024
rect 105918 81088 106234 81089
rect 105918 81024 105924 81088
rect 105988 81024 106004 81088
rect 106068 81024 106084 81088
rect 106148 81024 106164 81088
rect 106228 81024 106234 81088
rect 105918 81023 106234 81024
rect 1301 81018 1367 81021
rect 0 81016 1367 81018
rect 0 80960 1306 81016
rect 1362 80960 1367 81016
rect 0 80958 1367 80960
rect 0 80928 800 80958
rect 1301 80955 1367 80958
rect 4870 80544 5186 80545
rect 4870 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5186 80544
rect 4870 80479 5186 80480
rect 106654 80544 106970 80545
rect 106654 80480 106660 80544
rect 106724 80480 106740 80544
rect 106804 80480 106820 80544
rect 106884 80480 106900 80544
rect 106964 80480 106970 80544
rect 106654 80479 106970 80480
rect 0 80338 800 80368
rect 1301 80338 1367 80341
rect 0 80336 1367 80338
rect 0 80280 1306 80336
rect 1362 80280 1367 80336
rect 0 80278 1367 80280
rect 0 80248 800 80278
rect 1301 80275 1367 80278
rect 4210 80000 4526 80001
rect 4210 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4526 80000
rect 4210 79935 4526 79936
rect 105918 80000 106234 80001
rect 105918 79936 105924 80000
rect 105988 79936 106004 80000
rect 106068 79936 106084 80000
rect 106148 79936 106164 80000
rect 106228 79936 106234 80000
rect 105918 79935 106234 79936
rect 8477 79930 8543 79933
rect 36261 79932 36327 79933
rect 38653 79932 38719 79933
rect 31608 79930 31614 79932
rect 8477 79928 31614 79930
rect 8477 79872 8482 79928
rect 8538 79872 31614 79928
rect 8477 79870 31614 79872
rect 8477 79867 8543 79870
rect 31608 79868 31614 79870
rect 31678 79868 31684 79932
rect 36261 79928 36286 79932
rect 36350 79930 36356 79932
rect 38616 79930 38622 79932
rect 36261 79872 36266 79928
rect 36261 79868 36286 79872
rect 36350 79870 36418 79930
rect 38562 79870 38622 79930
rect 38686 79928 38719 79932
rect 38714 79872 38719 79928
rect 36350 79868 36356 79870
rect 38616 79868 38622 79870
rect 38686 79868 38719 79872
rect 36261 79867 36327 79868
rect 38653 79867 38719 79868
rect 39757 79932 39823 79933
rect 40953 79932 41019 79933
rect 39757 79928 39790 79932
rect 39854 79930 39860 79932
rect 39757 79872 39762 79928
rect 39757 79868 39790 79872
rect 39854 79870 39914 79930
rect 39854 79868 39860 79870
rect 40952 79868 40958 79932
rect 41022 79930 41028 79932
rect 90633 79930 90699 79933
rect 90808 79930 90814 79932
rect 41022 79870 41110 79930
rect 90633 79928 90814 79930
rect 90633 79872 90638 79928
rect 90694 79872 90814 79928
rect 90633 79870 90814 79872
rect 41022 79868 41028 79870
rect 39757 79867 39823 79868
rect 40953 79867 41019 79868
rect 90633 79867 90699 79870
rect 90808 79868 90814 79870
rect 90878 79868 90884 79932
rect 8661 79794 8727 79797
rect 30440 79794 30446 79796
rect 8661 79792 30446 79794
rect 8661 79736 8666 79792
rect 8722 79736 30446 79792
rect 8661 79734 30446 79736
rect 8661 79731 8727 79734
rect 30440 79732 30446 79734
rect 30510 79732 30516 79796
rect 32305 79794 32371 79797
rect 32776 79794 32782 79796
rect 32305 79792 32782 79794
rect 32305 79736 32310 79792
rect 32366 79736 32782 79792
rect 32305 79734 32782 79736
rect 32305 79731 32371 79734
rect 32776 79732 32782 79734
rect 32846 79732 32852 79796
rect 0 79658 800 79688
rect 1209 79658 1275 79661
rect 0 79656 1275 79658
rect 0 79600 1214 79656
rect 1270 79600 1275 79656
rect 0 79598 1275 79600
rect 0 79568 800 79598
rect 1209 79595 1275 79598
rect 5625 79658 5691 79661
rect 25768 79658 25774 79660
rect 5625 79656 25774 79658
rect 5625 79600 5630 79656
rect 5686 79600 25774 79656
rect 5625 79598 25774 79600
rect 5625 79595 5691 79598
rect 25768 79596 25774 79598
rect 25838 79658 25844 79660
rect 27613 79658 27679 79661
rect 25838 79656 27679 79658
rect 25838 79600 27618 79656
rect 27674 79600 27679 79656
rect 25838 79598 27679 79600
rect 25838 79596 25844 79598
rect 27613 79595 27679 79598
rect 36997 79658 37063 79661
rect 37448 79658 37454 79660
rect 36997 79656 37454 79658
rect 36997 79600 37002 79656
rect 37058 79600 37454 79656
rect 36997 79598 37454 79600
rect 36997 79595 37063 79598
rect 37448 79596 37454 79598
rect 37518 79596 37524 79660
rect 5533 79522 5599 79525
rect 24669 79524 24735 79525
rect 24600 79522 24606 79524
rect 5533 79520 24606 79522
rect 5533 79464 5538 79520
rect 5594 79464 24606 79520
rect 5533 79462 24606 79464
rect 5533 79459 5599 79462
rect 24600 79460 24606 79462
rect 24670 79522 24735 79524
rect 24670 79520 24798 79522
rect 24670 79464 24674 79520
rect 24730 79464 24798 79520
rect 24670 79462 24798 79464
rect 24670 79460 24735 79462
rect 29272 79460 29278 79524
rect 29342 79522 29348 79524
rect 29545 79522 29611 79525
rect 30465 79524 30531 79525
rect 30440 79522 30446 79524
rect 29342 79520 29611 79522
rect 29342 79464 29550 79520
rect 29606 79464 29611 79520
rect 29342 79462 29611 79464
rect 30374 79462 30446 79522
rect 30510 79520 30531 79524
rect 30526 79464 30531 79520
rect 29342 79460 29348 79462
rect 24669 79459 24735 79460
rect 29545 79459 29611 79462
rect 30440 79460 30446 79462
rect 30510 79460 30531 79464
rect 30465 79459 30531 79460
rect 31569 79524 31635 79525
rect 33961 79524 34027 79525
rect 31569 79520 31614 79524
rect 31678 79522 31684 79524
rect 31569 79464 31574 79520
rect 31569 79460 31614 79464
rect 31678 79462 31726 79522
rect 31678 79460 31684 79462
rect 33944 79460 33950 79524
rect 34014 79522 34027 79524
rect 34697 79522 34763 79525
rect 42149 79524 42215 79525
rect 35106 79522 35112 79524
rect 34014 79520 34106 79522
rect 34022 79464 34106 79520
rect 34014 79462 34106 79464
rect 34697 79520 35112 79522
rect 34697 79464 34702 79520
rect 34758 79464 35112 79520
rect 34697 79462 35112 79464
rect 34014 79460 34027 79462
rect 31569 79459 31635 79460
rect 33961 79459 34027 79460
rect 34697 79459 34763 79462
rect 35106 79460 35112 79462
rect 35176 79460 35182 79524
rect 42120 79522 42126 79524
rect 42058 79462 42126 79522
rect 42190 79520 42215 79524
rect 42210 79464 42215 79520
rect 42120 79460 42126 79462
rect 42190 79460 42215 79464
rect 42149 79459 42215 79460
rect 43253 79524 43319 79525
rect 43253 79520 43294 79524
rect 43358 79522 43364 79524
rect 43253 79464 43258 79520
rect 43253 79460 43294 79464
rect 43358 79462 43410 79522
rect 43358 79460 43364 79462
rect 90674 79460 90680 79524
rect 90744 79522 90750 79524
rect 90909 79522 90975 79525
rect 90744 79520 90975 79522
rect 90744 79464 90914 79520
rect 90970 79464 90975 79520
rect 90744 79462 90975 79464
rect 90744 79460 90750 79462
rect 43253 79459 43319 79460
rect 90909 79459 90975 79462
rect 4870 79456 5186 79457
rect 4870 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5186 79456
rect 4870 79391 5186 79392
rect 106654 79456 106970 79457
rect 106654 79392 106660 79456
rect 106724 79392 106740 79456
rect 106804 79392 106820 79456
rect 106884 79392 106900 79456
rect 106964 79392 106970 79456
rect 106654 79391 106970 79392
rect 9397 79386 9463 79389
rect 26785 79386 26851 79389
rect 26918 79386 26924 79388
rect 9397 79384 26924 79386
rect 9397 79328 9402 79384
rect 9458 79328 26790 79384
rect 26846 79328 26924 79384
rect 9397 79326 26924 79328
rect 9397 79323 9463 79326
rect 26785 79323 26851 79326
rect 26918 79324 26924 79326
rect 26988 79324 26994 79388
rect 7557 79250 7623 79253
rect 23422 79250 23428 79252
rect 7557 79248 23428 79250
rect 7557 79192 7562 79248
rect 7618 79192 23428 79248
rect 7557 79190 23428 79192
rect 7557 79187 7623 79190
rect 23422 79188 23428 79190
rect 23492 79188 23498 79252
rect 0 78978 800 79008
rect 1301 78978 1367 78981
rect 0 78976 1367 78978
rect 0 78920 1306 78976
rect 1362 78920 1367 78976
rect 0 78918 1367 78920
rect 0 78888 800 78918
rect 1301 78915 1367 78918
rect 108481 78978 108547 78981
rect 109200 78978 110000 79008
rect 108481 78976 110000 78978
rect 108481 78920 108486 78976
rect 108542 78920 110000 78976
rect 108481 78918 110000 78920
rect 108481 78915 108547 78918
rect 4210 78912 4526 78913
rect 4210 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4526 78912
rect 4210 78847 4526 78848
rect 105918 78912 106234 78913
rect 105918 78848 105924 78912
rect 105988 78848 106004 78912
rect 106068 78848 106084 78912
rect 106148 78848 106164 78912
rect 106228 78848 106234 78912
rect 109200 78888 110000 78918
rect 105918 78847 106234 78848
rect 23422 78780 23428 78844
rect 23492 78842 23498 78844
rect 24761 78842 24827 78845
rect 23492 78840 24827 78842
rect 23492 78784 24766 78840
rect 24822 78784 24827 78840
rect 23492 78782 24827 78784
rect 23492 78780 23498 78782
rect 24761 78779 24827 78782
rect 8017 78570 8083 78573
rect 32949 78570 33015 78573
rect 8017 78568 33015 78570
rect 8017 78512 8022 78568
rect 8078 78512 32954 78568
rect 33010 78512 33015 78568
rect 8017 78510 33015 78512
rect 8017 78507 8083 78510
rect 32949 78507 33015 78510
rect 63309 78570 63375 78573
rect 96521 78570 96587 78573
rect 63309 78568 96587 78570
rect 63309 78512 63314 78568
rect 63370 78512 96526 78568
rect 96582 78512 96587 78568
rect 63309 78510 96587 78512
rect 63309 78507 63375 78510
rect 96521 78507 96587 78510
rect 78765 78434 78831 78437
rect 103881 78434 103947 78437
rect 78765 78432 103947 78434
rect 78765 78376 78770 78432
rect 78826 78376 103886 78432
rect 103942 78376 103947 78432
rect 78765 78374 103947 78376
rect 78765 78371 78831 78374
rect 103881 78371 103947 78374
rect 4870 78368 5186 78369
rect 0 78298 800 78328
rect 4870 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5186 78368
rect 4870 78303 5186 78304
rect 106654 78368 106970 78369
rect 106654 78304 106660 78368
rect 106724 78304 106740 78368
rect 106804 78304 106820 78368
rect 106884 78304 106900 78368
rect 106964 78304 106970 78368
rect 106654 78303 106970 78304
rect 1301 78298 1367 78301
rect 0 78296 1367 78298
rect 0 78240 1306 78296
rect 1362 78240 1367 78296
rect 0 78238 1367 78240
rect 0 78208 800 78238
rect 1301 78235 1367 78238
rect 9581 78298 9647 78301
rect 35341 78298 35407 78301
rect 9581 78296 35407 78298
rect 9581 78240 9586 78296
rect 9642 78240 35346 78296
rect 35402 78240 35407 78296
rect 9581 78238 35407 78240
rect 9581 78235 9647 78238
rect 35341 78235 35407 78238
rect 76189 78298 76255 78301
rect 102501 78298 102567 78301
rect 76189 78296 102567 78298
rect 76189 78240 76194 78296
rect 76250 78240 102506 78296
rect 102562 78240 102567 78296
rect 76189 78238 102567 78240
rect 76189 78235 76255 78238
rect 102501 78235 102567 78238
rect 108481 78298 108547 78301
rect 109200 78298 110000 78328
rect 108481 78296 110000 78298
rect 108481 78240 108486 78296
rect 108542 78240 110000 78296
rect 108481 78238 110000 78240
rect 108481 78235 108547 78238
rect 109200 78208 110000 78238
rect 8201 78162 8267 78165
rect 37733 78162 37799 78165
rect 8201 78160 37799 78162
rect 8201 78104 8206 78160
rect 8262 78104 37738 78160
rect 37794 78104 37799 78160
rect 8201 78102 37799 78104
rect 8201 78099 8267 78102
rect 37733 78099 37799 78102
rect 73981 78162 74047 78165
rect 103697 78162 103763 78165
rect 73981 78160 103763 78162
rect 73981 78104 73986 78160
rect 74042 78104 103702 78160
rect 103758 78104 103763 78160
rect 73981 78102 103763 78104
rect 73981 78099 74047 78102
rect 103697 78099 103763 78102
rect 16021 78028 16087 78029
rect 16021 78024 16068 78028
rect 16132 78026 16138 78028
rect 40125 78026 40191 78029
rect 40861 78026 40927 78029
rect 16021 77968 16026 78024
rect 16021 77964 16068 77968
rect 16132 77966 16178 78026
rect 16530 78024 40927 78026
rect 16530 77968 40130 78024
rect 40186 77968 40866 78024
rect 40922 77968 40927 78024
rect 16530 77966 40927 77968
rect 16132 77964 16138 77966
rect 16021 77963 16087 77964
rect 8109 77890 8175 77893
rect 16530 77890 16590 77966
rect 40125 77963 40191 77966
rect 40861 77963 40927 77966
rect 70945 78026 71011 78029
rect 71681 78026 71747 78029
rect 103605 78026 103671 78029
rect 70945 78024 103671 78026
rect 70945 77968 70950 78024
rect 71006 77968 71686 78024
rect 71742 77968 103610 78024
rect 103666 77968 103671 78024
rect 70945 77966 103671 77968
rect 70945 77963 71011 77966
rect 71681 77963 71747 77966
rect 103605 77963 103671 77966
rect 31201 77890 31267 77893
rect 8109 77888 16590 77890
rect 8109 77832 8114 77888
rect 8170 77832 16590 77888
rect 8109 77830 16590 77832
rect 26190 77888 31267 77890
rect 26190 77832 31206 77888
rect 31262 77832 31267 77888
rect 26190 77830 31267 77832
rect 8109 77827 8175 77830
rect 4210 77824 4526 77825
rect 4210 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4526 77824
rect 4210 77759 4526 77760
rect 7925 77754 7991 77757
rect 26190 77754 26250 77830
rect 31201 77827 31267 77830
rect 34930 77824 35246 77825
rect 34930 77760 34936 77824
rect 35000 77760 35016 77824
rect 35080 77760 35096 77824
rect 35160 77760 35176 77824
rect 35240 77760 35246 77824
rect 34930 77759 35246 77760
rect 65650 77824 65966 77825
rect 65650 77760 65656 77824
rect 65720 77760 65736 77824
rect 65800 77760 65816 77824
rect 65880 77760 65896 77824
rect 65960 77760 65966 77824
rect 65650 77759 65966 77760
rect 96370 77824 96686 77825
rect 96370 77760 96376 77824
rect 96440 77760 96456 77824
rect 96520 77760 96536 77824
rect 96600 77760 96616 77824
rect 96680 77760 96686 77824
rect 96370 77759 96686 77760
rect 105918 77824 106234 77825
rect 105918 77760 105924 77824
rect 105988 77760 106004 77824
rect 106068 77760 106084 77824
rect 106148 77760 106164 77824
rect 106228 77760 106234 77824
rect 105918 77759 106234 77760
rect 28165 77756 28231 77757
rect 28165 77754 28212 77756
rect 7925 77752 26250 77754
rect 7925 77696 7930 77752
rect 7986 77696 26250 77752
rect 7925 77694 26250 77696
rect 28120 77752 28212 77754
rect 28120 77696 28170 77752
rect 28120 77694 28212 77696
rect 7925 77691 7991 77694
rect 28165 77692 28212 77694
rect 28276 77692 28282 77756
rect 28165 77691 28231 77692
rect 0 77618 800 77648
rect 1301 77618 1367 77621
rect 0 77616 1367 77618
rect 0 77560 1306 77616
rect 1362 77560 1367 77616
rect 0 77558 1367 77560
rect 0 77528 800 77558
rect 1301 77555 1367 77558
rect 9489 77618 9555 77621
rect 42885 77618 42951 77621
rect 9489 77616 42951 77618
rect 9489 77560 9494 77616
rect 9550 77560 42890 77616
rect 42946 77560 42951 77616
rect 9489 77558 42951 77560
rect 9489 77555 9555 77558
rect 42885 77555 42951 77558
rect 68461 77618 68527 77621
rect 102317 77618 102383 77621
rect 68461 77616 102383 77618
rect 68461 77560 68466 77616
rect 68522 77560 102322 77616
rect 102378 77560 102383 77616
rect 68461 77558 102383 77560
rect 68461 77555 68527 77558
rect 102317 77555 102383 77558
rect 108481 77618 108547 77621
rect 109200 77618 110000 77648
rect 108481 77616 110000 77618
rect 108481 77560 108486 77616
rect 108542 77560 110000 77616
rect 108481 77558 110000 77560
rect 108481 77555 108547 77558
rect 109200 77528 110000 77558
rect 40033 77482 40099 77485
rect 43621 77482 43687 77485
rect 40033 77480 43687 77482
rect 40033 77424 40038 77480
rect 40094 77424 43626 77480
rect 43682 77424 43687 77480
rect 40033 77422 43687 77424
rect 40033 77419 40099 77422
rect 43621 77419 43687 77422
rect 65885 77482 65951 77485
rect 103973 77482 104039 77485
rect 65885 77480 104039 77482
rect 65885 77424 65890 77480
rect 65946 77424 103978 77480
rect 104034 77424 104039 77480
rect 65885 77422 104039 77424
rect 65885 77419 65951 77422
rect 103973 77419 104039 77422
rect 35985 77346 36051 77349
rect 37917 77346 37983 77349
rect 35985 77344 37983 77346
rect 35985 77288 35990 77344
rect 36046 77288 37922 77344
rect 37978 77288 37983 77344
rect 35985 77286 37983 77288
rect 35985 77283 36051 77286
rect 37917 77283 37983 77286
rect 39941 77346 40007 77349
rect 42425 77346 42491 77349
rect 39941 77344 42491 77346
rect 39941 77288 39946 77344
rect 40002 77288 42430 77344
rect 42486 77288 42491 77344
rect 39941 77286 42491 77288
rect 39941 77283 40007 77286
rect 42425 77283 42491 77286
rect 4870 77280 5186 77281
rect 4870 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5186 77280
rect 4870 77215 5186 77216
rect 35590 77280 35906 77281
rect 35590 77216 35596 77280
rect 35660 77216 35676 77280
rect 35740 77216 35756 77280
rect 35820 77216 35836 77280
rect 35900 77216 35906 77280
rect 35590 77215 35906 77216
rect 66310 77280 66626 77281
rect 66310 77216 66316 77280
rect 66380 77216 66396 77280
rect 66460 77216 66476 77280
rect 66540 77216 66556 77280
rect 66620 77216 66626 77280
rect 66310 77215 66626 77216
rect 97030 77280 97346 77281
rect 97030 77216 97036 77280
rect 97100 77216 97116 77280
rect 97180 77216 97196 77280
rect 97260 77216 97276 77280
rect 97340 77216 97346 77280
rect 97030 77215 97346 77216
rect 106654 77280 106970 77281
rect 106654 77216 106660 77280
rect 106724 77216 106740 77280
rect 106804 77216 106820 77280
rect 106884 77216 106900 77280
rect 106964 77216 106970 77280
rect 106654 77215 106970 77216
rect 90398 77148 90404 77212
rect 90468 77210 90474 77212
rect 90541 77210 90607 77213
rect 90468 77208 90607 77210
rect 90468 77152 90546 77208
rect 90602 77152 90607 77208
rect 90468 77150 90607 77152
rect 90468 77148 90474 77150
rect 90541 77147 90607 77150
rect 0 76938 800 76968
rect 1209 76938 1275 76941
rect 0 76936 1275 76938
rect 0 76880 1214 76936
rect 1270 76880 1275 76936
rect 0 76878 1275 76880
rect 0 76848 800 76878
rect 1209 76875 1275 76878
rect 108481 76938 108547 76941
rect 109200 76938 110000 76968
rect 108481 76936 110000 76938
rect 108481 76880 108486 76936
rect 108542 76880 110000 76936
rect 108481 76878 110000 76880
rect 108481 76875 108547 76878
rect 109200 76848 110000 76878
rect 4210 76736 4526 76737
rect 4210 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4526 76736
rect 4210 76671 4526 76672
rect 34930 76736 35246 76737
rect 34930 76672 34936 76736
rect 35000 76672 35016 76736
rect 35080 76672 35096 76736
rect 35160 76672 35176 76736
rect 35240 76672 35246 76736
rect 34930 76671 35246 76672
rect 65650 76736 65966 76737
rect 65650 76672 65656 76736
rect 65720 76672 65736 76736
rect 65800 76672 65816 76736
rect 65880 76672 65896 76736
rect 65960 76672 65966 76736
rect 65650 76671 65966 76672
rect 96370 76736 96686 76737
rect 96370 76672 96376 76736
rect 96440 76672 96456 76736
rect 96520 76672 96536 76736
rect 96600 76672 96616 76736
rect 96680 76672 96686 76736
rect 96370 76671 96686 76672
rect 841 76394 907 76397
rect 798 76392 907 76394
rect 798 76336 846 76392
rect 902 76336 907 76392
rect 798 76331 907 76336
rect 798 76288 858 76331
rect 0 76198 858 76288
rect 108481 76258 108547 76261
rect 109200 76258 110000 76288
rect 108481 76256 110000 76258
rect 108481 76200 108486 76256
rect 108542 76200 110000 76256
rect 108481 76198 110000 76200
rect 0 76168 800 76198
rect 108481 76195 108547 76198
rect 4870 76192 5186 76193
rect 4870 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5186 76192
rect 4870 76127 5186 76128
rect 35590 76192 35906 76193
rect 35590 76128 35596 76192
rect 35660 76128 35676 76192
rect 35740 76128 35756 76192
rect 35820 76128 35836 76192
rect 35900 76128 35906 76192
rect 35590 76127 35906 76128
rect 66310 76192 66626 76193
rect 66310 76128 66316 76192
rect 66380 76128 66396 76192
rect 66460 76128 66476 76192
rect 66540 76128 66556 76192
rect 66620 76128 66626 76192
rect 66310 76127 66626 76128
rect 97030 76192 97346 76193
rect 97030 76128 97036 76192
rect 97100 76128 97116 76192
rect 97180 76128 97196 76192
rect 97260 76128 97276 76192
rect 97340 76128 97346 76192
rect 109200 76168 110000 76198
rect 97030 76127 97346 76128
rect 4210 75648 4526 75649
rect 0 75578 800 75608
rect 4210 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4526 75648
rect 4210 75583 4526 75584
rect 34930 75648 35246 75649
rect 34930 75584 34936 75648
rect 35000 75584 35016 75648
rect 35080 75584 35096 75648
rect 35160 75584 35176 75648
rect 35240 75584 35246 75648
rect 34930 75583 35246 75584
rect 65650 75648 65966 75649
rect 65650 75584 65656 75648
rect 65720 75584 65736 75648
rect 65800 75584 65816 75648
rect 65880 75584 65896 75648
rect 65960 75584 65966 75648
rect 65650 75583 65966 75584
rect 96370 75648 96686 75649
rect 96370 75584 96376 75648
rect 96440 75584 96456 75648
rect 96520 75584 96536 75648
rect 96600 75584 96616 75648
rect 96680 75584 96686 75648
rect 96370 75583 96686 75584
rect 1393 75578 1459 75581
rect 0 75576 1459 75578
rect 0 75520 1398 75576
rect 1454 75520 1459 75576
rect 0 75518 1459 75520
rect 0 75488 800 75518
rect 1393 75515 1459 75518
rect 108481 75578 108547 75581
rect 109200 75578 110000 75608
rect 108481 75576 110000 75578
rect 108481 75520 108486 75576
rect 108542 75520 110000 75576
rect 108481 75518 110000 75520
rect 108481 75515 108547 75518
rect 109200 75488 110000 75518
rect 4870 75104 5186 75105
rect 4870 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5186 75104
rect 4870 75039 5186 75040
rect 35590 75104 35906 75105
rect 35590 75040 35596 75104
rect 35660 75040 35676 75104
rect 35740 75040 35756 75104
rect 35820 75040 35836 75104
rect 35900 75040 35906 75104
rect 35590 75039 35906 75040
rect 66310 75104 66626 75105
rect 66310 75040 66316 75104
rect 66380 75040 66396 75104
rect 66460 75040 66476 75104
rect 66540 75040 66556 75104
rect 66620 75040 66626 75104
rect 66310 75039 66626 75040
rect 97030 75104 97346 75105
rect 97030 75040 97036 75104
rect 97100 75040 97116 75104
rect 97180 75040 97196 75104
rect 97260 75040 97276 75104
rect 97340 75040 97346 75104
rect 97030 75039 97346 75040
rect 841 75034 907 75037
rect 798 75032 907 75034
rect 798 74976 846 75032
rect 902 74976 907 75032
rect 798 74971 907 74976
rect 798 74928 858 74971
rect 0 74838 858 74928
rect 108481 74898 108547 74901
rect 109200 74898 110000 74928
rect 108481 74896 110000 74898
rect 108481 74840 108486 74896
rect 108542 74840 110000 74896
rect 108481 74838 110000 74840
rect 0 74808 800 74838
rect 108481 74835 108547 74838
rect 109200 74808 110000 74838
rect 4210 74560 4526 74561
rect 4210 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4526 74560
rect 4210 74495 4526 74496
rect 34930 74560 35246 74561
rect 34930 74496 34936 74560
rect 35000 74496 35016 74560
rect 35080 74496 35096 74560
rect 35160 74496 35176 74560
rect 35240 74496 35246 74560
rect 34930 74495 35246 74496
rect 65650 74560 65966 74561
rect 65650 74496 65656 74560
rect 65720 74496 65736 74560
rect 65800 74496 65816 74560
rect 65880 74496 65896 74560
rect 65960 74496 65966 74560
rect 65650 74495 65966 74496
rect 96370 74560 96686 74561
rect 96370 74496 96376 74560
rect 96440 74496 96456 74560
rect 96520 74496 96536 74560
rect 96600 74496 96616 74560
rect 96680 74496 96686 74560
rect 96370 74495 96686 74496
rect 841 74354 907 74357
rect 798 74352 907 74354
rect 798 74296 846 74352
rect 902 74296 907 74352
rect 798 74291 907 74296
rect 798 74248 858 74291
rect 0 74158 858 74248
rect 108481 74218 108547 74221
rect 109200 74218 110000 74248
rect 108481 74216 110000 74218
rect 108481 74160 108486 74216
rect 108542 74160 110000 74216
rect 108481 74158 110000 74160
rect 0 74128 800 74158
rect 108481 74155 108547 74158
rect 109200 74128 110000 74158
rect 4870 74016 5186 74017
rect 4870 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5186 74016
rect 4870 73951 5186 73952
rect 35590 74016 35906 74017
rect 35590 73952 35596 74016
rect 35660 73952 35676 74016
rect 35740 73952 35756 74016
rect 35820 73952 35836 74016
rect 35900 73952 35906 74016
rect 35590 73951 35906 73952
rect 66310 74016 66626 74017
rect 66310 73952 66316 74016
rect 66380 73952 66396 74016
rect 66460 73952 66476 74016
rect 66540 73952 66556 74016
rect 66620 73952 66626 74016
rect 66310 73951 66626 73952
rect 97030 74016 97346 74017
rect 97030 73952 97036 74016
rect 97100 73952 97116 74016
rect 97180 73952 97196 74016
rect 97260 73952 97276 74016
rect 97340 73952 97346 74016
rect 97030 73951 97346 73952
rect 841 73674 907 73677
rect 798 73672 907 73674
rect 798 73616 846 73672
rect 902 73616 907 73672
rect 798 73611 907 73616
rect 798 73568 858 73611
rect 0 73478 858 73568
rect 108481 73538 108547 73541
rect 109200 73538 110000 73568
rect 108481 73536 110000 73538
rect 108481 73480 108486 73536
rect 108542 73480 110000 73536
rect 108481 73478 110000 73480
rect 0 73448 800 73478
rect 108481 73475 108547 73478
rect 4210 73472 4526 73473
rect 4210 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4526 73472
rect 4210 73407 4526 73408
rect 34930 73472 35246 73473
rect 34930 73408 34936 73472
rect 35000 73408 35016 73472
rect 35080 73408 35096 73472
rect 35160 73408 35176 73472
rect 35240 73408 35246 73472
rect 34930 73407 35246 73408
rect 65650 73472 65966 73473
rect 65650 73408 65656 73472
rect 65720 73408 65736 73472
rect 65800 73408 65816 73472
rect 65880 73408 65896 73472
rect 65960 73408 65966 73472
rect 65650 73407 65966 73408
rect 96370 73472 96686 73473
rect 96370 73408 96376 73472
rect 96440 73408 96456 73472
rect 96520 73408 96536 73472
rect 96600 73408 96616 73472
rect 96680 73408 96686 73472
rect 109200 73448 110000 73478
rect 96370 73407 96686 73408
rect 841 72994 907 72997
rect 798 72992 907 72994
rect 798 72936 846 72992
rect 902 72936 907 72992
rect 798 72931 907 72936
rect 798 72888 858 72931
rect 0 72798 858 72888
rect 4870 72928 5186 72929
rect 4870 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5186 72928
rect 4870 72863 5186 72864
rect 35590 72928 35906 72929
rect 35590 72864 35596 72928
rect 35660 72864 35676 72928
rect 35740 72864 35756 72928
rect 35820 72864 35836 72928
rect 35900 72864 35906 72928
rect 35590 72863 35906 72864
rect 66310 72928 66626 72929
rect 66310 72864 66316 72928
rect 66380 72864 66396 72928
rect 66460 72864 66476 72928
rect 66540 72864 66556 72928
rect 66620 72864 66626 72928
rect 66310 72863 66626 72864
rect 97030 72928 97346 72929
rect 97030 72864 97036 72928
rect 97100 72864 97116 72928
rect 97180 72864 97196 72928
rect 97260 72864 97276 72928
rect 97340 72864 97346 72928
rect 97030 72863 97346 72864
rect 108481 72858 108547 72861
rect 109200 72858 110000 72888
rect 108481 72856 110000 72858
rect 108481 72800 108486 72856
rect 108542 72800 110000 72856
rect 108481 72798 110000 72800
rect 0 72768 800 72798
rect 108481 72795 108547 72798
rect 109200 72768 110000 72798
rect 4210 72384 4526 72385
rect 4210 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4526 72384
rect 4210 72319 4526 72320
rect 34930 72384 35246 72385
rect 34930 72320 34936 72384
rect 35000 72320 35016 72384
rect 35080 72320 35096 72384
rect 35160 72320 35176 72384
rect 35240 72320 35246 72384
rect 34930 72319 35246 72320
rect 65650 72384 65966 72385
rect 65650 72320 65656 72384
rect 65720 72320 65736 72384
rect 65800 72320 65816 72384
rect 65880 72320 65896 72384
rect 65960 72320 65966 72384
rect 65650 72319 65966 72320
rect 96370 72384 96686 72385
rect 96370 72320 96376 72384
rect 96440 72320 96456 72384
rect 96520 72320 96536 72384
rect 96600 72320 96616 72384
rect 96680 72320 96686 72384
rect 96370 72319 96686 72320
rect 0 72178 800 72208
rect 1117 72178 1183 72181
rect 0 72176 1183 72178
rect 0 72120 1122 72176
rect 1178 72120 1183 72176
rect 0 72118 1183 72120
rect 0 72088 800 72118
rect 1117 72115 1183 72118
rect 4870 71840 5186 71841
rect 4870 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5186 71840
rect 4870 71775 5186 71776
rect 35590 71840 35906 71841
rect 35590 71776 35596 71840
rect 35660 71776 35676 71840
rect 35740 71776 35756 71840
rect 35820 71776 35836 71840
rect 35900 71776 35906 71840
rect 35590 71775 35906 71776
rect 66310 71840 66626 71841
rect 66310 71776 66316 71840
rect 66380 71776 66396 71840
rect 66460 71776 66476 71840
rect 66540 71776 66556 71840
rect 66620 71776 66626 71840
rect 66310 71775 66626 71776
rect 97030 71840 97346 71841
rect 97030 71776 97036 71840
rect 97100 71776 97116 71840
rect 97180 71776 97196 71840
rect 97260 71776 97276 71840
rect 97340 71776 97346 71840
rect 97030 71775 97346 71776
rect 4210 71296 4526 71297
rect 4210 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4526 71296
rect 4210 71231 4526 71232
rect 34930 71296 35246 71297
rect 34930 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35246 71296
rect 34930 71231 35246 71232
rect 65650 71296 65966 71297
rect 65650 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65966 71296
rect 65650 71231 65966 71232
rect 96370 71296 96686 71297
rect 96370 71232 96376 71296
rect 96440 71232 96456 71296
rect 96520 71232 96536 71296
rect 96600 71232 96616 71296
rect 96680 71232 96686 71296
rect 96370 71231 96686 71232
rect 4870 70752 5186 70753
rect 4870 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5186 70752
rect 4870 70687 5186 70688
rect 35590 70752 35906 70753
rect 35590 70688 35596 70752
rect 35660 70688 35676 70752
rect 35740 70688 35756 70752
rect 35820 70688 35836 70752
rect 35900 70688 35906 70752
rect 35590 70687 35906 70688
rect 66310 70752 66626 70753
rect 66310 70688 66316 70752
rect 66380 70688 66396 70752
rect 66460 70688 66476 70752
rect 66540 70688 66556 70752
rect 66620 70688 66626 70752
rect 66310 70687 66626 70688
rect 97030 70752 97346 70753
rect 97030 70688 97036 70752
rect 97100 70688 97116 70752
rect 97180 70688 97196 70752
rect 97260 70688 97276 70752
rect 97340 70688 97346 70752
rect 97030 70687 97346 70688
rect 4210 70208 4526 70209
rect 4210 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4526 70208
rect 4210 70143 4526 70144
rect 34930 70208 35246 70209
rect 34930 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35246 70208
rect 34930 70143 35246 70144
rect 65650 70208 65966 70209
rect 65650 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65966 70208
rect 65650 70143 65966 70144
rect 96370 70208 96686 70209
rect 96370 70144 96376 70208
rect 96440 70144 96456 70208
rect 96520 70144 96536 70208
rect 96600 70144 96616 70208
rect 96680 70144 96686 70208
rect 96370 70143 96686 70144
rect 4870 69664 5186 69665
rect 4870 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5186 69664
rect 4870 69599 5186 69600
rect 35590 69664 35906 69665
rect 35590 69600 35596 69664
rect 35660 69600 35676 69664
rect 35740 69600 35756 69664
rect 35820 69600 35836 69664
rect 35900 69600 35906 69664
rect 35590 69599 35906 69600
rect 66310 69664 66626 69665
rect 66310 69600 66316 69664
rect 66380 69600 66396 69664
rect 66460 69600 66476 69664
rect 66540 69600 66556 69664
rect 66620 69600 66626 69664
rect 66310 69599 66626 69600
rect 97030 69664 97346 69665
rect 97030 69600 97036 69664
rect 97100 69600 97116 69664
rect 97180 69600 97196 69664
rect 97260 69600 97276 69664
rect 97340 69600 97346 69664
rect 97030 69599 97346 69600
rect 4210 69120 4526 69121
rect 4210 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4526 69120
rect 4210 69055 4526 69056
rect 34930 69120 35246 69121
rect 34930 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35246 69120
rect 34930 69055 35246 69056
rect 65650 69120 65966 69121
rect 65650 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65966 69120
rect 65650 69055 65966 69056
rect 96370 69120 96686 69121
rect 96370 69056 96376 69120
rect 96440 69056 96456 69120
rect 96520 69056 96536 69120
rect 96600 69056 96616 69120
rect 96680 69056 96686 69120
rect 96370 69055 96686 69056
rect 87270 68988 87276 69052
rect 87340 69050 87346 69052
rect 87689 69050 87755 69053
rect 87340 69048 87755 69050
rect 87340 68992 87694 69048
rect 87750 68992 87755 69048
rect 87340 68990 87755 68992
rect 87340 68988 87346 68990
rect 87689 68987 87755 68990
rect 4870 68576 5186 68577
rect 4870 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5186 68576
rect 4870 68511 5186 68512
rect 35590 68576 35906 68577
rect 35590 68512 35596 68576
rect 35660 68512 35676 68576
rect 35740 68512 35756 68576
rect 35820 68512 35836 68576
rect 35900 68512 35906 68576
rect 35590 68511 35906 68512
rect 66310 68576 66626 68577
rect 66310 68512 66316 68576
rect 66380 68512 66396 68576
rect 66460 68512 66476 68576
rect 66540 68512 66556 68576
rect 66620 68512 66626 68576
rect 66310 68511 66626 68512
rect 97030 68576 97346 68577
rect 97030 68512 97036 68576
rect 97100 68512 97116 68576
rect 97180 68512 97196 68576
rect 97260 68512 97276 68576
rect 97340 68512 97346 68576
rect 97030 68511 97346 68512
rect 4210 68032 4526 68033
rect 4210 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4526 68032
rect 4210 67967 4526 67968
rect 34930 68032 35246 68033
rect 34930 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35246 68032
rect 34930 67967 35246 67968
rect 65650 68032 65966 68033
rect 65650 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65966 68032
rect 65650 67967 65966 67968
rect 96370 68032 96686 68033
rect 96370 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96686 68032
rect 96370 67967 96686 67968
rect 4870 67488 5186 67489
rect 4870 67424 4876 67488
rect 4940 67424 4956 67488
rect 5020 67424 5036 67488
rect 5100 67424 5116 67488
rect 5180 67424 5186 67488
rect 4870 67423 5186 67424
rect 35590 67488 35906 67489
rect 35590 67424 35596 67488
rect 35660 67424 35676 67488
rect 35740 67424 35756 67488
rect 35820 67424 35836 67488
rect 35900 67424 35906 67488
rect 35590 67423 35906 67424
rect 66310 67488 66626 67489
rect 66310 67424 66316 67488
rect 66380 67424 66396 67488
rect 66460 67424 66476 67488
rect 66540 67424 66556 67488
rect 66620 67424 66626 67488
rect 66310 67423 66626 67424
rect 97030 67488 97346 67489
rect 97030 67424 97036 67488
rect 97100 67424 97116 67488
rect 97180 67424 97196 67488
rect 97260 67424 97276 67488
rect 97340 67424 97346 67488
rect 97030 67423 97346 67424
rect 108481 67418 108547 67421
rect 109200 67418 110000 67448
rect 108481 67416 110000 67418
rect 108481 67360 108486 67416
rect 108542 67360 110000 67416
rect 108481 67358 110000 67360
rect 108481 67355 108547 67358
rect 109200 67328 110000 67358
rect 4210 66944 4526 66945
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 34930 66944 35246 66945
rect 34930 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35246 66944
rect 34930 66879 35246 66880
rect 65650 66944 65966 66945
rect 65650 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65966 66944
rect 65650 66879 65966 66880
rect 96370 66944 96686 66945
rect 96370 66880 96376 66944
rect 96440 66880 96456 66944
rect 96520 66880 96536 66944
rect 96600 66880 96616 66944
rect 96680 66880 96686 66944
rect 96370 66879 96686 66880
rect 4870 66400 5186 66401
rect 4870 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5186 66400
rect 4870 66335 5186 66336
rect 35590 66400 35906 66401
rect 35590 66336 35596 66400
rect 35660 66336 35676 66400
rect 35740 66336 35756 66400
rect 35820 66336 35836 66400
rect 35900 66336 35906 66400
rect 35590 66335 35906 66336
rect 66310 66400 66626 66401
rect 66310 66336 66316 66400
rect 66380 66336 66396 66400
rect 66460 66336 66476 66400
rect 66540 66336 66556 66400
rect 66620 66336 66626 66400
rect 66310 66335 66626 66336
rect 97030 66400 97346 66401
rect 97030 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97346 66400
rect 97030 66335 97346 66336
rect 106654 66400 106970 66401
rect 106654 66336 106660 66400
rect 106724 66336 106740 66400
rect 106804 66336 106820 66400
rect 106884 66336 106900 66400
rect 106964 66336 106970 66400
rect 106654 66335 106970 66336
rect 89437 66330 89503 66333
rect 91001 66330 91067 66333
rect 89437 66328 91067 66330
rect 89437 66272 89442 66328
rect 89498 66272 91006 66328
rect 91062 66272 91067 66328
rect 89437 66270 91067 66272
rect 89437 66267 89503 66270
rect 91001 66267 91067 66270
rect 36077 66196 36143 66197
rect 38469 66196 38535 66197
rect 41137 66196 41203 66197
rect 36077 66192 36124 66196
rect 36188 66194 36194 66196
rect 36077 66136 36082 66192
rect 36077 66132 36124 66136
rect 36188 66134 36234 66194
rect 38469 66192 38516 66196
rect 38580 66194 38586 66196
rect 41086 66194 41092 66196
rect 38469 66136 38474 66192
rect 36188 66132 36194 66134
rect 38469 66132 38516 66136
rect 38580 66134 38626 66194
rect 41046 66134 41092 66194
rect 41156 66192 41203 66196
rect 41198 66136 41203 66192
rect 38580 66132 38586 66134
rect 41086 66132 41092 66134
rect 41156 66132 41203 66136
rect 36077 66131 36143 66132
rect 38469 66131 38535 66132
rect 41137 66131 41203 66132
rect 43621 66196 43687 66197
rect 46105 66196 46171 66197
rect 43621 66192 43668 66196
rect 43732 66194 43738 66196
rect 46054 66194 46060 66196
rect 43621 66136 43626 66192
rect 43621 66132 43668 66136
rect 43732 66134 43778 66194
rect 46014 66134 46060 66194
rect 46124 66192 46171 66196
rect 46166 66136 46171 66192
rect 43732 66132 43738 66134
rect 46054 66132 46060 66134
rect 46124 66132 46171 66136
rect 43621 66131 43687 66132
rect 46105 66131 46171 66132
rect 48589 66196 48655 66197
rect 51073 66196 51139 66197
rect 48589 66192 48636 66196
rect 48700 66194 48706 66196
rect 51022 66194 51028 66196
rect 48589 66136 48594 66192
rect 48589 66132 48636 66136
rect 48700 66134 48746 66194
rect 50982 66134 51028 66194
rect 51092 66192 51139 66196
rect 51134 66136 51139 66192
rect 48700 66132 48706 66134
rect 51022 66132 51028 66134
rect 51092 66132 51139 66136
rect 48589 66131 48655 66132
rect 51073 66131 51139 66132
rect 53557 66196 53623 66197
rect 53557 66192 53604 66196
rect 53668 66194 53674 66196
rect 53557 66136 53562 66192
rect 53557 66132 53604 66136
rect 53668 66134 53714 66194
rect 53668 66132 53674 66134
rect 55990 66132 55996 66196
rect 56060 66194 56066 66196
rect 56133 66194 56199 66197
rect 58617 66196 58683 66197
rect 58566 66194 58572 66196
rect 56060 66192 56199 66194
rect 56060 66136 56138 66192
rect 56194 66136 56199 66192
rect 56060 66134 56199 66136
rect 58526 66134 58572 66194
rect 58636 66192 58683 66196
rect 58678 66136 58683 66192
rect 56060 66132 56066 66134
rect 53557 66131 53623 66132
rect 56133 66131 56199 66134
rect 58566 66132 58572 66134
rect 58636 66132 58683 66136
rect 58617 66131 58683 66132
rect 61101 66196 61167 66197
rect 63585 66196 63651 66197
rect 61101 66192 61148 66196
rect 61212 66194 61218 66196
rect 63534 66194 63540 66196
rect 61101 66136 61106 66192
rect 61101 66132 61148 66136
rect 61212 66134 61258 66194
rect 63494 66134 63540 66194
rect 63604 66192 63651 66196
rect 63646 66136 63651 66192
rect 61212 66132 61218 66134
rect 63534 66132 63540 66134
rect 63604 66132 63651 66136
rect 61101 66131 61167 66132
rect 63585 66131 63651 66132
rect 66069 66196 66135 66197
rect 68553 66196 68619 66197
rect 66069 66192 66116 66196
rect 66180 66194 66186 66196
rect 68502 66194 68508 66196
rect 66069 66136 66074 66192
rect 66069 66132 66116 66136
rect 66180 66134 66226 66194
rect 68462 66134 68508 66194
rect 68572 66192 68619 66196
rect 68614 66136 68619 66192
rect 66180 66132 66186 66134
rect 68502 66132 68508 66134
rect 68572 66132 68619 66136
rect 66069 66131 66135 66132
rect 68553 66131 68619 66132
rect 71037 66196 71103 66197
rect 73521 66196 73587 66197
rect 71037 66192 71084 66196
rect 71148 66194 71154 66196
rect 73470 66194 73476 66196
rect 71037 66136 71042 66192
rect 71037 66132 71084 66136
rect 71148 66134 71194 66194
rect 73430 66134 73476 66194
rect 73540 66192 73587 66196
rect 73582 66136 73587 66192
rect 71148 66132 71154 66134
rect 73470 66132 73476 66134
rect 73540 66132 73587 66136
rect 86166 66132 86172 66196
rect 86236 66194 86242 66196
rect 86309 66194 86375 66197
rect 86236 66192 86375 66194
rect 86236 66136 86314 66192
rect 86370 66136 86375 66192
rect 86236 66134 86375 66136
rect 86236 66132 86242 66134
rect 71037 66131 71103 66132
rect 73521 66131 73587 66132
rect 86309 66131 86375 66134
rect 89345 66194 89411 66197
rect 91921 66194 91987 66197
rect 89345 66192 91987 66194
rect 89345 66136 89350 66192
rect 89406 66136 91926 66192
rect 91982 66136 91987 66192
rect 89345 66134 91987 66136
rect 89345 66131 89411 66134
rect 91921 66131 91987 66134
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 34930 65856 35246 65857
rect 34930 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35246 65856
rect 34930 65791 35246 65792
rect 65650 65856 65966 65857
rect 65650 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65966 65856
rect 65650 65791 65966 65792
rect 96370 65856 96686 65857
rect 96370 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96686 65856
rect 96370 65791 96686 65792
rect 105918 65856 106234 65857
rect 105918 65792 105924 65856
rect 105988 65792 106004 65856
rect 106068 65792 106084 65856
rect 106148 65792 106164 65856
rect 106228 65792 106234 65856
rect 105918 65791 106234 65792
rect 4870 65312 5186 65313
rect 4870 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5186 65312
rect 4870 65247 5186 65248
rect 106654 65312 106970 65313
rect 106654 65248 106660 65312
rect 106724 65248 106740 65312
rect 106804 65248 106820 65312
rect 106884 65248 106900 65312
rect 106964 65248 106970 65312
rect 106654 65247 106970 65248
rect 4210 64768 4526 64769
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 105918 64768 106234 64769
rect 105918 64704 105924 64768
rect 105988 64704 106004 64768
rect 106068 64704 106084 64768
rect 106148 64704 106164 64768
rect 106228 64704 106234 64768
rect 105918 64703 106234 64704
rect 4870 64224 5186 64225
rect 4870 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5186 64224
rect 4870 64159 5186 64160
rect 106654 64224 106970 64225
rect 106654 64160 106660 64224
rect 106724 64160 106740 64224
rect 106804 64160 106820 64224
rect 106884 64160 106900 64224
rect 106964 64160 106970 64224
rect 106654 64159 106970 64160
rect 95877 64156 95943 64157
rect 95852 64092 95858 64156
rect 95922 64154 95943 64156
rect 95922 64152 96014 64154
rect 95938 64096 96014 64152
rect 95922 64094 96014 64096
rect 95922 64092 95943 64094
rect 95877 64091 95943 64092
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 105918 63680 106234 63681
rect 105918 63616 105924 63680
rect 105988 63616 106004 63680
rect 106068 63616 106084 63680
rect 106148 63616 106164 63680
rect 106228 63616 106234 63680
rect 105918 63615 106234 63616
rect 4870 63136 5186 63137
rect 4870 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5186 63136
rect 4870 63071 5186 63072
rect 106654 63136 106970 63137
rect 106654 63072 106660 63136
rect 106724 63072 106740 63136
rect 106804 63072 106820 63136
rect 106884 63072 106900 63136
rect 106964 63072 106970 63136
rect 106654 63071 106970 63072
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 4210 62527 4526 62528
rect 105918 62592 106234 62593
rect 105918 62528 105924 62592
rect 105988 62528 106004 62592
rect 106068 62528 106084 62592
rect 106148 62528 106164 62592
rect 106228 62528 106234 62592
rect 105918 62527 106234 62528
rect 4870 62048 5186 62049
rect 4870 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5186 62048
rect 4870 61983 5186 61984
rect 106654 62048 106970 62049
rect 106654 61984 106660 62048
rect 106724 61984 106740 62048
rect 106804 61984 106820 62048
rect 106884 61984 106900 62048
rect 106964 61984 106970 62048
rect 106654 61983 106970 61984
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 105918 61504 106234 61505
rect 105918 61440 105924 61504
rect 105988 61440 106004 61504
rect 106068 61440 106084 61504
rect 106148 61440 106164 61504
rect 106228 61440 106234 61504
rect 105918 61439 106234 61440
rect 4870 60960 5186 60961
rect 4870 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5186 60960
rect 4870 60895 5186 60896
rect 106654 60960 106970 60961
rect 106654 60896 106660 60960
rect 106724 60896 106740 60960
rect 106804 60896 106820 60960
rect 106884 60896 106900 60960
rect 106964 60896 106970 60960
rect 106654 60895 106970 60896
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 105918 60416 106234 60417
rect 105918 60352 105924 60416
rect 105988 60352 106004 60416
rect 106068 60352 106084 60416
rect 106148 60352 106164 60416
rect 106228 60352 106234 60416
rect 105918 60351 106234 60352
rect 4870 59872 5186 59873
rect 4870 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5186 59872
rect 4870 59807 5186 59808
rect 106654 59872 106970 59873
rect 106654 59808 106660 59872
rect 106724 59808 106740 59872
rect 106804 59808 106820 59872
rect 106884 59808 106900 59872
rect 106964 59808 106970 59872
rect 106654 59807 106970 59808
rect 104341 59802 104407 59805
rect 102550 59800 104407 59802
rect 102550 59768 104346 59800
rect 101948 59744 104346 59768
rect 104402 59744 104407 59800
rect 101948 59742 104407 59744
rect 101948 59708 102610 59742
rect 104341 59739 104407 59742
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 105918 59328 106234 59329
rect 105918 59264 105924 59328
rect 105988 59264 106004 59328
rect 106068 59264 106084 59328
rect 106148 59264 106164 59328
rect 106228 59264 106234 59328
rect 105918 59263 106234 59264
rect 4870 58784 5186 58785
rect 4870 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5186 58784
rect 4870 58719 5186 58720
rect 106654 58784 106970 58785
rect 106654 58720 106660 58784
rect 106724 58720 106740 58784
rect 106804 58720 106820 58784
rect 106884 58720 106900 58784
rect 106964 58720 106970 58784
rect 106654 58719 106970 58720
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 105918 58240 106234 58241
rect 105918 58176 105924 58240
rect 105988 58176 106004 58240
rect 106068 58176 106084 58240
rect 106148 58176 106164 58240
rect 106228 58176 106234 58240
rect 105918 58175 106234 58176
rect 4870 57696 5186 57697
rect 4870 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5186 57696
rect 4870 57631 5186 57632
rect 106654 57696 106970 57697
rect 106654 57632 106660 57696
rect 106724 57632 106740 57696
rect 106804 57632 106820 57696
rect 106884 57632 106900 57696
rect 106964 57632 106970 57696
rect 106654 57631 106970 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 105918 57152 106234 57153
rect 105918 57088 105924 57152
rect 105988 57088 106004 57152
rect 106068 57088 106084 57152
rect 106148 57088 106164 57152
rect 106228 57088 106234 57152
rect 105918 57087 106234 57088
rect 4870 56608 5186 56609
rect 4870 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5186 56608
rect 4870 56543 5186 56544
rect 106654 56608 106970 56609
rect 106654 56544 106660 56608
rect 106724 56544 106740 56608
rect 106804 56544 106820 56608
rect 106884 56544 106900 56608
rect 106964 56544 106970 56608
rect 106654 56543 106970 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 105918 56064 106234 56065
rect 105918 56000 105924 56064
rect 105988 56000 106004 56064
rect 106068 56000 106084 56064
rect 106148 56000 106164 56064
rect 106228 56000 106234 56064
rect 105918 55999 106234 56000
rect 4870 55520 5186 55521
rect 4870 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5186 55520
rect 4870 55455 5186 55456
rect 106654 55520 106970 55521
rect 106654 55456 106660 55520
rect 106724 55456 106740 55520
rect 106804 55456 106820 55520
rect 106884 55456 106900 55520
rect 106964 55456 106970 55520
rect 106654 55455 106970 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 105918 54976 106234 54977
rect 105918 54912 105924 54976
rect 105988 54912 106004 54976
rect 106068 54912 106084 54976
rect 106148 54912 106164 54976
rect 106228 54912 106234 54976
rect 105918 54911 106234 54912
rect 4870 54432 5186 54433
rect 4870 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5186 54432
rect 4870 54367 5186 54368
rect 106654 54432 106970 54433
rect 106654 54368 106660 54432
rect 106724 54368 106740 54432
rect 106804 54368 106820 54432
rect 106884 54368 106900 54432
rect 106964 54368 106970 54432
rect 106654 54367 106970 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 105918 53888 106234 53889
rect 105918 53824 105924 53888
rect 105988 53824 106004 53888
rect 106068 53824 106084 53888
rect 106148 53824 106164 53888
rect 106228 53824 106234 53888
rect 105918 53823 106234 53824
rect 4870 53344 5186 53345
rect 4870 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5186 53344
rect 4870 53279 5186 53280
rect 106654 53344 106970 53345
rect 106654 53280 106660 53344
rect 106724 53280 106740 53344
rect 106804 53280 106820 53344
rect 106884 53280 106900 53344
rect 106964 53280 106970 53344
rect 106654 53279 106970 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 105918 52800 106234 52801
rect 105918 52736 105924 52800
rect 105988 52736 106004 52800
rect 106068 52736 106084 52800
rect 106148 52736 106164 52800
rect 106228 52736 106234 52800
rect 105918 52735 106234 52736
rect 4870 52256 5186 52257
rect 4870 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5186 52256
rect 4870 52191 5186 52192
rect 106654 52256 106970 52257
rect 106654 52192 106660 52256
rect 106724 52192 106740 52256
rect 106804 52192 106820 52256
rect 106884 52192 106900 52256
rect 106964 52192 106970 52256
rect 106654 52191 106970 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 105918 51712 106234 51713
rect 105918 51648 105924 51712
rect 105988 51648 106004 51712
rect 106068 51648 106084 51712
rect 106148 51648 106164 51712
rect 106228 51648 106234 51712
rect 105918 51647 106234 51648
rect 4870 51168 5186 51169
rect 4870 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5186 51168
rect 4870 51103 5186 51104
rect 106654 51168 106970 51169
rect 106654 51104 106660 51168
rect 106724 51104 106740 51168
rect 106804 51104 106820 51168
rect 106884 51104 106900 51168
rect 106964 51104 106970 51168
rect 106654 51103 106970 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 105918 50624 106234 50625
rect 105918 50560 105924 50624
rect 105988 50560 106004 50624
rect 106068 50560 106084 50624
rect 106148 50560 106164 50624
rect 106228 50560 106234 50624
rect 105918 50559 106234 50560
rect 4870 50080 5186 50081
rect 4870 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5186 50080
rect 4870 50015 5186 50016
rect 106654 50080 106970 50081
rect 106654 50016 106660 50080
rect 106724 50016 106740 50080
rect 106804 50016 106820 50080
rect 106884 50016 106900 50080
rect 106964 50016 106970 50080
rect 106654 50015 106970 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 105918 49536 106234 49537
rect 105918 49472 105924 49536
rect 105988 49472 106004 49536
rect 106068 49472 106084 49536
rect 106148 49472 106164 49536
rect 106228 49472 106234 49536
rect 105918 49471 106234 49472
rect 4870 48992 5186 48993
rect 4870 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5186 48992
rect 4870 48927 5186 48928
rect 106654 48992 106970 48993
rect 106654 48928 106660 48992
rect 106724 48928 106740 48992
rect 106804 48928 106820 48992
rect 106884 48928 106900 48992
rect 106964 48928 106970 48992
rect 106654 48927 106970 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 105918 48448 106234 48449
rect 105918 48384 105924 48448
rect 105988 48384 106004 48448
rect 106068 48384 106084 48448
rect 106148 48384 106164 48448
rect 106228 48384 106234 48448
rect 105918 48383 106234 48384
rect 4870 47904 5186 47905
rect 4870 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5186 47904
rect 4870 47839 5186 47840
rect 106654 47904 106970 47905
rect 106654 47840 106660 47904
rect 106724 47840 106740 47904
rect 106804 47840 106820 47904
rect 106884 47840 106900 47904
rect 106964 47840 106970 47904
rect 106654 47839 106970 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 105918 47360 106234 47361
rect 105918 47296 105924 47360
rect 105988 47296 106004 47360
rect 106068 47296 106084 47360
rect 106148 47296 106164 47360
rect 106228 47296 106234 47360
rect 105918 47295 106234 47296
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 106654 46816 106970 46817
rect 106654 46752 106660 46816
rect 106724 46752 106740 46816
rect 106804 46752 106820 46816
rect 106884 46752 106900 46816
rect 106964 46752 106970 46816
rect 106654 46751 106970 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 105918 46272 106234 46273
rect 105918 46208 105924 46272
rect 105988 46208 106004 46272
rect 106068 46208 106084 46272
rect 106148 46208 106164 46272
rect 106228 46208 106234 46272
rect 105918 46207 106234 46208
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 106654 45728 106970 45729
rect 106654 45664 106660 45728
rect 106724 45664 106740 45728
rect 106804 45664 106820 45728
rect 106884 45664 106900 45728
rect 106964 45664 106970 45728
rect 106654 45663 106970 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 105918 45184 106234 45185
rect 105918 45120 105924 45184
rect 105988 45120 106004 45184
rect 106068 45120 106084 45184
rect 106148 45120 106164 45184
rect 106228 45120 106234 45184
rect 105918 45119 106234 45120
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 106654 44640 106970 44641
rect 106654 44576 106660 44640
rect 106724 44576 106740 44640
rect 106804 44576 106820 44640
rect 106884 44576 106900 44640
rect 106964 44576 106970 44640
rect 106654 44575 106970 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 105918 44096 106234 44097
rect 105918 44032 105924 44096
rect 105988 44032 106004 44096
rect 106068 44032 106084 44096
rect 106148 44032 106164 44096
rect 106228 44032 106234 44096
rect 105918 44031 106234 44032
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 106654 43552 106970 43553
rect 106654 43488 106660 43552
rect 106724 43488 106740 43552
rect 106804 43488 106820 43552
rect 106884 43488 106900 43552
rect 106964 43488 106970 43552
rect 106654 43487 106970 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 105918 43008 106234 43009
rect 105918 42944 105924 43008
rect 105988 42944 106004 43008
rect 106068 42944 106084 43008
rect 106148 42944 106164 43008
rect 106228 42944 106234 43008
rect 105918 42943 106234 42944
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 106654 42464 106970 42465
rect 106654 42400 106660 42464
rect 106724 42400 106740 42464
rect 106804 42400 106820 42464
rect 106884 42400 106900 42464
rect 106964 42400 106970 42464
rect 106654 42399 106970 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 105918 41920 106234 41921
rect 105918 41856 105924 41920
rect 105988 41856 106004 41920
rect 106068 41856 106084 41920
rect 106148 41856 106164 41920
rect 106228 41856 106234 41920
rect 105918 41855 106234 41856
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 106654 41376 106970 41377
rect 106654 41312 106660 41376
rect 106724 41312 106740 41376
rect 106804 41312 106820 41376
rect 106884 41312 106900 41376
rect 106964 41312 106970 41376
rect 106654 41311 106970 41312
rect 7557 41306 7623 41309
rect 7557 41304 9506 41306
rect 7557 41248 7562 41304
rect 7618 41254 9506 41304
rect 7618 41248 10028 41254
rect 7557 41246 10028 41248
rect 7557 41243 7623 41246
rect 9446 41194 10028 41246
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 105918 40832 106234 40833
rect 105918 40768 105924 40832
rect 105988 40768 106004 40832
rect 106068 40768 106084 40832
rect 106148 40768 106164 40832
rect 106228 40768 106234 40832
rect 105918 40767 106234 40768
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 106654 40288 106970 40289
rect 106654 40224 106660 40288
rect 106724 40224 106740 40288
rect 106804 40224 106820 40288
rect 106884 40224 106900 40288
rect 106964 40224 106970 40288
rect 106654 40223 106970 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 105918 39744 106234 39745
rect 105918 39680 105924 39744
rect 105988 39680 106004 39744
rect 106068 39680 106084 39744
rect 106148 39680 106164 39744
rect 106228 39680 106234 39744
rect 105918 39679 106234 39680
rect 7281 39538 7347 39541
rect 9446 39538 10028 39554
rect 7281 39536 10028 39538
rect 7281 39480 7286 39536
rect 7342 39494 10028 39536
rect 7342 39480 9506 39494
rect 7281 39478 9506 39480
rect 7281 39475 7347 39478
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 106654 39200 106970 39201
rect 106654 39136 106660 39200
rect 106724 39136 106740 39200
rect 106804 39136 106820 39200
rect 106884 39136 106900 39200
rect 106964 39136 106970 39200
rect 106654 39135 106970 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 105918 38656 106234 38657
rect 105918 38592 105924 38656
rect 105988 38592 106004 38656
rect 106068 38592 106084 38656
rect 106148 38592 106164 38656
rect 106228 38592 106234 38656
rect 105918 38591 106234 38592
rect 7557 38450 7623 38453
rect 7557 38448 9506 38450
rect 7557 38392 7562 38448
rect 7618 38426 9506 38448
rect 7618 38392 10028 38426
rect 7557 38390 10028 38392
rect 7557 38387 7623 38390
rect 9446 38366 10028 38390
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 106654 38112 106970 38113
rect 106654 38048 106660 38112
rect 106724 38048 106740 38112
rect 106804 38048 106820 38112
rect 106884 38048 106900 38112
rect 106964 38048 106970 38112
rect 106654 38047 106970 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 105918 37568 106234 37569
rect 105918 37504 105924 37568
rect 105988 37504 106004 37568
rect 106068 37504 106084 37568
rect 106148 37504 106164 37568
rect 106228 37504 106234 37568
rect 105918 37503 106234 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 106654 37024 106970 37025
rect 106654 36960 106660 37024
rect 106724 36960 106740 37024
rect 106804 36960 106820 37024
rect 106884 36960 106900 37024
rect 106964 36960 106970 37024
rect 106654 36959 106970 36960
rect 7557 36682 7623 36685
rect 9446 36682 10028 36726
rect 7557 36680 10028 36682
rect 7557 36624 7562 36680
rect 7618 36666 10028 36680
rect 7618 36624 9506 36666
rect 7557 36622 9506 36624
rect 7557 36619 7623 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 105918 36480 106234 36481
rect 105918 36416 105924 36480
rect 105988 36416 106004 36480
rect 106068 36416 106084 36480
rect 106148 36416 106164 36480
rect 106228 36416 106234 36480
rect 105918 36415 106234 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 106654 35936 106970 35937
rect 106654 35872 106660 35936
rect 106724 35872 106740 35936
rect 106804 35872 106820 35936
rect 106884 35872 106900 35936
rect 106964 35872 106970 35936
rect 106654 35871 106970 35872
rect 7465 35594 7531 35597
rect 9446 35594 10028 35643
rect 7465 35592 10028 35594
rect 7465 35536 7470 35592
rect 7526 35583 10028 35592
rect 7526 35536 9506 35583
rect 7465 35534 9506 35536
rect 7465 35531 7531 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 105918 35392 106234 35393
rect 105918 35328 105924 35392
rect 105988 35328 106004 35392
rect 106068 35328 106084 35392
rect 106148 35328 106164 35392
rect 106228 35328 106234 35392
rect 105918 35327 106234 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 106654 34848 106970 34849
rect 106654 34784 106660 34848
rect 106724 34784 106740 34848
rect 106804 34784 106820 34848
rect 106884 34784 106900 34848
rect 106964 34784 106970 34848
rect 106654 34783 106970 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 105918 34304 106234 34305
rect 105918 34240 105924 34304
rect 105988 34240 106004 34304
rect 106068 34240 106084 34304
rect 106148 34240 106164 34304
rect 106228 34240 106234 34304
rect 105918 34239 106234 34240
rect 7557 33962 7623 33965
rect 9446 33962 10028 33963
rect 7557 33960 10028 33962
rect 7557 33904 7562 33960
rect 7618 33904 10028 33960
rect 7557 33903 10028 33904
rect 7557 33902 9506 33903
rect 7557 33899 7623 33902
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 106654 33760 106970 33761
rect 106654 33696 106660 33760
rect 106724 33696 106740 33760
rect 106804 33696 106820 33760
rect 106884 33696 106900 33760
rect 106964 33696 106970 33760
rect 106654 33695 106970 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 105918 33216 106234 33217
rect 105918 33152 105924 33216
rect 105988 33152 106004 33216
rect 106068 33152 106084 33216
rect 106148 33152 106164 33216
rect 106228 33152 106234 33216
rect 105918 33151 106234 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 106654 32672 106970 32673
rect 106654 32608 106660 32672
rect 106724 32608 106740 32672
rect 106804 32608 106820 32672
rect 106884 32608 106900 32672
rect 106964 32608 106970 32672
rect 106654 32607 106970 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 105918 32128 106234 32129
rect 105918 32064 105924 32128
rect 105988 32064 106004 32128
rect 106068 32064 106084 32128
rect 106148 32064 106164 32128
rect 106228 32064 106234 32128
rect 105918 32063 106234 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 106654 31584 106970 31585
rect 106654 31520 106660 31584
rect 106724 31520 106740 31584
rect 106804 31520 106820 31584
rect 106884 31520 106900 31584
rect 106964 31520 106970 31584
rect 106654 31519 106970 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 105918 31040 106234 31041
rect 105918 30976 105924 31040
rect 105988 30976 106004 31040
rect 106068 30976 106084 31040
rect 106148 30976 106164 31040
rect 106228 30976 106234 31040
rect 105918 30975 106234 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 106654 30496 106970 30497
rect 106654 30432 106660 30496
rect 106724 30432 106740 30496
rect 106804 30432 106820 30496
rect 106884 30432 106900 30496
rect 106964 30432 106970 30496
rect 106654 30431 106970 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 105918 29952 106234 29953
rect 105918 29888 105924 29952
rect 105988 29888 106004 29952
rect 106068 29888 106084 29952
rect 106148 29888 106164 29952
rect 106228 29888 106234 29952
rect 105918 29887 106234 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 106654 29408 106970 29409
rect 106654 29344 106660 29408
rect 106724 29344 106740 29408
rect 106804 29344 106820 29408
rect 106884 29344 106900 29408
rect 106964 29344 106970 29408
rect 106654 29343 106970 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 105918 28864 106234 28865
rect 105918 28800 105924 28864
rect 105988 28800 106004 28864
rect 106068 28800 106084 28864
rect 106148 28800 106164 28864
rect 106228 28800 106234 28864
rect 105918 28799 106234 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 106654 28320 106970 28321
rect 106654 28256 106660 28320
rect 106724 28256 106740 28320
rect 106804 28256 106820 28320
rect 106884 28256 106900 28320
rect 106964 28256 106970 28320
rect 106654 28255 106970 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 105918 27776 106234 27777
rect 105918 27712 105924 27776
rect 105988 27712 106004 27776
rect 106068 27712 106084 27776
rect 106148 27712 106164 27776
rect 106228 27712 106234 27776
rect 105918 27711 106234 27712
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 106654 27232 106970 27233
rect 106654 27168 106660 27232
rect 106724 27168 106740 27232
rect 106804 27168 106820 27232
rect 106884 27168 106900 27232
rect 106964 27168 106970 27232
rect 106654 27167 106970 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 105918 26688 106234 26689
rect 105918 26624 105924 26688
rect 105988 26624 106004 26688
rect 106068 26624 106084 26688
rect 106148 26624 106164 26688
rect 106228 26624 106234 26688
rect 105918 26623 106234 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 106654 26144 106970 26145
rect 106654 26080 106660 26144
rect 106724 26080 106740 26144
rect 106804 26080 106820 26144
rect 106884 26080 106900 26144
rect 106964 26080 106970 26144
rect 106654 26079 106970 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 105918 25600 106234 25601
rect 105918 25536 105924 25600
rect 105988 25536 106004 25600
rect 106068 25536 106084 25600
rect 106148 25536 106164 25600
rect 106228 25536 106234 25600
rect 105918 25535 106234 25536
rect 102593 25122 102659 25125
rect 102550 25120 102659 25122
rect 102225 25090 102291 25093
rect 102550 25090 102598 25120
rect 101948 25088 102598 25090
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 101948 25032 102230 25088
rect 102286 25064 102598 25088
rect 102654 25064 102659 25120
rect 102286 25059 102659 25064
rect 102286 25032 102610 25059
rect 101948 25030 102610 25032
rect 106654 25056 106970 25057
rect 102225 25027 102291 25030
rect 4870 24991 5186 24992
rect 106654 24992 106660 25056
rect 106724 24992 106740 25056
rect 106804 24992 106820 25056
rect 106884 24992 106900 25056
rect 106964 24992 106970 25056
rect 106654 24991 106970 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 105918 24512 106234 24513
rect 105918 24448 105924 24512
rect 105988 24448 106004 24512
rect 106068 24448 106084 24512
rect 106148 24448 106164 24512
rect 106228 24448 106234 24512
rect 105918 24447 106234 24448
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 106654 23968 106970 23969
rect 106654 23904 106660 23968
rect 106724 23904 106740 23968
rect 106804 23904 106820 23968
rect 106884 23904 106900 23968
rect 106964 23904 106970 23968
rect 106654 23903 106970 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 105918 23424 106234 23425
rect 102041 23390 102107 23393
rect 4210 23359 4526 23360
rect 101948 23388 102107 23390
rect 101948 23332 102046 23388
rect 102102 23332 102107 23388
rect 105918 23360 105924 23424
rect 105988 23360 106004 23424
rect 106068 23360 106084 23424
rect 106148 23360 106164 23424
rect 106228 23360 106234 23424
rect 105918 23359 106234 23360
rect 101948 23330 102107 23332
rect 102041 23327 102107 23330
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 106654 22880 106970 22881
rect 106654 22816 106660 22880
rect 106724 22816 106740 22880
rect 106804 22816 106820 22880
rect 106884 22816 106900 22880
rect 106964 22816 106970 22880
rect 106654 22815 106970 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 105918 22336 106234 22337
rect 105918 22272 105924 22336
rect 105988 22272 106004 22336
rect 106068 22272 106084 22336
rect 106148 22272 106164 22336
rect 106228 22272 106234 22336
rect 105918 22271 106234 22272
rect 102317 22262 102383 22265
rect 101948 22260 102383 22262
rect 101948 22204 102322 22260
rect 102378 22204 102383 22260
rect 101948 22202 102383 22204
rect 102317 22199 102383 22202
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 106654 21792 106970 21793
rect 106654 21728 106660 21792
rect 106724 21728 106740 21792
rect 106804 21728 106820 21792
rect 106884 21728 106900 21792
rect 106964 21728 106970 21792
rect 106654 21727 106970 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 105918 21248 106234 21249
rect 105918 21184 105924 21248
rect 105988 21184 106004 21248
rect 106068 21184 106084 21248
rect 106148 21184 106164 21248
rect 106228 21184 106234 21248
rect 105918 21183 106234 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 106654 20704 106970 20705
rect 106654 20640 106660 20704
rect 106724 20640 106740 20704
rect 106804 20640 106820 20704
rect 106884 20640 106900 20704
rect 106964 20640 106970 20704
rect 106654 20639 106970 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 105918 20160 106234 20161
rect 105918 20096 105924 20160
rect 105988 20096 106004 20160
rect 106068 20096 106084 20160
rect 106148 20096 106164 20160
rect 106228 20096 106234 20160
rect 105918 20095 106234 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 106654 19616 106970 19617
rect 106654 19552 106660 19616
rect 106724 19552 106740 19616
rect 106804 19552 106820 19616
rect 106884 19552 106900 19616
rect 106964 19552 106970 19616
rect 106654 19551 106970 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 105918 19072 106234 19073
rect 105918 19008 105924 19072
rect 105988 19008 106004 19072
rect 106068 19008 106084 19072
rect 106148 19008 106164 19072
rect 106228 19008 106234 19072
rect 105918 19007 106234 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 106654 18528 106970 18529
rect 106654 18464 106660 18528
rect 106724 18464 106740 18528
rect 106804 18464 106820 18528
rect 106884 18464 106900 18528
rect 106964 18464 106970 18528
rect 106654 18463 106970 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 105918 17984 106234 17985
rect 105918 17920 105924 17984
rect 105988 17920 106004 17984
rect 106068 17920 106084 17984
rect 106148 17920 106164 17984
rect 106228 17920 106234 17984
rect 105918 17919 106234 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 106654 17440 106970 17441
rect 106654 17376 106660 17440
rect 106724 17376 106740 17440
rect 106804 17376 106820 17440
rect 106884 17376 106900 17440
rect 106964 17376 106970 17440
rect 106654 17375 106970 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 105918 16896 106234 16897
rect 105918 16832 105924 16896
rect 105988 16832 106004 16896
rect 106068 16832 106084 16896
rect 106148 16832 106164 16896
rect 106228 16832 106234 16896
rect 105918 16831 106234 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 106654 16352 106970 16353
rect 106654 16288 106660 16352
rect 106724 16288 106740 16352
rect 106804 16288 106820 16352
rect 106884 16288 106900 16352
rect 106964 16288 106970 16352
rect 106654 16287 106970 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 105918 15808 106234 15809
rect 105918 15744 105924 15808
rect 105988 15744 106004 15808
rect 106068 15744 106084 15808
rect 106148 15744 106164 15808
rect 106228 15744 106234 15808
rect 105918 15743 106234 15744
rect 7465 15466 7531 15469
rect 9446 15466 10028 15483
rect 7465 15464 10028 15466
rect 7465 15408 7470 15464
rect 7526 15423 10028 15464
rect 7526 15408 9506 15423
rect 7465 15406 9506 15408
rect 7465 15403 7531 15406
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 106654 15264 106970 15265
rect 106654 15200 106660 15264
rect 106724 15200 106740 15264
rect 106804 15200 106820 15264
rect 106884 15200 106900 15264
rect 106964 15200 106970 15264
rect 106654 15199 106970 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 105918 14720 106234 14721
rect 105918 14656 105924 14720
rect 105988 14656 106004 14720
rect 106068 14656 106084 14720
rect 106148 14656 106164 14720
rect 106228 14656 106234 14720
rect 105918 14655 106234 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 106654 14176 106970 14177
rect 106654 14112 106660 14176
rect 106724 14112 106740 14176
rect 106804 14112 106820 14176
rect 106884 14112 106900 14176
rect 106964 14112 106970 14176
rect 106654 14111 106970 14112
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 105918 13632 106234 13633
rect 105918 13568 105924 13632
rect 105988 13568 106004 13632
rect 106068 13568 106084 13632
rect 106148 13568 106164 13632
rect 106228 13568 106234 13632
rect 105918 13567 106234 13568
rect 4870 13088 5186 13089
rect 0 13018 800 13048
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 106654 13088 106970 13089
rect 106654 13024 106660 13088
rect 106724 13024 106740 13088
rect 106804 13024 106820 13088
rect 106884 13024 106900 13088
rect 106964 13024 106970 13088
rect 106654 13023 106970 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 105918 12544 106234 12545
rect 105918 12480 105924 12544
rect 105988 12480 106004 12544
rect 106068 12480 106084 12544
rect 106148 12480 106164 12544
rect 106228 12480 106234 12544
rect 105918 12479 106234 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 106654 12000 106970 12001
rect 106654 11936 106660 12000
rect 106724 11936 106740 12000
rect 106804 11936 106820 12000
rect 106884 11936 106900 12000
rect 106964 11936 106970 12000
rect 106654 11935 106970 11936
rect 0 11658 800 11688
rect 1209 11658 1275 11661
rect 0 11656 1275 11658
rect 0 11600 1214 11656
rect 1270 11600 1275 11656
rect 0 11598 1275 11600
rect 0 11568 800 11598
rect 1209 11595 1275 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 105918 11456 106234 11457
rect 105918 11392 105924 11456
rect 105988 11392 106004 11456
rect 106068 11392 106084 11456
rect 106148 11392 106164 11456
rect 106228 11392 106234 11456
rect 105918 11391 106234 11392
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 106654 10912 106970 10913
rect 106654 10848 106660 10912
rect 106724 10848 106740 10912
rect 106804 10848 106820 10912
rect 106884 10848 106900 10912
rect 106964 10848 106970 10912
rect 106654 10847 106970 10848
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 105918 10368 106234 10369
rect 105918 10304 105924 10368
rect 105988 10304 106004 10368
rect 106068 10304 106084 10368
rect 106148 10304 106164 10368
rect 106228 10304 106234 10368
rect 105918 10303 106234 10304
rect 1301 10298 1367 10301
rect 0 10296 1367 10298
rect 0 10240 1306 10296
rect 1362 10240 1367 10296
rect 0 10238 1367 10240
rect 0 10208 800 10238
rect 1301 10235 1367 10238
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 106654 9824 106970 9825
rect 106654 9760 106660 9824
rect 106724 9760 106740 9824
rect 106804 9760 106820 9824
rect 106884 9760 106900 9824
rect 106964 9760 106970 9824
rect 106654 9759 106970 9760
rect 23473 9756 23539 9757
rect 25773 9756 25839 9757
rect 28165 9756 28231 9757
rect 23432 9692 23438 9756
rect 23502 9754 23539 9756
rect 25768 9754 25774 9756
rect 23502 9752 23594 9754
rect 23534 9696 23594 9752
rect 23502 9694 23594 9696
rect 25686 9694 25774 9754
rect 23502 9692 23539 9694
rect 25768 9692 25774 9694
rect 25838 9692 25844 9756
rect 28114 9692 28120 9756
rect 28184 9754 28231 9756
rect 28184 9752 28276 9754
rect 28226 9696 28276 9752
rect 28184 9694 28276 9696
rect 28184 9692 28231 9694
rect 29272 9692 29278 9756
rect 29342 9754 29348 9756
rect 29545 9754 29611 9757
rect 30465 9756 30531 9757
rect 90541 9756 90607 9757
rect 29342 9752 29611 9754
rect 29342 9696 29550 9752
rect 29606 9696 29611 9752
rect 29342 9694 29611 9696
rect 29342 9692 29348 9694
rect 23473 9691 23539 9692
rect 25773 9691 25839 9692
rect 28165 9691 28231 9692
rect 29545 9691 29611 9694
rect 30440 9692 30446 9756
rect 30510 9754 30531 9756
rect 90521 9754 90527 9756
rect 30510 9752 30602 9754
rect 30526 9696 30602 9752
rect 30510 9694 30602 9696
rect 90450 9694 90527 9754
rect 90591 9752 90607 9756
rect 90602 9696 90607 9752
rect 30510 9692 30531 9694
rect 90521 9692 90527 9694
rect 90591 9692 90607 9696
rect 30465 9691 30531 9692
rect 90541 9691 90607 9692
rect 90909 9756 90975 9757
rect 90909 9752 90956 9756
rect 91020 9754 91026 9756
rect 90909 9696 90914 9752
rect 90909 9692 90956 9696
rect 91020 9694 91066 9754
rect 91020 9692 91026 9694
rect 90909 9691 90975 9692
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 16021 9620 16087 9621
rect 24669 9620 24735 9621
rect 90725 9620 90791 9621
rect 16021 9616 16058 9620
rect 16122 9618 16128 9620
rect 24618 9618 24624 9620
rect 16021 9560 16026 9616
rect 16021 9556 16058 9560
rect 16122 9558 16178 9618
rect 24578 9558 24624 9618
rect 24688 9616 24735 9620
rect 90674 9618 90680 9620
rect 24730 9560 24735 9616
rect 16122 9556 16128 9558
rect 24618 9556 24624 9558
rect 24688 9556 24735 9560
rect 90634 9558 90680 9618
rect 90744 9616 90791 9620
rect 90786 9560 90791 9616
rect 90674 9556 90680 9558
rect 90744 9556 90791 9560
rect 16021 9555 16087 9556
rect 24669 9555 24735 9556
rect 90725 9555 90791 9556
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 105918 9280 106234 9281
rect 105918 9216 105924 9280
rect 105988 9216 106004 9280
rect 106068 9216 106084 9280
rect 106148 9216 106164 9280
rect 106228 9216 106234 9280
rect 105918 9215 106234 9216
rect 0 8938 800 8968
rect 1301 8938 1367 8941
rect 0 8936 1367 8938
rect 0 8880 1306 8936
rect 1362 8880 1367 8936
rect 0 8878 1367 8880
rect 0 8848 800 8878
rect 1301 8875 1367 8878
rect 26693 8938 26759 8941
rect 26918 8938 26924 8940
rect 26693 8936 26924 8938
rect 26693 8880 26698 8936
rect 26754 8880 26924 8936
rect 26693 8878 26924 8880
rect 26693 8875 26759 8878
rect 26918 8876 26924 8878
rect 26988 8876 26994 8940
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 106654 8736 106970 8737
rect 106654 8672 106660 8736
rect 106724 8672 106740 8736
rect 106804 8672 106820 8736
rect 106884 8672 106900 8736
rect 106964 8672 106970 8736
rect 106654 8671 106970 8672
rect 0 8258 800 8288
rect 1945 8258 2011 8261
rect 31661 8260 31727 8261
rect 31661 8258 31708 8260
rect 0 8256 2011 8258
rect 0 8200 1950 8256
rect 2006 8200 2011 8256
rect 0 8198 2011 8200
rect 31616 8256 31708 8258
rect 31616 8200 31666 8256
rect 31616 8198 31708 8200
rect 0 8168 800 8198
rect 1945 8195 2011 8198
rect 31661 8196 31708 8198
rect 31772 8196 31778 8260
rect 32806 8196 32812 8260
rect 32876 8258 32882 8260
rect 32949 8258 33015 8261
rect 32876 8256 33015 8258
rect 32876 8200 32954 8256
rect 33010 8200 33015 8256
rect 32876 8198 33015 8200
rect 32876 8196 32882 8198
rect 31661 8195 31727 8196
rect 32949 8195 33015 8198
rect 33910 8196 33916 8260
rect 33980 8258 33986 8260
rect 34237 8258 34303 8261
rect 33980 8256 34303 8258
rect 33980 8200 34242 8256
rect 34298 8200 34303 8256
rect 33980 8198 34303 8200
rect 33980 8196 33986 8198
rect 34237 8195 34303 8198
rect 35198 8196 35204 8260
rect 35268 8258 35274 8260
rect 35433 8258 35499 8261
rect 36353 8260 36419 8261
rect 37457 8260 37523 8261
rect 38745 8260 38811 8261
rect 36302 8258 36308 8260
rect 35268 8256 35499 8258
rect 35268 8200 35438 8256
rect 35494 8200 35499 8256
rect 35268 8198 35499 8200
rect 36262 8198 36308 8258
rect 36372 8256 36419 8260
rect 37406 8258 37412 8260
rect 36414 8200 36419 8256
rect 35268 8196 35274 8198
rect 35433 8195 35499 8198
rect 36302 8196 36308 8198
rect 36372 8196 36419 8200
rect 37366 8198 37412 8258
rect 37476 8256 37523 8260
rect 38694 8258 38700 8260
rect 37518 8200 37523 8256
rect 37406 8196 37412 8198
rect 37476 8196 37523 8200
rect 38654 8198 38700 8258
rect 38764 8256 38811 8260
rect 38806 8200 38811 8256
rect 38694 8196 38700 8198
rect 38764 8196 38811 8200
rect 40902 8196 40908 8260
rect 40972 8258 40978 8260
rect 41321 8258 41387 8261
rect 40972 8256 41387 8258
rect 40972 8200 41326 8256
rect 41382 8200 41387 8256
rect 40972 8198 41387 8200
rect 40972 8196 40978 8198
rect 36353 8195 36419 8196
rect 37457 8195 37523 8196
rect 38745 8195 38811 8196
rect 41321 8195 41387 8198
rect 42149 8260 42215 8261
rect 42149 8256 42196 8260
rect 42260 8258 42266 8260
rect 42149 8200 42154 8256
rect 42149 8196 42196 8200
rect 42260 8198 42306 8258
rect 42260 8196 42266 8198
rect 43294 8196 43300 8260
rect 43364 8258 43370 8260
rect 43437 8258 43503 8261
rect 43364 8256 43503 8258
rect 43364 8200 43442 8256
rect 43498 8200 43503 8256
rect 43364 8198 43503 8200
rect 43364 8196 43370 8198
rect 42149 8195 42215 8196
rect 43437 8195 43503 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 105918 8192 106234 8193
rect 105918 8128 105924 8192
rect 105988 8128 106004 8192
rect 106068 8128 106084 8192
rect 106148 8128 106164 8192
rect 106228 8128 106234 8192
rect 105918 8127 106234 8128
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 66310 7648 66626 7649
rect 66310 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66626 7648
rect 66310 7583 66626 7584
rect 97030 7648 97346 7649
rect 97030 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97346 7648
rect 97030 7583 97346 7584
rect 106654 7648 106970 7649
rect 106654 7584 106660 7648
rect 106724 7584 106740 7648
rect 106804 7584 106820 7648
rect 106884 7584 106900 7648
rect 106964 7584 106970 7648
rect 106654 7583 106970 7584
rect 1301 7578 1367 7581
rect 0 7576 1367 7578
rect 0 7520 1306 7576
rect 1362 7520 1367 7576
rect 0 7518 1367 7520
rect 0 7488 800 7518
rect 1301 7515 1367 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 96370 7104 96686 7105
rect 96370 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96686 7104
rect 96370 7039 96686 7040
rect 105918 7104 106234 7105
rect 105918 7040 105924 7104
rect 105988 7040 106004 7104
rect 106068 7040 106084 7104
rect 106148 7040 106164 7104
rect 106228 7040 106234 7104
rect 105918 7039 106234 7040
rect 0 6898 800 6928
rect 1301 6898 1367 6901
rect 0 6896 1367 6898
rect 0 6840 1306 6896
rect 1362 6840 1367 6896
rect 0 6838 1367 6840
rect 0 6808 800 6838
rect 1301 6835 1367 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 66310 6560 66626 6561
rect 66310 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66626 6560
rect 66310 6495 66626 6496
rect 97030 6560 97346 6561
rect 97030 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97346 6560
rect 97030 6495 97346 6496
rect 0 6218 800 6248
rect 1209 6218 1275 6221
rect 0 6216 1275 6218
rect 0 6160 1214 6216
rect 1270 6160 1275 6216
rect 0 6158 1275 6160
rect 0 6128 800 6158
rect 1209 6155 1275 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 96370 6016 96686 6017
rect 96370 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96686 6016
rect 96370 5951 96686 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 66310 5472 66626 5473
rect 66310 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66626 5472
rect 66310 5407 66626 5408
rect 97030 5472 97346 5473
rect 97030 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97346 5472
rect 97030 5407 97346 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 96370 4928 96686 4929
rect 96370 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96686 4928
rect 96370 4863 96686 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 39798 4524 39804 4588
rect 39868 4586 39874 4588
rect 39941 4586 40007 4589
rect 39868 4584 40007 4586
rect 39868 4528 39946 4584
rect 40002 4528 40007 4584
rect 39868 4526 40007 4528
rect 39868 4524 39874 4526
rect 39941 4523 40007 4526
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 66310 4384 66626 4385
rect 66310 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66626 4384
rect 66310 4319 66626 4320
rect 97030 4384 97346 4385
rect 97030 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97346 4384
rect 97030 4319 97346 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 96370 3840 96686 3841
rect 96370 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96686 3840
rect 96370 3775 96686 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 66310 3296 66626 3297
rect 66310 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66626 3296
rect 66310 3231 66626 3232
rect 97030 3296 97346 3297
rect 97030 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97346 3296
rect 97030 3231 97346 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 96370 2752 96686 2753
rect 96370 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96686 2752
rect 96370 2687 96686 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 66310 2208 66626 2209
rect 66310 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66626 2208
rect 66310 2143 66626 2144
rect 97030 2208 97346 2209
rect 97030 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97346 2208
rect 97030 2143 97346 2144
<< via3 >>
rect 4216 147452 4280 147456
rect 4216 147396 4220 147452
rect 4220 147396 4276 147452
rect 4276 147396 4280 147452
rect 4216 147392 4280 147396
rect 4296 147452 4360 147456
rect 4296 147396 4300 147452
rect 4300 147396 4356 147452
rect 4356 147396 4360 147452
rect 4296 147392 4360 147396
rect 4376 147452 4440 147456
rect 4376 147396 4380 147452
rect 4380 147396 4436 147452
rect 4436 147396 4440 147452
rect 4376 147392 4440 147396
rect 4456 147452 4520 147456
rect 4456 147396 4460 147452
rect 4460 147396 4516 147452
rect 4516 147396 4520 147452
rect 4456 147392 4520 147396
rect 34936 147452 35000 147456
rect 34936 147396 34940 147452
rect 34940 147396 34996 147452
rect 34996 147396 35000 147452
rect 34936 147392 35000 147396
rect 35016 147452 35080 147456
rect 35016 147396 35020 147452
rect 35020 147396 35076 147452
rect 35076 147396 35080 147452
rect 35016 147392 35080 147396
rect 35096 147452 35160 147456
rect 35096 147396 35100 147452
rect 35100 147396 35156 147452
rect 35156 147396 35160 147452
rect 35096 147392 35160 147396
rect 35176 147452 35240 147456
rect 35176 147396 35180 147452
rect 35180 147396 35236 147452
rect 35236 147396 35240 147452
rect 35176 147392 35240 147396
rect 65656 147452 65720 147456
rect 65656 147396 65660 147452
rect 65660 147396 65716 147452
rect 65716 147396 65720 147452
rect 65656 147392 65720 147396
rect 65736 147452 65800 147456
rect 65736 147396 65740 147452
rect 65740 147396 65796 147452
rect 65796 147396 65800 147452
rect 65736 147392 65800 147396
rect 65816 147452 65880 147456
rect 65816 147396 65820 147452
rect 65820 147396 65876 147452
rect 65876 147396 65880 147452
rect 65816 147392 65880 147396
rect 65896 147452 65960 147456
rect 65896 147396 65900 147452
rect 65900 147396 65956 147452
rect 65956 147396 65960 147452
rect 65896 147392 65960 147396
rect 96376 147452 96440 147456
rect 96376 147396 96380 147452
rect 96380 147396 96436 147452
rect 96436 147396 96440 147452
rect 96376 147392 96440 147396
rect 96456 147452 96520 147456
rect 96456 147396 96460 147452
rect 96460 147396 96516 147452
rect 96516 147396 96520 147452
rect 96456 147392 96520 147396
rect 96536 147452 96600 147456
rect 96536 147396 96540 147452
rect 96540 147396 96596 147452
rect 96596 147396 96600 147452
rect 96536 147392 96600 147396
rect 96616 147452 96680 147456
rect 96616 147396 96620 147452
rect 96620 147396 96676 147452
rect 96676 147396 96680 147452
rect 96616 147392 96680 147396
rect 4876 146908 4940 146912
rect 4876 146852 4880 146908
rect 4880 146852 4936 146908
rect 4936 146852 4940 146908
rect 4876 146848 4940 146852
rect 4956 146908 5020 146912
rect 4956 146852 4960 146908
rect 4960 146852 5016 146908
rect 5016 146852 5020 146908
rect 4956 146848 5020 146852
rect 5036 146908 5100 146912
rect 5036 146852 5040 146908
rect 5040 146852 5096 146908
rect 5096 146852 5100 146908
rect 5036 146848 5100 146852
rect 5116 146908 5180 146912
rect 5116 146852 5120 146908
rect 5120 146852 5176 146908
rect 5176 146852 5180 146908
rect 5116 146848 5180 146852
rect 35596 146908 35660 146912
rect 35596 146852 35600 146908
rect 35600 146852 35656 146908
rect 35656 146852 35660 146908
rect 35596 146848 35660 146852
rect 35676 146908 35740 146912
rect 35676 146852 35680 146908
rect 35680 146852 35736 146908
rect 35736 146852 35740 146908
rect 35676 146848 35740 146852
rect 35756 146908 35820 146912
rect 35756 146852 35760 146908
rect 35760 146852 35816 146908
rect 35816 146852 35820 146908
rect 35756 146848 35820 146852
rect 35836 146908 35900 146912
rect 35836 146852 35840 146908
rect 35840 146852 35896 146908
rect 35896 146852 35900 146908
rect 35836 146848 35900 146852
rect 66316 146908 66380 146912
rect 66316 146852 66320 146908
rect 66320 146852 66376 146908
rect 66376 146852 66380 146908
rect 66316 146848 66380 146852
rect 66396 146908 66460 146912
rect 66396 146852 66400 146908
rect 66400 146852 66456 146908
rect 66456 146852 66460 146908
rect 66396 146848 66460 146852
rect 66476 146908 66540 146912
rect 66476 146852 66480 146908
rect 66480 146852 66536 146908
rect 66536 146852 66540 146908
rect 66476 146848 66540 146852
rect 66556 146908 66620 146912
rect 66556 146852 66560 146908
rect 66560 146852 66616 146908
rect 66616 146852 66620 146908
rect 66556 146848 66620 146852
rect 97036 146908 97100 146912
rect 97036 146852 97040 146908
rect 97040 146852 97096 146908
rect 97096 146852 97100 146908
rect 97036 146848 97100 146852
rect 97116 146908 97180 146912
rect 97116 146852 97120 146908
rect 97120 146852 97176 146908
rect 97176 146852 97180 146908
rect 97116 146848 97180 146852
rect 97196 146908 97260 146912
rect 97196 146852 97200 146908
rect 97200 146852 97256 146908
rect 97256 146852 97260 146908
rect 97196 146848 97260 146852
rect 97276 146908 97340 146912
rect 97276 146852 97280 146908
rect 97280 146852 97336 146908
rect 97336 146852 97340 146908
rect 97276 146848 97340 146852
rect 4216 146364 4280 146368
rect 4216 146308 4220 146364
rect 4220 146308 4276 146364
rect 4276 146308 4280 146364
rect 4216 146304 4280 146308
rect 4296 146364 4360 146368
rect 4296 146308 4300 146364
rect 4300 146308 4356 146364
rect 4356 146308 4360 146364
rect 4296 146304 4360 146308
rect 4376 146364 4440 146368
rect 4376 146308 4380 146364
rect 4380 146308 4436 146364
rect 4436 146308 4440 146364
rect 4376 146304 4440 146308
rect 4456 146364 4520 146368
rect 4456 146308 4460 146364
rect 4460 146308 4516 146364
rect 4516 146308 4520 146364
rect 4456 146304 4520 146308
rect 34936 146364 35000 146368
rect 34936 146308 34940 146364
rect 34940 146308 34996 146364
rect 34996 146308 35000 146364
rect 34936 146304 35000 146308
rect 35016 146364 35080 146368
rect 35016 146308 35020 146364
rect 35020 146308 35076 146364
rect 35076 146308 35080 146364
rect 35016 146304 35080 146308
rect 35096 146364 35160 146368
rect 35096 146308 35100 146364
rect 35100 146308 35156 146364
rect 35156 146308 35160 146364
rect 35096 146304 35160 146308
rect 35176 146364 35240 146368
rect 35176 146308 35180 146364
rect 35180 146308 35236 146364
rect 35236 146308 35240 146364
rect 35176 146304 35240 146308
rect 65656 146364 65720 146368
rect 65656 146308 65660 146364
rect 65660 146308 65716 146364
rect 65716 146308 65720 146364
rect 65656 146304 65720 146308
rect 65736 146364 65800 146368
rect 65736 146308 65740 146364
rect 65740 146308 65796 146364
rect 65796 146308 65800 146364
rect 65736 146304 65800 146308
rect 65816 146364 65880 146368
rect 65816 146308 65820 146364
rect 65820 146308 65876 146364
rect 65876 146308 65880 146364
rect 65816 146304 65880 146308
rect 65896 146364 65960 146368
rect 65896 146308 65900 146364
rect 65900 146308 65956 146364
rect 65956 146308 65960 146364
rect 65896 146304 65960 146308
rect 96376 146364 96440 146368
rect 96376 146308 96380 146364
rect 96380 146308 96436 146364
rect 96436 146308 96440 146364
rect 96376 146304 96440 146308
rect 96456 146364 96520 146368
rect 96456 146308 96460 146364
rect 96460 146308 96516 146364
rect 96516 146308 96520 146364
rect 96456 146304 96520 146308
rect 96536 146364 96600 146368
rect 96536 146308 96540 146364
rect 96540 146308 96596 146364
rect 96596 146308 96600 146364
rect 96536 146304 96600 146308
rect 96616 146364 96680 146368
rect 96616 146308 96620 146364
rect 96620 146308 96676 146364
rect 96676 146308 96680 146364
rect 96616 146304 96680 146308
rect 4876 145820 4940 145824
rect 4876 145764 4880 145820
rect 4880 145764 4936 145820
rect 4936 145764 4940 145820
rect 4876 145760 4940 145764
rect 4956 145820 5020 145824
rect 4956 145764 4960 145820
rect 4960 145764 5016 145820
rect 5016 145764 5020 145820
rect 4956 145760 5020 145764
rect 5036 145820 5100 145824
rect 5036 145764 5040 145820
rect 5040 145764 5096 145820
rect 5096 145764 5100 145820
rect 5036 145760 5100 145764
rect 5116 145820 5180 145824
rect 5116 145764 5120 145820
rect 5120 145764 5176 145820
rect 5176 145764 5180 145820
rect 5116 145760 5180 145764
rect 35596 145820 35660 145824
rect 35596 145764 35600 145820
rect 35600 145764 35656 145820
rect 35656 145764 35660 145820
rect 35596 145760 35660 145764
rect 35676 145820 35740 145824
rect 35676 145764 35680 145820
rect 35680 145764 35736 145820
rect 35736 145764 35740 145820
rect 35676 145760 35740 145764
rect 35756 145820 35820 145824
rect 35756 145764 35760 145820
rect 35760 145764 35816 145820
rect 35816 145764 35820 145820
rect 35756 145760 35820 145764
rect 35836 145820 35900 145824
rect 35836 145764 35840 145820
rect 35840 145764 35896 145820
rect 35896 145764 35900 145820
rect 35836 145760 35900 145764
rect 66316 145820 66380 145824
rect 66316 145764 66320 145820
rect 66320 145764 66376 145820
rect 66376 145764 66380 145820
rect 66316 145760 66380 145764
rect 66396 145820 66460 145824
rect 66396 145764 66400 145820
rect 66400 145764 66456 145820
rect 66456 145764 66460 145820
rect 66396 145760 66460 145764
rect 66476 145820 66540 145824
rect 66476 145764 66480 145820
rect 66480 145764 66536 145820
rect 66536 145764 66540 145820
rect 66476 145760 66540 145764
rect 66556 145820 66620 145824
rect 66556 145764 66560 145820
rect 66560 145764 66616 145820
rect 66616 145764 66620 145820
rect 66556 145760 66620 145764
rect 97036 145820 97100 145824
rect 97036 145764 97040 145820
rect 97040 145764 97096 145820
rect 97096 145764 97100 145820
rect 97036 145760 97100 145764
rect 97116 145820 97180 145824
rect 97116 145764 97120 145820
rect 97120 145764 97176 145820
rect 97176 145764 97180 145820
rect 97116 145760 97180 145764
rect 97196 145820 97260 145824
rect 97196 145764 97200 145820
rect 97200 145764 97256 145820
rect 97256 145764 97260 145820
rect 97196 145760 97260 145764
rect 97276 145820 97340 145824
rect 97276 145764 97280 145820
rect 97280 145764 97336 145820
rect 97336 145764 97340 145820
rect 97276 145760 97340 145764
rect 4216 145276 4280 145280
rect 4216 145220 4220 145276
rect 4220 145220 4276 145276
rect 4276 145220 4280 145276
rect 4216 145216 4280 145220
rect 4296 145276 4360 145280
rect 4296 145220 4300 145276
rect 4300 145220 4356 145276
rect 4356 145220 4360 145276
rect 4296 145216 4360 145220
rect 4376 145276 4440 145280
rect 4376 145220 4380 145276
rect 4380 145220 4436 145276
rect 4436 145220 4440 145276
rect 4376 145216 4440 145220
rect 4456 145276 4520 145280
rect 4456 145220 4460 145276
rect 4460 145220 4516 145276
rect 4516 145220 4520 145276
rect 4456 145216 4520 145220
rect 34936 145276 35000 145280
rect 34936 145220 34940 145276
rect 34940 145220 34996 145276
rect 34996 145220 35000 145276
rect 34936 145216 35000 145220
rect 35016 145276 35080 145280
rect 35016 145220 35020 145276
rect 35020 145220 35076 145276
rect 35076 145220 35080 145276
rect 35016 145216 35080 145220
rect 35096 145276 35160 145280
rect 35096 145220 35100 145276
rect 35100 145220 35156 145276
rect 35156 145220 35160 145276
rect 35096 145216 35160 145220
rect 35176 145276 35240 145280
rect 35176 145220 35180 145276
rect 35180 145220 35236 145276
rect 35236 145220 35240 145276
rect 35176 145216 35240 145220
rect 65656 145276 65720 145280
rect 65656 145220 65660 145276
rect 65660 145220 65716 145276
rect 65716 145220 65720 145276
rect 65656 145216 65720 145220
rect 65736 145276 65800 145280
rect 65736 145220 65740 145276
rect 65740 145220 65796 145276
rect 65796 145220 65800 145276
rect 65736 145216 65800 145220
rect 65816 145276 65880 145280
rect 65816 145220 65820 145276
rect 65820 145220 65876 145276
rect 65876 145220 65880 145276
rect 65816 145216 65880 145220
rect 65896 145276 65960 145280
rect 65896 145220 65900 145276
rect 65900 145220 65956 145276
rect 65956 145220 65960 145276
rect 65896 145216 65960 145220
rect 96376 145276 96440 145280
rect 96376 145220 96380 145276
rect 96380 145220 96436 145276
rect 96436 145220 96440 145276
rect 96376 145216 96440 145220
rect 96456 145276 96520 145280
rect 96456 145220 96460 145276
rect 96460 145220 96516 145276
rect 96516 145220 96520 145276
rect 96456 145216 96520 145220
rect 96536 145276 96600 145280
rect 96536 145220 96540 145276
rect 96540 145220 96596 145276
rect 96596 145220 96600 145276
rect 96536 145216 96600 145220
rect 96616 145276 96680 145280
rect 96616 145220 96620 145276
rect 96620 145220 96676 145276
rect 96676 145220 96680 145276
rect 96616 145216 96680 145220
rect 4876 144732 4940 144736
rect 4876 144676 4880 144732
rect 4880 144676 4936 144732
rect 4936 144676 4940 144732
rect 4876 144672 4940 144676
rect 4956 144732 5020 144736
rect 4956 144676 4960 144732
rect 4960 144676 5016 144732
rect 5016 144676 5020 144732
rect 4956 144672 5020 144676
rect 5036 144732 5100 144736
rect 5036 144676 5040 144732
rect 5040 144676 5096 144732
rect 5096 144676 5100 144732
rect 5036 144672 5100 144676
rect 5116 144732 5180 144736
rect 5116 144676 5120 144732
rect 5120 144676 5176 144732
rect 5176 144676 5180 144732
rect 5116 144672 5180 144676
rect 35596 144732 35660 144736
rect 35596 144676 35600 144732
rect 35600 144676 35656 144732
rect 35656 144676 35660 144732
rect 35596 144672 35660 144676
rect 35676 144732 35740 144736
rect 35676 144676 35680 144732
rect 35680 144676 35736 144732
rect 35736 144676 35740 144732
rect 35676 144672 35740 144676
rect 35756 144732 35820 144736
rect 35756 144676 35760 144732
rect 35760 144676 35816 144732
rect 35816 144676 35820 144732
rect 35756 144672 35820 144676
rect 35836 144732 35900 144736
rect 35836 144676 35840 144732
rect 35840 144676 35896 144732
rect 35896 144676 35900 144732
rect 35836 144672 35900 144676
rect 66316 144732 66380 144736
rect 66316 144676 66320 144732
rect 66320 144676 66376 144732
rect 66376 144676 66380 144732
rect 66316 144672 66380 144676
rect 66396 144732 66460 144736
rect 66396 144676 66400 144732
rect 66400 144676 66456 144732
rect 66456 144676 66460 144732
rect 66396 144672 66460 144676
rect 66476 144732 66540 144736
rect 66476 144676 66480 144732
rect 66480 144676 66536 144732
rect 66536 144676 66540 144732
rect 66476 144672 66540 144676
rect 66556 144732 66620 144736
rect 66556 144676 66560 144732
rect 66560 144676 66616 144732
rect 66616 144676 66620 144732
rect 66556 144672 66620 144676
rect 97036 144732 97100 144736
rect 97036 144676 97040 144732
rect 97040 144676 97096 144732
rect 97096 144676 97100 144732
rect 97036 144672 97100 144676
rect 97116 144732 97180 144736
rect 97116 144676 97120 144732
rect 97120 144676 97176 144732
rect 97176 144676 97180 144732
rect 97116 144672 97180 144676
rect 97196 144732 97260 144736
rect 97196 144676 97200 144732
rect 97200 144676 97256 144732
rect 97256 144676 97260 144732
rect 97196 144672 97260 144676
rect 97276 144732 97340 144736
rect 97276 144676 97280 144732
rect 97280 144676 97336 144732
rect 97336 144676 97340 144732
rect 97276 144672 97340 144676
rect 4216 144188 4280 144192
rect 4216 144132 4220 144188
rect 4220 144132 4276 144188
rect 4276 144132 4280 144188
rect 4216 144128 4280 144132
rect 4296 144188 4360 144192
rect 4296 144132 4300 144188
rect 4300 144132 4356 144188
rect 4356 144132 4360 144188
rect 4296 144128 4360 144132
rect 4376 144188 4440 144192
rect 4376 144132 4380 144188
rect 4380 144132 4436 144188
rect 4436 144132 4440 144188
rect 4376 144128 4440 144132
rect 4456 144188 4520 144192
rect 4456 144132 4460 144188
rect 4460 144132 4516 144188
rect 4516 144132 4520 144188
rect 4456 144128 4520 144132
rect 34936 144188 35000 144192
rect 34936 144132 34940 144188
rect 34940 144132 34996 144188
rect 34996 144132 35000 144188
rect 34936 144128 35000 144132
rect 35016 144188 35080 144192
rect 35016 144132 35020 144188
rect 35020 144132 35076 144188
rect 35076 144132 35080 144188
rect 35016 144128 35080 144132
rect 35096 144188 35160 144192
rect 35096 144132 35100 144188
rect 35100 144132 35156 144188
rect 35156 144132 35160 144188
rect 35096 144128 35160 144132
rect 35176 144188 35240 144192
rect 35176 144132 35180 144188
rect 35180 144132 35236 144188
rect 35236 144132 35240 144188
rect 35176 144128 35240 144132
rect 65656 144188 65720 144192
rect 65656 144132 65660 144188
rect 65660 144132 65716 144188
rect 65716 144132 65720 144188
rect 65656 144128 65720 144132
rect 65736 144188 65800 144192
rect 65736 144132 65740 144188
rect 65740 144132 65796 144188
rect 65796 144132 65800 144188
rect 65736 144128 65800 144132
rect 65816 144188 65880 144192
rect 65816 144132 65820 144188
rect 65820 144132 65876 144188
rect 65876 144132 65880 144188
rect 65816 144128 65880 144132
rect 65896 144188 65960 144192
rect 65896 144132 65900 144188
rect 65900 144132 65956 144188
rect 65956 144132 65960 144188
rect 65896 144128 65960 144132
rect 96376 144188 96440 144192
rect 96376 144132 96380 144188
rect 96380 144132 96436 144188
rect 96436 144132 96440 144188
rect 96376 144128 96440 144132
rect 96456 144188 96520 144192
rect 96456 144132 96460 144188
rect 96460 144132 96516 144188
rect 96516 144132 96520 144188
rect 96456 144128 96520 144132
rect 96536 144188 96600 144192
rect 96536 144132 96540 144188
rect 96540 144132 96596 144188
rect 96596 144132 96600 144188
rect 96536 144128 96600 144132
rect 96616 144188 96680 144192
rect 96616 144132 96620 144188
rect 96620 144132 96676 144188
rect 96676 144132 96680 144188
rect 96616 144128 96680 144132
rect 4876 143644 4940 143648
rect 4876 143588 4880 143644
rect 4880 143588 4936 143644
rect 4936 143588 4940 143644
rect 4876 143584 4940 143588
rect 4956 143644 5020 143648
rect 4956 143588 4960 143644
rect 4960 143588 5016 143644
rect 5016 143588 5020 143644
rect 4956 143584 5020 143588
rect 5036 143644 5100 143648
rect 5036 143588 5040 143644
rect 5040 143588 5096 143644
rect 5096 143588 5100 143644
rect 5036 143584 5100 143588
rect 5116 143644 5180 143648
rect 5116 143588 5120 143644
rect 5120 143588 5176 143644
rect 5176 143588 5180 143644
rect 5116 143584 5180 143588
rect 35596 143644 35660 143648
rect 35596 143588 35600 143644
rect 35600 143588 35656 143644
rect 35656 143588 35660 143644
rect 35596 143584 35660 143588
rect 35676 143644 35740 143648
rect 35676 143588 35680 143644
rect 35680 143588 35736 143644
rect 35736 143588 35740 143644
rect 35676 143584 35740 143588
rect 35756 143644 35820 143648
rect 35756 143588 35760 143644
rect 35760 143588 35816 143644
rect 35816 143588 35820 143644
rect 35756 143584 35820 143588
rect 35836 143644 35900 143648
rect 35836 143588 35840 143644
rect 35840 143588 35896 143644
rect 35896 143588 35900 143644
rect 35836 143584 35900 143588
rect 66316 143644 66380 143648
rect 66316 143588 66320 143644
rect 66320 143588 66376 143644
rect 66376 143588 66380 143644
rect 66316 143584 66380 143588
rect 66396 143644 66460 143648
rect 66396 143588 66400 143644
rect 66400 143588 66456 143644
rect 66456 143588 66460 143644
rect 66396 143584 66460 143588
rect 66476 143644 66540 143648
rect 66476 143588 66480 143644
rect 66480 143588 66536 143644
rect 66536 143588 66540 143644
rect 66476 143584 66540 143588
rect 66556 143644 66620 143648
rect 66556 143588 66560 143644
rect 66560 143588 66616 143644
rect 66616 143588 66620 143644
rect 66556 143584 66620 143588
rect 97036 143644 97100 143648
rect 97036 143588 97040 143644
rect 97040 143588 97096 143644
rect 97096 143588 97100 143644
rect 97036 143584 97100 143588
rect 97116 143644 97180 143648
rect 97116 143588 97120 143644
rect 97120 143588 97176 143644
rect 97176 143588 97180 143644
rect 97116 143584 97180 143588
rect 97196 143644 97260 143648
rect 97196 143588 97200 143644
rect 97200 143588 97256 143644
rect 97256 143588 97260 143644
rect 97196 143584 97260 143588
rect 97276 143644 97340 143648
rect 97276 143588 97280 143644
rect 97280 143588 97336 143644
rect 97336 143588 97340 143644
rect 97276 143584 97340 143588
rect 4216 143100 4280 143104
rect 4216 143044 4220 143100
rect 4220 143044 4276 143100
rect 4276 143044 4280 143100
rect 4216 143040 4280 143044
rect 4296 143100 4360 143104
rect 4296 143044 4300 143100
rect 4300 143044 4356 143100
rect 4356 143044 4360 143100
rect 4296 143040 4360 143044
rect 4376 143100 4440 143104
rect 4376 143044 4380 143100
rect 4380 143044 4436 143100
rect 4436 143044 4440 143100
rect 4376 143040 4440 143044
rect 4456 143100 4520 143104
rect 4456 143044 4460 143100
rect 4460 143044 4516 143100
rect 4516 143044 4520 143100
rect 4456 143040 4520 143044
rect 34936 143100 35000 143104
rect 34936 143044 34940 143100
rect 34940 143044 34996 143100
rect 34996 143044 35000 143100
rect 34936 143040 35000 143044
rect 35016 143100 35080 143104
rect 35016 143044 35020 143100
rect 35020 143044 35076 143100
rect 35076 143044 35080 143100
rect 35016 143040 35080 143044
rect 35096 143100 35160 143104
rect 35096 143044 35100 143100
rect 35100 143044 35156 143100
rect 35156 143044 35160 143100
rect 35096 143040 35160 143044
rect 35176 143100 35240 143104
rect 35176 143044 35180 143100
rect 35180 143044 35236 143100
rect 35236 143044 35240 143100
rect 35176 143040 35240 143044
rect 65656 143100 65720 143104
rect 65656 143044 65660 143100
rect 65660 143044 65716 143100
rect 65716 143044 65720 143100
rect 65656 143040 65720 143044
rect 65736 143100 65800 143104
rect 65736 143044 65740 143100
rect 65740 143044 65796 143100
rect 65796 143044 65800 143100
rect 65736 143040 65800 143044
rect 65816 143100 65880 143104
rect 65816 143044 65820 143100
rect 65820 143044 65876 143100
rect 65876 143044 65880 143100
rect 65816 143040 65880 143044
rect 65896 143100 65960 143104
rect 65896 143044 65900 143100
rect 65900 143044 65956 143100
rect 65956 143044 65960 143100
rect 65896 143040 65960 143044
rect 96376 143100 96440 143104
rect 96376 143044 96380 143100
rect 96380 143044 96436 143100
rect 96436 143044 96440 143100
rect 96376 143040 96440 143044
rect 96456 143100 96520 143104
rect 96456 143044 96460 143100
rect 96460 143044 96516 143100
rect 96516 143044 96520 143100
rect 96456 143040 96520 143044
rect 96536 143100 96600 143104
rect 96536 143044 96540 143100
rect 96540 143044 96596 143100
rect 96596 143044 96600 143100
rect 96536 143040 96600 143044
rect 96616 143100 96680 143104
rect 96616 143044 96620 143100
rect 96620 143044 96676 143100
rect 96676 143044 96680 143100
rect 96616 143040 96680 143044
rect 4876 142556 4940 142560
rect 4876 142500 4880 142556
rect 4880 142500 4936 142556
rect 4936 142500 4940 142556
rect 4876 142496 4940 142500
rect 4956 142556 5020 142560
rect 4956 142500 4960 142556
rect 4960 142500 5016 142556
rect 5016 142500 5020 142556
rect 4956 142496 5020 142500
rect 5036 142556 5100 142560
rect 5036 142500 5040 142556
rect 5040 142500 5096 142556
rect 5096 142500 5100 142556
rect 5036 142496 5100 142500
rect 5116 142556 5180 142560
rect 5116 142500 5120 142556
rect 5120 142500 5176 142556
rect 5176 142500 5180 142556
rect 5116 142496 5180 142500
rect 35596 142556 35660 142560
rect 35596 142500 35600 142556
rect 35600 142500 35656 142556
rect 35656 142500 35660 142556
rect 35596 142496 35660 142500
rect 35676 142556 35740 142560
rect 35676 142500 35680 142556
rect 35680 142500 35736 142556
rect 35736 142500 35740 142556
rect 35676 142496 35740 142500
rect 35756 142556 35820 142560
rect 35756 142500 35760 142556
rect 35760 142500 35816 142556
rect 35816 142500 35820 142556
rect 35756 142496 35820 142500
rect 35836 142556 35900 142560
rect 35836 142500 35840 142556
rect 35840 142500 35896 142556
rect 35896 142500 35900 142556
rect 35836 142496 35900 142500
rect 66316 142556 66380 142560
rect 66316 142500 66320 142556
rect 66320 142500 66376 142556
rect 66376 142500 66380 142556
rect 66316 142496 66380 142500
rect 66396 142556 66460 142560
rect 66396 142500 66400 142556
rect 66400 142500 66456 142556
rect 66456 142500 66460 142556
rect 66396 142496 66460 142500
rect 66476 142556 66540 142560
rect 66476 142500 66480 142556
rect 66480 142500 66536 142556
rect 66536 142500 66540 142556
rect 66476 142496 66540 142500
rect 66556 142556 66620 142560
rect 66556 142500 66560 142556
rect 66560 142500 66616 142556
rect 66616 142500 66620 142556
rect 66556 142496 66620 142500
rect 97036 142556 97100 142560
rect 97036 142500 97040 142556
rect 97040 142500 97096 142556
rect 97096 142500 97100 142556
rect 97036 142496 97100 142500
rect 97116 142556 97180 142560
rect 97116 142500 97120 142556
rect 97120 142500 97176 142556
rect 97176 142500 97180 142556
rect 97116 142496 97180 142500
rect 97196 142556 97260 142560
rect 97196 142500 97200 142556
rect 97200 142500 97256 142556
rect 97256 142500 97260 142556
rect 97196 142496 97260 142500
rect 97276 142556 97340 142560
rect 97276 142500 97280 142556
rect 97280 142500 97336 142556
rect 97336 142500 97340 142556
rect 97276 142496 97340 142500
rect 4216 142012 4280 142016
rect 4216 141956 4220 142012
rect 4220 141956 4276 142012
rect 4276 141956 4280 142012
rect 4216 141952 4280 141956
rect 4296 142012 4360 142016
rect 4296 141956 4300 142012
rect 4300 141956 4356 142012
rect 4356 141956 4360 142012
rect 4296 141952 4360 141956
rect 4376 142012 4440 142016
rect 4376 141956 4380 142012
rect 4380 141956 4436 142012
rect 4436 141956 4440 142012
rect 4376 141952 4440 141956
rect 4456 142012 4520 142016
rect 4456 141956 4460 142012
rect 4460 141956 4516 142012
rect 4516 141956 4520 142012
rect 4456 141952 4520 141956
rect 34936 142012 35000 142016
rect 34936 141956 34940 142012
rect 34940 141956 34996 142012
rect 34996 141956 35000 142012
rect 34936 141952 35000 141956
rect 35016 142012 35080 142016
rect 35016 141956 35020 142012
rect 35020 141956 35076 142012
rect 35076 141956 35080 142012
rect 35016 141952 35080 141956
rect 35096 142012 35160 142016
rect 35096 141956 35100 142012
rect 35100 141956 35156 142012
rect 35156 141956 35160 142012
rect 35096 141952 35160 141956
rect 35176 142012 35240 142016
rect 35176 141956 35180 142012
rect 35180 141956 35236 142012
rect 35236 141956 35240 142012
rect 35176 141952 35240 141956
rect 65656 142012 65720 142016
rect 65656 141956 65660 142012
rect 65660 141956 65716 142012
rect 65716 141956 65720 142012
rect 65656 141952 65720 141956
rect 65736 142012 65800 142016
rect 65736 141956 65740 142012
rect 65740 141956 65796 142012
rect 65796 141956 65800 142012
rect 65736 141952 65800 141956
rect 65816 142012 65880 142016
rect 65816 141956 65820 142012
rect 65820 141956 65876 142012
rect 65876 141956 65880 142012
rect 65816 141952 65880 141956
rect 65896 142012 65960 142016
rect 65896 141956 65900 142012
rect 65900 141956 65956 142012
rect 65956 141956 65960 142012
rect 65896 141952 65960 141956
rect 96376 142012 96440 142016
rect 96376 141956 96380 142012
rect 96380 141956 96436 142012
rect 96436 141956 96440 142012
rect 96376 141952 96440 141956
rect 96456 142012 96520 142016
rect 96456 141956 96460 142012
rect 96460 141956 96516 142012
rect 96516 141956 96520 142012
rect 96456 141952 96520 141956
rect 96536 142012 96600 142016
rect 96536 141956 96540 142012
rect 96540 141956 96596 142012
rect 96596 141956 96600 142012
rect 96536 141952 96600 141956
rect 96616 142012 96680 142016
rect 96616 141956 96620 142012
rect 96620 141956 96676 142012
rect 96676 141956 96680 142012
rect 96616 141952 96680 141956
rect 4876 141468 4940 141472
rect 4876 141412 4880 141468
rect 4880 141412 4936 141468
rect 4936 141412 4940 141468
rect 4876 141408 4940 141412
rect 4956 141468 5020 141472
rect 4956 141412 4960 141468
rect 4960 141412 5016 141468
rect 5016 141412 5020 141468
rect 4956 141408 5020 141412
rect 5036 141468 5100 141472
rect 5036 141412 5040 141468
rect 5040 141412 5096 141468
rect 5096 141412 5100 141468
rect 5036 141408 5100 141412
rect 5116 141468 5180 141472
rect 5116 141412 5120 141468
rect 5120 141412 5176 141468
rect 5176 141412 5180 141468
rect 5116 141408 5180 141412
rect 35596 141468 35660 141472
rect 35596 141412 35600 141468
rect 35600 141412 35656 141468
rect 35656 141412 35660 141468
rect 35596 141408 35660 141412
rect 35676 141468 35740 141472
rect 35676 141412 35680 141468
rect 35680 141412 35736 141468
rect 35736 141412 35740 141468
rect 35676 141408 35740 141412
rect 35756 141468 35820 141472
rect 35756 141412 35760 141468
rect 35760 141412 35816 141468
rect 35816 141412 35820 141468
rect 35756 141408 35820 141412
rect 35836 141468 35900 141472
rect 35836 141412 35840 141468
rect 35840 141412 35896 141468
rect 35896 141412 35900 141468
rect 35836 141408 35900 141412
rect 66316 141468 66380 141472
rect 66316 141412 66320 141468
rect 66320 141412 66376 141468
rect 66376 141412 66380 141468
rect 66316 141408 66380 141412
rect 66396 141468 66460 141472
rect 66396 141412 66400 141468
rect 66400 141412 66456 141468
rect 66456 141412 66460 141468
rect 66396 141408 66460 141412
rect 66476 141468 66540 141472
rect 66476 141412 66480 141468
rect 66480 141412 66536 141468
rect 66536 141412 66540 141468
rect 66476 141408 66540 141412
rect 66556 141468 66620 141472
rect 66556 141412 66560 141468
rect 66560 141412 66616 141468
rect 66616 141412 66620 141468
rect 66556 141408 66620 141412
rect 97036 141468 97100 141472
rect 97036 141412 97040 141468
rect 97040 141412 97096 141468
rect 97096 141412 97100 141468
rect 97036 141408 97100 141412
rect 97116 141468 97180 141472
rect 97116 141412 97120 141468
rect 97120 141412 97176 141468
rect 97176 141412 97180 141468
rect 97116 141408 97180 141412
rect 97196 141468 97260 141472
rect 97196 141412 97200 141468
rect 97200 141412 97256 141468
rect 97256 141412 97260 141468
rect 97196 141408 97260 141412
rect 97276 141468 97340 141472
rect 97276 141412 97280 141468
rect 97280 141412 97336 141468
rect 97336 141412 97340 141468
rect 97276 141408 97340 141412
rect 4216 140924 4280 140928
rect 4216 140868 4220 140924
rect 4220 140868 4276 140924
rect 4276 140868 4280 140924
rect 4216 140864 4280 140868
rect 4296 140924 4360 140928
rect 4296 140868 4300 140924
rect 4300 140868 4356 140924
rect 4356 140868 4360 140924
rect 4296 140864 4360 140868
rect 4376 140924 4440 140928
rect 4376 140868 4380 140924
rect 4380 140868 4436 140924
rect 4436 140868 4440 140924
rect 4376 140864 4440 140868
rect 4456 140924 4520 140928
rect 4456 140868 4460 140924
rect 4460 140868 4516 140924
rect 4516 140868 4520 140924
rect 4456 140864 4520 140868
rect 34936 140924 35000 140928
rect 34936 140868 34940 140924
rect 34940 140868 34996 140924
rect 34996 140868 35000 140924
rect 34936 140864 35000 140868
rect 35016 140924 35080 140928
rect 35016 140868 35020 140924
rect 35020 140868 35076 140924
rect 35076 140868 35080 140924
rect 35016 140864 35080 140868
rect 35096 140924 35160 140928
rect 35096 140868 35100 140924
rect 35100 140868 35156 140924
rect 35156 140868 35160 140924
rect 35096 140864 35160 140868
rect 35176 140924 35240 140928
rect 35176 140868 35180 140924
rect 35180 140868 35236 140924
rect 35236 140868 35240 140924
rect 35176 140864 35240 140868
rect 65656 140924 65720 140928
rect 65656 140868 65660 140924
rect 65660 140868 65716 140924
rect 65716 140868 65720 140924
rect 65656 140864 65720 140868
rect 65736 140924 65800 140928
rect 65736 140868 65740 140924
rect 65740 140868 65796 140924
rect 65796 140868 65800 140924
rect 65736 140864 65800 140868
rect 65816 140924 65880 140928
rect 65816 140868 65820 140924
rect 65820 140868 65876 140924
rect 65876 140868 65880 140924
rect 65816 140864 65880 140868
rect 65896 140924 65960 140928
rect 65896 140868 65900 140924
rect 65900 140868 65956 140924
rect 65956 140868 65960 140924
rect 65896 140864 65960 140868
rect 96376 140924 96440 140928
rect 96376 140868 96380 140924
rect 96380 140868 96436 140924
rect 96436 140868 96440 140924
rect 96376 140864 96440 140868
rect 96456 140924 96520 140928
rect 96456 140868 96460 140924
rect 96460 140868 96516 140924
rect 96516 140868 96520 140924
rect 96456 140864 96520 140868
rect 96536 140924 96600 140928
rect 96536 140868 96540 140924
rect 96540 140868 96596 140924
rect 96596 140868 96600 140924
rect 96536 140864 96600 140868
rect 96616 140924 96680 140928
rect 96616 140868 96620 140924
rect 96620 140868 96676 140924
rect 96676 140868 96680 140924
rect 96616 140864 96680 140868
rect 4876 140380 4940 140384
rect 4876 140324 4880 140380
rect 4880 140324 4936 140380
rect 4936 140324 4940 140380
rect 4876 140320 4940 140324
rect 4956 140380 5020 140384
rect 4956 140324 4960 140380
rect 4960 140324 5016 140380
rect 5016 140324 5020 140380
rect 4956 140320 5020 140324
rect 5036 140380 5100 140384
rect 5036 140324 5040 140380
rect 5040 140324 5096 140380
rect 5096 140324 5100 140380
rect 5036 140320 5100 140324
rect 5116 140380 5180 140384
rect 5116 140324 5120 140380
rect 5120 140324 5176 140380
rect 5176 140324 5180 140380
rect 5116 140320 5180 140324
rect 35596 140380 35660 140384
rect 35596 140324 35600 140380
rect 35600 140324 35656 140380
rect 35656 140324 35660 140380
rect 35596 140320 35660 140324
rect 35676 140380 35740 140384
rect 35676 140324 35680 140380
rect 35680 140324 35736 140380
rect 35736 140324 35740 140380
rect 35676 140320 35740 140324
rect 35756 140380 35820 140384
rect 35756 140324 35760 140380
rect 35760 140324 35816 140380
rect 35816 140324 35820 140380
rect 35756 140320 35820 140324
rect 35836 140380 35900 140384
rect 35836 140324 35840 140380
rect 35840 140324 35896 140380
rect 35896 140324 35900 140380
rect 35836 140320 35900 140324
rect 66316 140380 66380 140384
rect 66316 140324 66320 140380
rect 66320 140324 66376 140380
rect 66376 140324 66380 140380
rect 66316 140320 66380 140324
rect 66396 140380 66460 140384
rect 66396 140324 66400 140380
rect 66400 140324 66456 140380
rect 66456 140324 66460 140380
rect 66396 140320 66460 140324
rect 66476 140380 66540 140384
rect 66476 140324 66480 140380
rect 66480 140324 66536 140380
rect 66536 140324 66540 140380
rect 66476 140320 66540 140324
rect 66556 140380 66620 140384
rect 66556 140324 66560 140380
rect 66560 140324 66616 140380
rect 66616 140324 66620 140380
rect 66556 140320 66620 140324
rect 97036 140380 97100 140384
rect 97036 140324 97040 140380
rect 97040 140324 97096 140380
rect 97096 140324 97100 140380
rect 97036 140320 97100 140324
rect 97116 140380 97180 140384
rect 97116 140324 97120 140380
rect 97120 140324 97176 140380
rect 97176 140324 97180 140380
rect 97116 140320 97180 140324
rect 97196 140380 97260 140384
rect 97196 140324 97200 140380
rect 97200 140324 97256 140380
rect 97256 140324 97260 140380
rect 97196 140320 97260 140324
rect 97276 140380 97340 140384
rect 97276 140324 97280 140380
rect 97280 140324 97336 140380
rect 97336 140324 97340 140380
rect 97276 140320 97340 140324
rect 4216 139836 4280 139840
rect 4216 139780 4220 139836
rect 4220 139780 4276 139836
rect 4276 139780 4280 139836
rect 4216 139776 4280 139780
rect 4296 139836 4360 139840
rect 4296 139780 4300 139836
rect 4300 139780 4356 139836
rect 4356 139780 4360 139836
rect 4296 139776 4360 139780
rect 4376 139836 4440 139840
rect 4376 139780 4380 139836
rect 4380 139780 4436 139836
rect 4436 139780 4440 139836
rect 4376 139776 4440 139780
rect 4456 139836 4520 139840
rect 4456 139780 4460 139836
rect 4460 139780 4516 139836
rect 4516 139780 4520 139836
rect 4456 139776 4520 139780
rect 34936 139836 35000 139840
rect 34936 139780 34940 139836
rect 34940 139780 34996 139836
rect 34996 139780 35000 139836
rect 34936 139776 35000 139780
rect 35016 139836 35080 139840
rect 35016 139780 35020 139836
rect 35020 139780 35076 139836
rect 35076 139780 35080 139836
rect 35016 139776 35080 139780
rect 35096 139836 35160 139840
rect 35096 139780 35100 139836
rect 35100 139780 35156 139836
rect 35156 139780 35160 139836
rect 35096 139776 35160 139780
rect 35176 139836 35240 139840
rect 35176 139780 35180 139836
rect 35180 139780 35236 139836
rect 35236 139780 35240 139836
rect 35176 139776 35240 139780
rect 65656 139836 65720 139840
rect 65656 139780 65660 139836
rect 65660 139780 65716 139836
rect 65716 139780 65720 139836
rect 65656 139776 65720 139780
rect 65736 139836 65800 139840
rect 65736 139780 65740 139836
rect 65740 139780 65796 139836
rect 65796 139780 65800 139836
rect 65736 139776 65800 139780
rect 65816 139836 65880 139840
rect 65816 139780 65820 139836
rect 65820 139780 65876 139836
rect 65876 139780 65880 139836
rect 65816 139776 65880 139780
rect 65896 139836 65960 139840
rect 65896 139780 65900 139836
rect 65900 139780 65956 139836
rect 65956 139780 65960 139836
rect 65896 139776 65960 139780
rect 96376 139836 96440 139840
rect 96376 139780 96380 139836
rect 96380 139780 96436 139836
rect 96436 139780 96440 139836
rect 96376 139776 96440 139780
rect 96456 139836 96520 139840
rect 96456 139780 96460 139836
rect 96460 139780 96516 139836
rect 96516 139780 96520 139836
rect 96456 139776 96520 139780
rect 96536 139836 96600 139840
rect 96536 139780 96540 139836
rect 96540 139780 96596 139836
rect 96596 139780 96600 139836
rect 96536 139776 96600 139780
rect 96616 139836 96680 139840
rect 96616 139780 96620 139836
rect 96620 139780 96676 139836
rect 96676 139780 96680 139836
rect 96616 139776 96680 139780
rect 4876 139292 4940 139296
rect 4876 139236 4880 139292
rect 4880 139236 4936 139292
rect 4936 139236 4940 139292
rect 4876 139232 4940 139236
rect 4956 139292 5020 139296
rect 4956 139236 4960 139292
rect 4960 139236 5016 139292
rect 5016 139236 5020 139292
rect 4956 139232 5020 139236
rect 5036 139292 5100 139296
rect 5036 139236 5040 139292
rect 5040 139236 5096 139292
rect 5096 139236 5100 139292
rect 5036 139232 5100 139236
rect 5116 139292 5180 139296
rect 5116 139236 5120 139292
rect 5120 139236 5176 139292
rect 5176 139236 5180 139292
rect 5116 139232 5180 139236
rect 35596 139292 35660 139296
rect 35596 139236 35600 139292
rect 35600 139236 35656 139292
rect 35656 139236 35660 139292
rect 35596 139232 35660 139236
rect 35676 139292 35740 139296
rect 35676 139236 35680 139292
rect 35680 139236 35736 139292
rect 35736 139236 35740 139292
rect 35676 139232 35740 139236
rect 35756 139292 35820 139296
rect 35756 139236 35760 139292
rect 35760 139236 35816 139292
rect 35816 139236 35820 139292
rect 35756 139232 35820 139236
rect 35836 139292 35900 139296
rect 35836 139236 35840 139292
rect 35840 139236 35896 139292
rect 35896 139236 35900 139292
rect 35836 139232 35900 139236
rect 66316 139292 66380 139296
rect 66316 139236 66320 139292
rect 66320 139236 66376 139292
rect 66376 139236 66380 139292
rect 66316 139232 66380 139236
rect 66396 139292 66460 139296
rect 66396 139236 66400 139292
rect 66400 139236 66456 139292
rect 66456 139236 66460 139292
rect 66396 139232 66460 139236
rect 66476 139292 66540 139296
rect 66476 139236 66480 139292
rect 66480 139236 66536 139292
rect 66536 139236 66540 139292
rect 66476 139232 66540 139236
rect 66556 139292 66620 139296
rect 66556 139236 66560 139292
rect 66560 139236 66616 139292
rect 66616 139236 66620 139292
rect 66556 139232 66620 139236
rect 97036 139292 97100 139296
rect 97036 139236 97040 139292
rect 97040 139236 97096 139292
rect 97096 139236 97100 139292
rect 97036 139232 97100 139236
rect 97116 139292 97180 139296
rect 97116 139236 97120 139292
rect 97120 139236 97176 139292
rect 97176 139236 97180 139292
rect 97116 139232 97180 139236
rect 97196 139292 97260 139296
rect 97196 139236 97200 139292
rect 97200 139236 97256 139292
rect 97256 139236 97260 139292
rect 97196 139232 97260 139236
rect 97276 139292 97340 139296
rect 97276 139236 97280 139292
rect 97280 139236 97336 139292
rect 97336 139236 97340 139292
rect 97276 139232 97340 139236
rect 4216 138748 4280 138752
rect 4216 138692 4220 138748
rect 4220 138692 4276 138748
rect 4276 138692 4280 138748
rect 4216 138688 4280 138692
rect 4296 138748 4360 138752
rect 4296 138692 4300 138748
rect 4300 138692 4356 138748
rect 4356 138692 4360 138748
rect 4296 138688 4360 138692
rect 4376 138748 4440 138752
rect 4376 138692 4380 138748
rect 4380 138692 4436 138748
rect 4436 138692 4440 138748
rect 4376 138688 4440 138692
rect 4456 138748 4520 138752
rect 4456 138692 4460 138748
rect 4460 138692 4516 138748
rect 4516 138692 4520 138748
rect 4456 138688 4520 138692
rect 34936 138748 35000 138752
rect 34936 138692 34940 138748
rect 34940 138692 34996 138748
rect 34996 138692 35000 138748
rect 34936 138688 35000 138692
rect 35016 138748 35080 138752
rect 35016 138692 35020 138748
rect 35020 138692 35076 138748
rect 35076 138692 35080 138748
rect 35016 138688 35080 138692
rect 35096 138748 35160 138752
rect 35096 138692 35100 138748
rect 35100 138692 35156 138748
rect 35156 138692 35160 138748
rect 35096 138688 35160 138692
rect 35176 138748 35240 138752
rect 35176 138692 35180 138748
rect 35180 138692 35236 138748
rect 35236 138692 35240 138748
rect 35176 138688 35240 138692
rect 65656 138748 65720 138752
rect 65656 138692 65660 138748
rect 65660 138692 65716 138748
rect 65716 138692 65720 138748
rect 65656 138688 65720 138692
rect 65736 138748 65800 138752
rect 65736 138692 65740 138748
rect 65740 138692 65796 138748
rect 65796 138692 65800 138748
rect 65736 138688 65800 138692
rect 65816 138748 65880 138752
rect 65816 138692 65820 138748
rect 65820 138692 65876 138748
rect 65876 138692 65880 138748
rect 65816 138688 65880 138692
rect 65896 138748 65960 138752
rect 65896 138692 65900 138748
rect 65900 138692 65956 138748
rect 65956 138692 65960 138748
rect 65896 138688 65960 138692
rect 96376 138748 96440 138752
rect 96376 138692 96380 138748
rect 96380 138692 96436 138748
rect 96436 138692 96440 138748
rect 96376 138688 96440 138692
rect 96456 138748 96520 138752
rect 96456 138692 96460 138748
rect 96460 138692 96516 138748
rect 96516 138692 96520 138748
rect 96456 138688 96520 138692
rect 96536 138748 96600 138752
rect 96536 138692 96540 138748
rect 96540 138692 96596 138748
rect 96596 138692 96600 138748
rect 96536 138688 96600 138692
rect 96616 138748 96680 138752
rect 96616 138692 96620 138748
rect 96620 138692 96676 138748
rect 96676 138692 96680 138748
rect 96616 138688 96680 138692
rect 4876 138204 4940 138208
rect 4876 138148 4880 138204
rect 4880 138148 4936 138204
rect 4936 138148 4940 138204
rect 4876 138144 4940 138148
rect 4956 138204 5020 138208
rect 4956 138148 4960 138204
rect 4960 138148 5016 138204
rect 5016 138148 5020 138204
rect 4956 138144 5020 138148
rect 5036 138204 5100 138208
rect 5036 138148 5040 138204
rect 5040 138148 5096 138204
rect 5096 138148 5100 138204
rect 5036 138144 5100 138148
rect 5116 138204 5180 138208
rect 5116 138148 5120 138204
rect 5120 138148 5176 138204
rect 5176 138148 5180 138204
rect 5116 138144 5180 138148
rect 35596 138204 35660 138208
rect 35596 138148 35600 138204
rect 35600 138148 35656 138204
rect 35656 138148 35660 138204
rect 35596 138144 35660 138148
rect 35676 138204 35740 138208
rect 35676 138148 35680 138204
rect 35680 138148 35736 138204
rect 35736 138148 35740 138204
rect 35676 138144 35740 138148
rect 35756 138204 35820 138208
rect 35756 138148 35760 138204
rect 35760 138148 35816 138204
rect 35816 138148 35820 138204
rect 35756 138144 35820 138148
rect 35836 138204 35900 138208
rect 35836 138148 35840 138204
rect 35840 138148 35896 138204
rect 35896 138148 35900 138204
rect 35836 138144 35900 138148
rect 66316 138204 66380 138208
rect 66316 138148 66320 138204
rect 66320 138148 66376 138204
rect 66376 138148 66380 138204
rect 66316 138144 66380 138148
rect 66396 138204 66460 138208
rect 66396 138148 66400 138204
rect 66400 138148 66456 138204
rect 66456 138148 66460 138204
rect 66396 138144 66460 138148
rect 66476 138204 66540 138208
rect 66476 138148 66480 138204
rect 66480 138148 66536 138204
rect 66536 138148 66540 138204
rect 66476 138144 66540 138148
rect 66556 138204 66620 138208
rect 66556 138148 66560 138204
rect 66560 138148 66616 138204
rect 66616 138148 66620 138204
rect 66556 138144 66620 138148
rect 97036 138204 97100 138208
rect 97036 138148 97040 138204
rect 97040 138148 97096 138204
rect 97096 138148 97100 138204
rect 97036 138144 97100 138148
rect 97116 138204 97180 138208
rect 97116 138148 97120 138204
rect 97120 138148 97176 138204
rect 97176 138148 97180 138204
rect 97116 138144 97180 138148
rect 97196 138204 97260 138208
rect 97196 138148 97200 138204
rect 97200 138148 97256 138204
rect 97256 138148 97260 138204
rect 97196 138144 97260 138148
rect 97276 138204 97340 138208
rect 97276 138148 97280 138204
rect 97280 138148 97336 138204
rect 97336 138148 97340 138204
rect 97276 138144 97340 138148
rect 4216 137660 4280 137664
rect 4216 137604 4220 137660
rect 4220 137604 4276 137660
rect 4276 137604 4280 137660
rect 4216 137600 4280 137604
rect 4296 137660 4360 137664
rect 4296 137604 4300 137660
rect 4300 137604 4356 137660
rect 4356 137604 4360 137660
rect 4296 137600 4360 137604
rect 4376 137660 4440 137664
rect 4376 137604 4380 137660
rect 4380 137604 4436 137660
rect 4436 137604 4440 137660
rect 4376 137600 4440 137604
rect 4456 137660 4520 137664
rect 4456 137604 4460 137660
rect 4460 137604 4516 137660
rect 4516 137604 4520 137660
rect 4456 137600 4520 137604
rect 34936 137660 35000 137664
rect 34936 137604 34940 137660
rect 34940 137604 34996 137660
rect 34996 137604 35000 137660
rect 34936 137600 35000 137604
rect 35016 137660 35080 137664
rect 35016 137604 35020 137660
rect 35020 137604 35076 137660
rect 35076 137604 35080 137660
rect 35016 137600 35080 137604
rect 35096 137660 35160 137664
rect 35096 137604 35100 137660
rect 35100 137604 35156 137660
rect 35156 137604 35160 137660
rect 35096 137600 35160 137604
rect 35176 137660 35240 137664
rect 35176 137604 35180 137660
rect 35180 137604 35236 137660
rect 35236 137604 35240 137660
rect 35176 137600 35240 137604
rect 65656 137660 65720 137664
rect 65656 137604 65660 137660
rect 65660 137604 65716 137660
rect 65716 137604 65720 137660
rect 65656 137600 65720 137604
rect 65736 137660 65800 137664
rect 65736 137604 65740 137660
rect 65740 137604 65796 137660
rect 65796 137604 65800 137660
rect 65736 137600 65800 137604
rect 65816 137660 65880 137664
rect 65816 137604 65820 137660
rect 65820 137604 65876 137660
rect 65876 137604 65880 137660
rect 65816 137600 65880 137604
rect 65896 137660 65960 137664
rect 65896 137604 65900 137660
rect 65900 137604 65956 137660
rect 65956 137604 65960 137660
rect 65896 137600 65960 137604
rect 96376 137660 96440 137664
rect 96376 137604 96380 137660
rect 96380 137604 96436 137660
rect 96436 137604 96440 137660
rect 96376 137600 96440 137604
rect 96456 137660 96520 137664
rect 96456 137604 96460 137660
rect 96460 137604 96516 137660
rect 96516 137604 96520 137660
rect 96456 137600 96520 137604
rect 96536 137660 96600 137664
rect 96536 137604 96540 137660
rect 96540 137604 96596 137660
rect 96596 137604 96600 137660
rect 96536 137600 96600 137604
rect 96616 137660 96680 137664
rect 96616 137604 96620 137660
rect 96620 137604 96676 137660
rect 96676 137604 96680 137660
rect 96616 137600 96680 137604
rect 4876 137116 4940 137120
rect 4876 137060 4880 137116
rect 4880 137060 4936 137116
rect 4936 137060 4940 137116
rect 4876 137056 4940 137060
rect 4956 137116 5020 137120
rect 4956 137060 4960 137116
rect 4960 137060 5016 137116
rect 5016 137060 5020 137116
rect 4956 137056 5020 137060
rect 5036 137116 5100 137120
rect 5036 137060 5040 137116
rect 5040 137060 5096 137116
rect 5096 137060 5100 137116
rect 5036 137056 5100 137060
rect 5116 137116 5180 137120
rect 5116 137060 5120 137116
rect 5120 137060 5176 137116
rect 5176 137060 5180 137116
rect 5116 137056 5180 137060
rect 35596 137116 35660 137120
rect 35596 137060 35600 137116
rect 35600 137060 35656 137116
rect 35656 137060 35660 137116
rect 35596 137056 35660 137060
rect 35676 137116 35740 137120
rect 35676 137060 35680 137116
rect 35680 137060 35736 137116
rect 35736 137060 35740 137116
rect 35676 137056 35740 137060
rect 35756 137116 35820 137120
rect 35756 137060 35760 137116
rect 35760 137060 35816 137116
rect 35816 137060 35820 137116
rect 35756 137056 35820 137060
rect 35836 137116 35900 137120
rect 35836 137060 35840 137116
rect 35840 137060 35896 137116
rect 35896 137060 35900 137116
rect 35836 137056 35900 137060
rect 66316 137116 66380 137120
rect 66316 137060 66320 137116
rect 66320 137060 66376 137116
rect 66376 137060 66380 137116
rect 66316 137056 66380 137060
rect 66396 137116 66460 137120
rect 66396 137060 66400 137116
rect 66400 137060 66456 137116
rect 66456 137060 66460 137116
rect 66396 137056 66460 137060
rect 66476 137116 66540 137120
rect 66476 137060 66480 137116
rect 66480 137060 66536 137116
rect 66536 137060 66540 137116
rect 66476 137056 66540 137060
rect 66556 137116 66620 137120
rect 66556 137060 66560 137116
rect 66560 137060 66616 137116
rect 66616 137060 66620 137116
rect 66556 137056 66620 137060
rect 97036 137116 97100 137120
rect 97036 137060 97040 137116
rect 97040 137060 97096 137116
rect 97096 137060 97100 137116
rect 97036 137056 97100 137060
rect 97116 137116 97180 137120
rect 97116 137060 97120 137116
rect 97120 137060 97176 137116
rect 97176 137060 97180 137116
rect 97116 137056 97180 137060
rect 97196 137116 97260 137120
rect 97196 137060 97200 137116
rect 97200 137060 97256 137116
rect 97256 137060 97260 137116
rect 97196 137056 97260 137060
rect 97276 137116 97340 137120
rect 97276 137060 97280 137116
rect 97280 137060 97336 137116
rect 97336 137060 97340 137116
rect 97276 137056 97340 137060
rect 4216 136572 4280 136576
rect 4216 136516 4220 136572
rect 4220 136516 4276 136572
rect 4276 136516 4280 136572
rect 4216 136512 4280 136516
rect 4296 136572 4360 136576
rect 4296 136516 4300 136572
rect 4300 136516 4356 136572
rect 4356 136516 4360 136572
rect 4296 136512 4360 136516
rect 4376 136572 4440 136576
rect 4376 136516 4380 136572
rect 4380 136516 4436 136572
rect 4436 136516 4440 136572
rect 4376 136512 4440 136516
rect 4456 136572 4520 136576
rect 4456 136516 4460 136572
rect 4460 136516 4516 136572
rect 4516 136516 4520 136572
rect 4456 136512 4520 136516
rect 34936 136572 35000 136576
rect 34936 136516 34940 136572
rect 34940 136516 34996 136572
rect 34996 136516 35000 136572
rect 34936 136512 35000 136516
rect 35016 136572 35080 136576
rect 35016 136516 35020 136572
rect 35020 136516 35076 136572
rect 35076 136516 35080 136572
rect 35016 136512 35080 136516
rect 35096 136572 35160 136576
rect 35096 136516 35100 136572
rect 35100 136516 35156 136572
rect 35156 136516 35160 136572
rect 35096 136512 35160 136516
rect 35176 136572 35240 136576
rect 35176 136516 35180 136572
rect 35180 136516 35236 136572
rect 35236 136516 35240 136572
rect 35176 136512 35240 136516
rect 65656 136572 65720 136576
rect 65656 136516 65660 136572
rect 65660 136516 65716 136572
rect 65716 136516 65720 136572
rect 65656 136512 65720 136516
rect 65736 136572 65800 136576
rect 65736 136516 65740 136572
rect 65740 136516 65796 136572
rect 65796 136516 65800 136572
rect 65736 136512 65800 136516
rect 65816 136572 65880 136576
rect 65816 136516 65820 136572
rect 65820 136516 65876 136572
rect 65876 136516 65880 136572
rect 65816 136512 65880 136516
rect 65896 136572 65960 136576
rect 65896 136516 65900 136572
rect 65900 136516 65956 136572
rect 65956 136516 65960 136572
rect 65896 136512 65960 136516
rect 96376 136572 96440 136576
rect 96376 136516 96380 136572
rect 96380 136516 96436 136572
rect 96436 136516 96440 136572
rect 96376 136512 96440 136516
rect 96456 136572 96520 136576
rect 96456 136516 96460 136572
rect 96460 136516 96516 136572
rect 96516 136516 96520 136572
rect 96456 136512 96520 136516
rect 96536 136572 96600 136576
rect 96536 136516 96540 136572
rect 96540 136516 96596 136572
rect 96596 136516 96600 136572
rect 96536 136512 96600 136516
rect 96616 136572 96680 136576
rect 96616 136516 96620 136572
rect 96620 136516 96676 136572
rect 96676 136516 96680 136572
rect 96616 136512 96680 136516
rect 105924 136572 105988 136576
rect 105924 136516 105928 136572
rect 105928 136516 105984 136572
rect 105984 136516 105988 136572
rect 105924 136512 105988 136516
rect 106004 136572 106068 136576
rect 106004 136516 106008 136572
rect 106008 136516 106064 136572
rect 106064 136516 106068 136572
rect 106004 136512 106068 136516
rect 106084 136572 106148 136576
rect 106084 136516 106088 136572
rect 106088 136516 106144 136572
rect 106144 136516 106148 136572
rect 106084 136512 106148 136516
rect 106164 136572 106228 136576
rect 106164 136516 106168 136572
rect 106168 136516 106224 136572
rect 106224 136516 106228 136572
rect 106164 136512 106228 136516
rect 4876 136028 4940 136032
rect 4876 135972 4880 136028
rect 4880 135972 4936 136028
rect 4936 135972 4940 136028
rect 4876 135968 4940 135972
rect 4956 136028 5020 136032
rect 4956 135972 4960 136028
rect 4960 135972 5016 136028
rect 5016 135972 5020 136028
rect 4956 135968 5020 135972
rect 5036 136028 5100 136032
rect 5036 135972 5040 136028
rect 5040 135972 5096 136028
rect 5096 135972 5100 136028
rect 5036 135968 5100 135972
rect 5116 136028 5180 136032
rect 5116 135972 5120 136028
rect 5120 135972 5176 136028
rect 5176 135972 5180 136028
rect 5116 135968 5180 135972
rect 35596 136028 35660 136032
rect 35596 135972 35600 136028
rect 35600 135972 35656 136028
rect 35656 135972 35660 136028
rect 35596 135968 35660 135972
rect 35676 136028 35740 136032
rect 35676 135972 35680 136028
rect 35680 135972 35736 136028
rect 35736 135972 35740 136028
rect 35676 135968 35740 135972
rect 35756 136028 35820 136032
rect 35756 135972 35760 136028
rect 35760 135972 35816 136028
rect 35816 135972 35820 136028
rect 35756 135968 35820 135972
rect 35836 136028 35900 136032
rect 35836 135972 35840 136028
rect 35840 135972 35896 136028
rect 35896 135972 35900 136028
rect 35836 135968 35900 135972
rect 66316 136028 66380 136032
rect 66316 135972 66320 136028
rect 66320 135972 66376 136028
rect 66376 135972 66380 136028
rect 66316 135968 66380 135972
rect 66396 136028 66460 136032
rect 66396 135972 66400 136028
rect 66400 135972 66456 136028
rect 66456 135972 66460 136028
rect 66396 135968 66460 135972
rect 66476 136028 66540 136032
rect 66476 135972 66480 136028
rect 66480 135972 66536 136028
rect 66536 135972 66540 136028
rect 66476 135968 66540 135972
rect 66556 136028 66620 136032
rect 66556 135972 66560 136028
rect 66560 135972 66616 136028
rect 66616 135972 66620 136028
rect 66556 135968 66620 135972
rect 97036 136028 97100 136032
rect 97036 135972 97040 136028
rect 97040 135972 97096 136028
rect 97096 135972 97100 136028
rect 97036 135968 97100 135972
rect 97116 136028 97180 136032
rect 97116 135972 97120 136028
rect 97120 135972 97176 136028
rect 97176 135972 97180 136028
rect 97116 135968 97180 135972
rect 97196 136028 97260 136032
rect 97196 135972 97200 136028
rect 97200 135972 97256 136028
rect 97256 135972 97260 136028
rect 97196 135968 97260 135972
rect 97276 136028 97340 136032
rect 97276 135972 97280 136028
rect 97280 135972 97336 136028
rect 97336 135972 97340 136028
rect 97276 135968 97340 135972
rect 106660 136028 106724 136032
rect 106660 135972 106664 136028
rect 106664 135972 106720 136028
rect 106720 135972 106724 136028
rect 106660 135968 106724 135972
rect 106740 136028 106804 136032
rect 106740 135972 106744 136028
rect 106744 135972 106800 136028
rect 106800 135972 106804 136028
rect 106740 135968 106804 135972
rect 106820 136028 106884 136032
rect 106820 135972 106824 136028
rect 106824 135972 106880 136028
rect 106880 135972 106884 136028
rect 106820 135968 106884 135972
rect 106900 136028 106964 136032
rect 106900 135972 106904 136028
rect 106904 135972 106960 136028
rect 106960 135972 106964 136028
rect 106900 135968 106964 135972
rect 4216 135484 4280 135488
rect 4216 135428 4220 135484
rect 4220 135428 4276 135484
rect 4276 135428 4280 135484
rect 4216 135424 4280 135428
rect 4296 135484 4360 135488
rect 4296 135428 4300 135484
rect 4300 135428 4356 135484
rect 4356 135428 4360 135484
rect 4296 135424 4360 135428
rect 4376 135484 4440 135488
rect 4376 135428 4380 135484
rect 4380 135428 4436 135484
rect 4436 135428 4440 135484
rect 4376 135424 4440 135428
rect 4456 135484 4520 135488
rect 4456 135428 4460 135484
rect 4460 135428 4516 135484
rect 4516 135428 4520 135484
rect 4456 135424 4520 135428
rect 105924 135484 105988 135488
rect 105924 135428 105928 135484
rect 105928 135428 105984 135484
rect 105984 135428 105988 135484
rect 105924 135424 105988 135428
rect 106004 135484 106068 135488
rect 106004 135428 106008 135484
rect 106008 135428 106064 135484
rect 106064 135428 106068 135484
rect 106004 135424 106068 135428
rect 106084 135484 106148 135488
rect 106084 135428 106088 135484
rect 106088 135428 106144 135484
rect 106144 135428 106148 135484
rect 106084 135424 106148 135428
rect 106164 135484 106228 135488
rect 106164 135428 106168 135484
rect 106168 135428 106224 135484
rect 106224 135428 106228 135484
rect 106164 135424 106228 135428
rect 58572 135220 58636 135284
rect 61148 135220 61212 135284
rect 66116 135220 66180 135284
rect 68508 135220 68572 135284
rect 71084 135220 71148 135284
rect 63540 135084 63604 135148
rect 4876 134940 4940 134944
rect 4876 134884 4880 134940
rect 4880 134884 4936 134940
rect 4936 134884 4940 134940
rect 4876 134880 4940 134884
rect 4956 134940 5020 134944
rect 4956 134884 4960 134940
rect 4960 134884 5016 134940
rect 5016 134884 5020 134940
rect 4956 134880 5020 134884
rect 5036 134940 5100 134944
rect 5036 134884 5040 134940
rect 5040 134884 5096 134940
rect 5096 134884 5100 134940
rect 5036 134880 5100 134884
rect 5116 134940 5180 134944
rect 5116 134884 5120 134940
rect 5120 134884 5176 134940
rect 5176 134884 5180 134940
rect 5116 134880 5180 134884
rect 106660 134940 106724 134944
rect 106660 134884 106664 134940
rect 106664 134884 106720 134940
rect 106720 134884 106724 134940
rect 106660 134880 106724 134884
rect 106740 134940 106804 134944
rect 106740 134884 106744 134940
rect 106744 134884 106800 134940
rect 106800 134884 106804 134940
rect 106740 134880 106804 134884
rect 106820 134940 106884 134944
rect 106820 134884 106824 134940
rect 106824 134884 106880 134940
rect 106880 134884 106884 134940
rect 106820 134880 106884 134884
rect 106900 134940 106964 134944
rect 106900 134884 106904 134940
rect 106904 134884 106960 134940
rect 106960 134884 106964 134940
rect 106900 134880 106964 134884
rect 95924 134464 95988 134468
rect 95924 134408 95974 134464
rect 95974 134408 95988 134464
rect 95924 134404 95988 134408
rect 4216 134396 4280 134400
rect 4216 134340 4220 134396
rect 4220 134340 4276 134396
rect 4276 134340 4280 134396
rect 4216 134336 4280 134340
rect 4296 134396 4360 134400
rect 4296 134340 4300 134396
rect 4300 134340 4356 134396
rect 4356 134340 4360 134396
rect 4296 134336 4360 134340
rect 4376 134396 4440 134400
rect 4376 134340 4380 134396
rect 4380 134340 4436 134396
rect 4436 134340 4440 134396
rect 4376 134336 4440 134340
rect 4456 134396 4520 134400
rect 4456 134340 4460 134396
rect 4460 134340 4516 134396
rect 4516 134340 4520 134396
rect 4456 134336 4520 134340
rect 105924 134396 105988 134400
rect 105924 134340 105928 134396
rect 105928 134340 105984 134396
rect 105984 134340 105988 134396
rect 105924 134336 105988 134340
rect 106004 134396 106068 134400
rect 106004 134340 106008 134396
rect 106008 134340 106064 134396
rect 106064 134340 106068 134396
rect 106004 134336 106068 134340
rect 106084 134396 106148 134400
rect 106084 134340 106088 134396
rect 106088 134340 106144 134396
rect 106144 134340 106148 134396
rect 106084 134336 106148 134340
rect 106164 134396 106228 134400
rect 106164 134340 106168 134396
rect 106168 134340 106224 134396
rect 106224 134340 106228 134396
rect 106164 134336 106228 134340
rect 38571 134132 38635 134196
rect 41067 134132 41131 134196
rect 51051 134132 51115 134196
rect 56043 134132 56107 134196
rect 73515 134132 73579 134196
rect 53547 133996 53611 134060
rect 36075 133920 36139 133924
rect 36075 133864 36082 133920
rect 36082 133864 36138 133920
rect 36138 133864 36139 133920
rect 36075 133860 36139 133864
rect 43563 133860 43627 133924
rect 46059 133920 46123 133924
rect 46059 133864 46074 133920
rect 46074 133864 46123 133920
rect 46059 133860 46123 133864
rect 48544 133920 48608 133924
rect 48544 133864 48558 133920
rect 48558 133864 48608 133920
rect 48544 133860 48608 133864
rect 86142 133920 86206 133924
rect 86142 133864 86186 133920
rect 86186 133864 86206 133920
rect 86142 133860 86206 133864
rect 87310 133920 87374 133924
rect 87310 133864 87326 133920
rect 87326 133864 87374 133920
rect 87310 133860 87374 133864
rect 4876 133852 4940 133856
rect 4876 133796 4880 133852
rect 4880 133796 4936 133852
rect 4936 133796 4940 133852
rect 4876 133792 4940 133796
rect 4956 133852 5020 133856
rect 4956 133796 4960 133852
rect 4960 133796 5016 133852
rect 5016 133796 5020 133852
rect 4956 133792 5020 133796
rect 5036 133852 5100 133856
rect 5036 133796 5040 133852
rect 5040 133796 5096 133852
rect 5096 133796 5100 133852
rect 5036 133792 5100 133796
rect 5116 133852 5180 133856
rect 5116 133796 5120 133852
rect 5120 133796 5176 133852
rect 5176 133796 5180 133852
rect 5116 133792 5180 133796
rect 106660 133852 106724 133856
rect 106660 133796 106664 133852
rect 106664 133796 106720 133852
rect 106720 133796 106724 133852
rect 106660 133792 106724 133796
rect 106740 133852 106804 133856
rect 106740 133796 106744 133852
rect 106744 133796 106800 133852
rect 106800 133796 106804 133852
rect 106740 133792 106804 133796
rect 106820 133852 106884 133856
rect 106820 133796 106824 133852
rect 106824 133796 106880 133852
rect 106880 133796 106884 133852
rect 106820 133792 106884 133796
rect 106900 133852 106964 133856
rect 106900 133796 106904 133852
rect 106904 133796 106960 133852
rect 106960 133796 106964 133852
rect 106900 133792 106964 133796
rect 4216 133308 4280 133312
rect 4216 133252 4220 133308
rect 4220 133252 4276 133308
rect 4276 133252 4280 133308
rect 4216 133248 4280 133252
rect 4296 133308 4360 133312
rect 4296 133252 4300 133308
rect 4300 133252 4356 133308
rect 4356 133252 4360 133308
rect 4296 133248 4360 133252
rect 4376 133308 4440 133312
rect 4376 133252 4380 133308
rect 4380 133252 4436 133308
rect 4436 133252 4440 133308
rect 4376 133248 4440 133252
rect 4456 133308 4520 133312
rect 4456 133252 4460 133308
rect 4460 133252 4516 133308
rect 4516 133252 4520 133308
rect 4456 133248 4520 133252
rect 105924 133308 105988 133312
rect 105924 133252 105928 133308
rect 105928 133252 105984 133308
rect 105984 133252 105988 133308
rect 105924 133248 105988 133252
rect 106004 133308 106068 133312
rect 106004 133252 106008 133308
rect 106008 133252 106064 133308
rect 106064 133252 106068 133308
rect 106004 133248 106068 133252
rect 106084 133308 106148 133312
rect 106084 133252 106088 133308
rect 106088 133252 106144 133308
rect 106144 133252 106148 133308
rect 106084 133248 106148 133252
rect 106164 133308 106228 133312
rect 106164 133252 106168 133308
rect 106168 133252 106224 133308
rect 106224 133252 106228 133308
rect 106164 133248 106228 133252
rect 4876 132764 4940 132768
rect 4876 132708 4880 132764
rect 4880 132708 4936 132764
rect 4936 132708 4940 132764
rect 4876 132704 4940 132708
rect 4956 132764 5020 132768
rect 4956 132708 4960 132764
rect 4960 132708 5016 132764
rect 5016 132708 5020 132764
rect 4956 132704 5020 132708
rect 5036 132764 5100 132768
rect 5036 132708 5040 132764
rect 5040 132708 5096 132764
rect 5096 132708 5100 132764
rect 5036 132704 5100 132708
rect 5116 132764 5180 132768
rect 5116 132708 5120 132764
rect 5120 132708 5176 132764
rect 5176 132708 5180 132764
rect 5116 132704 5180 132708
rect 106660 132764 106724 132768
rect 106660 132708 106664 132764
rect 106664 132708 106720 132764
rect 106720 132708 106724 132764
rect 106660 132704 106724 132708
rect 106740 132764 106804 132768
rect 106740 132708 106744 132764
rect 106744 132708 106800 132764
rect 106800 132708 106804 132764
rect 106740 132704 106804 132708
rect 106820 132764 106884 132768
rect 106820 132708 106824 132764
rect 106824 132708 106880 132764
rect 106880 132708 106884 132764
rect 106820 132704 106884 132708
rect 106900 132764 106964 132768
rect 106900 132708 106904 132764
rect 106904 132708 106960 132764
rect 106960 132708 106964 132764
rect 106900 132704 106964 132708
rect 4216 132220 4280 132224
rect 4216 132164 4220 132220
rect 4220 132164 4276 132220
rect 4276 132164 4280 132220
rect 4216 132160 4280 132164
rect 4296 132220 4360 132224
rect 4296 132164 4300 132220
rect 4300 132164 4356 132220
rect 4356 132164 4360 132220
rect 4296 132160 4360 132164
rect 4376 132220 4440 132224
rect 4376 132164 4380 132220
rect 4380 132164 4436 132220
rect 4436 132164 4440 132220
rect 4376 132160 4440 132164
rect 4456 132220 4520 132224
rect 4456 132164 4460 132220
rect 4460 132164 4516 132220
rect 4516 132164 4520 132220
rect 4456 132160 4520 132164
rect 105924 132220 105988 132224
rect 105924 132164 105928 132220
rect 105928 132164 105984 132220
rect 105984 132164 105988 132220
rect 105924 132160 105988 132164
rect 106004 132220 106068 132224
rect 106004 132164 106008 132220
rect 106008 132164 106064 132220
rect 106064 132164 106068 132220
rect 106004 132160 106068 132164
rect 106084 132220 106148 132224
rect 106084 132164 106088 132220
rect 106088 132164 106144 132220
rect 106144 132164 106148 132220
rect 106084 132160 106148 132164
rect 106164 132220 106228 132224
rect 106164 132164 106168 132220
rect 106168 132164 106224 132220
rect 106224 132164 106228 132220
rect 106164 132160 106228 132164
rect 4876 131676 4940 131680
rect 4876 131620 4880 131676
rect 4880 131620 4936 131676
rect 4936 131620 4940 131676
rect 4876 131616 4940 131620
rect 4956 131676 5020 131680
rect 4956 131620 4960 131676
rect 4960 131620 5016 131676
rect 5016 131620 5020 131676
rect 4956 131616 5020 131620
rect 5036 131676 5100 131680
rect 5036 131620 5040 131676
rect 5040 131620 5096 131676
rect 5096 131620 5100 131676
rect 5036 131616 5100 131620
rect 5116 131676 5180 131680
rect 5116 131620 5120 131676
rect 5120 131620 5176 131676
rect 5176 131620 5180 131676
rect 5116 131616 5180 131620
rect 106660 131676 106724 131680
rect 106660 131620 106664 131676
rect 106664 131620 106720 131676
rect 106720 131620 106724 131676
rect 106660 131616 106724 131620
rect 106740 131676 106804 131680
rect 106740 131620 106744 131676
rect 106744 131620 106800 131676
rect 106800 131620 106804 131676
rect 106740 131616 106804 131620
rect 106820 131676 106884 131680
rect 106820 131620 106824 131676
rect 106824 131620 106880 131676
rect 106880 131620 106884 131676
rect 106820 131616 106884 131620
rect 106900 131676 106964 131680
rect 106900 131620 106904 131676
rect 106904 131620 106960 131676
rect 106960 131620 106964 131676
rect 106900 131616 106964 131620
rect 4216 131132 4280 131136
rect 4216 131076 4220 131132
rect 4220 131076 4276 131132
rect 4276 131076 4280 131132
rect 4216 131072 4280 131076
rect 4296 131132 4360 131136
rect 4296 131076 4300 131132
rect 4300 131076 4356 131132
rect 4356 131076 4360 131132
rect 4296 131072 4360 131076
rect 4376 131132 4440 131136
rect 4376 131076 4380 131132
rect 4380 131076 4436 131132
rect 4436 131076 4440 131132
rect 4376 131072 4440 131076
rect 4456 131132 4520 131136
rect 4456 131076 4460 131132
rect 4460 131076 4516 131132
rect 4516 131076 4520 131132
rect 4456 131072 4520 131076
rect 105924 131132 105988 131136
rect 105924 131076 105928 131132
rect 105928 131076 105984 131132
rect 105984 131076 105988 131132
rect 105924 131072 105988 131076
rect 106004 131132 106068 131136
rect 106004 131076 106008 131132
rect 106008 131076 106064 131132
rect 106064 131076 106068 131132
rect 106004 131072 106068 131076
rect 106084 131132 106148 131136
rect 106084 131076 106088 131132
rect 106088 131076 106144 131132
rect 106144 131076 106148 131132
rect 106084 131072 106148 131076
rect 106164 131132 106228 131136
rect 106164 131076 106168 131132
rect 106168 131076 106224 131132
rect 106224 131076 106228 131132
rect 106164 131072 106228 131076
rect 4876 130588 4940 130592
rect 4876 130532 4880 130588
rect 4880 130532 4936 130588
rect 4936 130532 4940 130588
rect 4876 130528 4940 130532
rect 4956 130588 5020 130592
rect 4956 130532 4960 130588
rect 4960 130532 5016 130588
rect 5016 130532 5020 130588
rect 4956 130528 5020 130532
rect 5036 130588 5100 130592
rect 5036 130532 5040 130588
rect 5040 130532 5096 130588
rect 5096 130532 5100 130588
rect 5036 130528 5100 130532
rect 5116 130588 5180 130592
rect 5116 130532 5120 130588
rect 5120 130532 5176 130588
rect 5176 130532 5180 130588
rect 5116 130528 5180 130532
rect 106660 130588 106724 130592
rect 106660 130532 106664 130588
rect 106664 130532 106720 130588
rect 106720 130532 106724 130588
rect 106660 130528 106724 130532
rect 106740 130588 106804 130592
rect 106740 130532 106744 130588
rect 106744 130532 106800 130588
rect 106800 130532 106804 130588
rect 106740 130528 106804 130532
rect 106820 130588 106884 130592
rect 106820 130532 106824 130588
rect 106824 130532 106880 130588
rect 106880 130532 106884 130588
rect 106820 130528 106884 130532
rect 106900 130588 106964 130592
rect 106900 130532 106904 130588
rect 106904 130532 106960 130588
rect 106960 130532 106964 130588
rect 106900 130528 106964 130532
rect 4216 130044 4280 130048
rect 4216 129988 4220 130044
rect 4220 129988 4276 130044
rect 4276 129988 4280 130044
rect 4216 129984 4280 129988
rect 4296 130044 4360 130048
rect 4296 129988 4300 130044
rect 4300 129988 4356 130044
rect 4356 129988 4360 130044
rect 4296 129984 4360 129988
rect 4376 130044 4440 130048
rect 4376 129988 4380 130044
rect 4380 129988 4436 130044
rect 4436 129988 4440 130044
rect 4376 129984 4440 129988
rect 4456 130044 4520 130048
rect 4456 129988 4460 130044
rect 4460 129988 4516 130044
rect 4516 129988 4520 130044
rect 4456 129984 4520 129988
rect 105924 130044 105988 130048
rect 105924 129988 105928 130044
rect 105928 129988 105984 130044
rect 105984 129988 105988 130044
rect 105924 129984 105988 129988
rect 106004 130044 106068 130048
rect 106004 129988 106008 130044
rect 106008 129988 106064 130044
rect 106064 129988 106068 130044
rect 106004 129984 106068 129988
rect 106084 130044 106148 130048
rect 106084 129988 106088 130044
rect 106088 129988 106144 130044
rect 106144 129988 106148 130044
rect 106084 129984 106148 129988
rect 106164 130044 106228 130048
rect 106164 129988 106168 130044
rect 106168 129988 106224 130044
rect 106224 129988 106228 130044
rect 106164 129984 106228 129988
rect 4876 129500 4940 129504
rect 4876 129444 4880 129500
rect 4880 129444 4936 129500
rect 4936 129444 4940 129500
rect 4876 129440 4940 129444
rect 4956 129500 5020 129504
rect 4956 129444 4960 129500
rect 4960 129444 5016 129500
rect 5016 129444 5020 129500
rect 4956 129440 5020 129444
rect 5036 129500 5100 129504
rect 5036 129444 5040 129500
rect 5040 129444 5096 129500
rect 5096 129444 5100 129500
rect 5036 129440 5100 129444
rect 5116 129500 5180 129504
rect 5116 129444 5120 129500
rect 5120 129444 5176 129500
rect 5176 129444 5180 129500
rect 5116 129440 5180 129444
rect 106660 129500 106724 129504
rect 106660 129444 106664 129500
rect 106664 129444 106720 129500
rect 106720 129444 106724 129500
rect 106660 129440 106724 129444
rect 106740 129500 106804 129504
rect 106740 129444 106744 129500
rect 106744 129444 106800 129500
rect 106800 129444 106804 129500
rect 106740 129440 106804 129444
rect 106820 129500 106884 129504
rect 106820 129444 106824 129500
rect 106824 129444 106880 129500
rect 106880 129444 106884 129500
rect 106820 129440 106884 129444
rect 106900 129500 106964 129504
rect 106900 129444 106904 129500
rect 106904 129444 106960 129500
rect 106960 129444 106964 129500
rect 106900 129440 106964 129444
rect 4216 128956 4280 128960
rect 4216 128900 4220 128956
rect 4220 128900 4276 128956
rect 4276 128900 4280 128956
rect 4216 128896 4280 128900
rect 4296 128956 4360 128960
rect 4296 128900 4300 128956
rect 4300 128900 4356 128956
rect 4356 128900 4360 128956
rect 4296 128896 4360 128900
rect 4376 128956 4440 128960
rect 4376 128900 4380 128956
rect 4380 128900 4436 128956
rect 4436 128900 4440 128956
rect 4376 128896 4440 128900
rect 4456 128956 4520 128960
rect 4456 128900 4460 128956
rect 4460 128900 4516 128956
rect 4516 128900 4520 128956
rect 4456 128896 4520 128900
rect 105924 128956 105988 128960
rect 105924 128900 105928 128956
rect 105928 128900 105984 128956
rect 105984 128900 105988 128956
rect 105924 128896 105988 128900
rect 106004 128956 106068 128960
rect 106004 128900 106008 128956
rect 106008 128900 106064 128956
rect 106064 128900 106068 128956
rect 106004 128896 106068 128900
rect 106084 128956 106148 128960
rect 106084 128900 106088 128956
rect 106088 128900 106144 128956
rect 106144 128900 106148 128956
rect 106084 128896 106148 128900
rect 106164 128956 106228 128960
rect 106164 128900 106168 128956
rect 106168 128900 106224 128956
rect 106224 128900 106228 128956
rect 106164 128896 106228 128900
rect 4876 128412 4940 128416
rect 4876 128356 4880 128412
rect 4880 128356 4936 128412
rect 4936 128356 4940 128412
rect 4876 128352 4940 128356
rect 4956 128412 5020 128416
rect 4956 128356 4960 128412
rect 4960 128356 5016 128412
rect 5016 128356 5020 128412
rect 4956 128352 5020 128356
rect 5036 128412 5100 128416
rect 5036 128356 5040 128412
rect 5040 128356 5096 128412
rect 5096 128356 5100 128412
rect 5036 128352 5100 128356
rect 5116 128412 5180 128416
rect 5116 128356 5120 128412
rect 5120 128356 5176 128412
rect 5176 128356 5180 128412
rect 5116 128352 5180 128356
rect 106660 128412 106724 128416
rect 106660 128356 106664 128412
rect 106664 128356 106720 128412
rect 106720 128356 106724 128412
rect 106660 128352 106724 128356
rect 106740 128412 106804 128416
rect 106740 128356 106744 128412
rect 106744 128356 106800 128412
rect 106800 128356 106804 128412
rect 106740 128352 106804 128356
rect 106820 128412 106884 128416
rect 106820 128356 106824 128412
rect 106824 128356 106880 128412
rect 106880 128356 106884 128412
rect 106820 128352 106884 128356
rect 106900 128412 106964 128416
rect 106900 128356 106904 128412
rect 106904 128356 106960 128412
rect 106960 128356 106964 128412
rect 106900 128352 106964 128356
rect 4216 127868 4280 127872
rect 4216 127812 4220 127868
rect 4220 127812 4276 127868
rect 4276 127812 4280 127868
rect 4216 127808 4280 127812
rect 4296 127868 4360 127872
rect 4296 127812 4300 127868
rect 4300 127812 4356 127868
rect 4356 127812 4360 127868
rect 4296 127808 4360 127812
rect 4376 127868 4440 127872
rect 4376 127812 4380 127868
rect 4380 127812 4436 127868
rect 4436 127812 4440 127868
rect 4376 127808 4440 127812
rect 4456 127868 4520 127872
rect 4456 127812 4460 127868
rect 4460 127812 4516 127868
rect 4516 127812 4520 127868
rect 4456 127808 4520 127812
rect 105924 127868 105988 127872
rect 105924 127812 105928 127868
rect 105928 127812 105984 127868
rect 105984 127812 105988 127868
rect 105924 127808 105988 127812
rect 106004 127868 106068 127872
rect 106004 127812 106008 127868
rect 106008 127812 106064 127868
rect 106064 127812 106068 127868
rect 106004 127808 106068 127812
rect 106084 127868 106148 127872
rect 106084 127812 106088 127868
rect 106088 127812 106144 127868
rect 106144 127812 106148 127868
rect 106084 127808 106148 127812
rect 106164 127868 106228 127872
rect 106164 127812 106168 127868
rect 106168 127812 106224 127868
rect 106224 127812 106228 127868
rect 106164 127808 106228 127812
rect 4876 127324 4940 127328
rect 4876 127268 4880 127324
rect 4880 127268 4936 127324
rect 4936 127268 4940 127324
rect 4876 127264 4940 127268
rect 4956 127324 5020 127328
rect 4956 127268 4960 127324
rect 4960 127268 5016 127324
rect 5016 127268 5020 127324
rect 4956 127264 5020 127268
rect 5036 127324 5100 127328
rect 5036 127268 5040 127324
rect 5040 127268 5096 127324
rect 5096 127268 5100 127324
rect 5036 127264 5100 127268
rect 5116 127324 5180 127328
rect 5116 127268 5120 127324
rect 5120 127268 5176 127324
rect 5176 127268 5180 127324
rect 5116 127264 5180 127268
rect 106660 127324 106724 127328
rect 106660 127268 106664 127324
rect 106664 127268 106720 127324
rect 106720 127268 106724 127324
rect 106660 127264 106724 127268
rect 106740 127324 106804 127328
rect 106740 127268 106744 127324
rect 106744 127268 106800 127324
rect 106800 127268 106804 127324
rect 106740 127264 106804 127268
rect 106820 127324 106884 127328
rect 106820 127268 106824 127324
rect 106824 127268 106880 127324
rect 106880 127268 106884 127324
rect 106820 127264 106884 127268
rect 106900 127324 106964 127328
rect 106900 127268 106904 127324
rect 106904 127268 106960 127324
rect 106960 127268 106964 127324
rect 106900 127264 106964 127268
rect 4216 126780 4280 126784
rect 4216 126724 4220 126780
rect 4220 126724 4276 126780
rect 4276 126724 4280 126780
rect 4216 126720 4280 126724
rect 4296 126780 4360 126784
rect 4296 126724 4300 126780
rect 4300 126724 4356 126780
rect 4356 126724 4360 126780
rect 4296 126720 4360 126724
rect 4376 126780 4440 126784
rect 4376 126724 4380 126780
rect 4380 126724 4436 126780
rect 4436 126724 4440 126780
rect 4376 126720 4440 126724
rect 4456 126780 4520 126784
rect 4456 126724 4460 126780
rect 4460 126724 4516 126780
rect 4516 126724 4520 126780
rect 4456 126720 4520 126724
rect 105924 126780 105988 126784
rect 105924 126724 105928 126780
rect 105928 126724 105984 126780
rect 105984 126724 105988 126780
rect 105924 126720 105988 126724
rect 106004 126780 106068 126784
rect 106004 126724 106008 126780
rect 106008 126724 106064 126780
rect 106064 126724 106068 126780
rect 106004 126720 106068 126724
rect 106084 126780 106148 126784
rect 106084 126724 106088 126780
rect 106088 126724 106144 126780
rect 106144 126724 106148 126780
rect 106084 126720 106148 126724
rect 106164 126780 106228 126784
rect 106164 126724 106168 126780
rect 106168 126724 106224 126780
rect 106224 126724 106228 126780
rect 106164 126720 106228 126724
rect 4876 126236 4940 126240
rect 4876 126180 4880 126236
rect 4880 126180 4936 126236
rect 4936 126180 4940 126236
rect 4876 126176 4940 126180
rect 4956 126236 5020 126240
rect 4956 126180 4960 126236
rect 4960 126180 5016 126236
rect 5016 126180 5020 126236
rect 4956 126176 5020 126180
rect 5036 126236 5100 126240
rect 5036 126180 5040 126236
rect 5040 126180 5096 126236
rect 5096 126180 5100 126236
rect 5036 126176 5100 126180
rect 5116 126236 5180 126240
rect 5116 126180 5120 126236
rect 5120 126180 5176 126236
rect 5176 126180 5180 126236
rect 5116 126176 5180 126180
rect 106660 126236 106724 126240
rect 106660 126180 106664 126236
rect 106664 126180 106720 126236
rect 106720 126180 106724 126236
rect 106660 126176 106724 126180
rect 106740 126236 106804 126240
rect 106740 126180 106744 126236
rect 106744 126180 106800 126236
rect 106800 126180 106804 126236
rect 106740 126176 106804 126180
rect 106820 126236 106884 126240
rect 106820 126180 106824 126236
rect 106824 126180 106880 126236
rect 106880 126180 106884 126236
rect 106820 126176 106884 126180
rect 106900 126236 106964 126240
rect 106900 126180 106904 126236
rect 106904 126180 106960 126236
rect 106960 126180 106964 126236
rect 106900 126176 106964 126180
rect 4216 125692 4280 125696
rect 4216 125636 4220 125692
rect 4220 125636 4276 125692
rect 4276 125636 4280 125692
rect 4216 125632 4280 125636
rect 4296 125692 4360 125696
rect 4296 125636 4300 125692
rect 4300 125636 4356 125692
rect 4356 125636 4360 125692
rect 4296 125632 4360 125636
rect 4376 125692 4440 125696
rect 4376 125636 4380 125692
rect 4380 125636 4436 125692
rect 4436 125636 4440 125692
rect 4376 125632 4440 125636
rect 4456 125692 4520 125696
rect 4456 125636 4460 125692
rect 4460 125636 4516 125692
rect 4516 125636 4520 125692
rect 4456 125632 4520 125636
rect 105924 125692 105988 125696
rect 105924 125636 105928 125692
rect 105928 125636 105984 125692
rect 105984 125636 105988 125692
rect 105924 125632 105988 125636
rect 106004 125692 106068 125696
rect 106004 125636 106008 125692
rect 106008 125636 106064 125692
rect 106064 125636 106068 125692
rect 106004 125632 106068 125636
rect 106084 125692 106148 125696
rect 106084 125636 106088 125692
rect 106088 125636 106144 125692
rect 106144 125636 106148 125692
rect 106084 125632 106148 125636
rect 106164 125692 106228 125696
rect 106164 125636 106168 125692
rect 106168 125636 106224 125692
rect 106224 125636 106228 125692
rect 106164 125632 106228 125636
rect 4876 125148 4940 125152
rect 4876 125092 4880 125148
rect 4880 125092 4936 125148
rect 4936 125092 4940 125148
rect 4876 125088 4940 125092
rect 4956 125148 5020 125152
rect 4956 125092 4960 125148
rect 4960 125092 5016 125148
rect 5016 125092 5020 125148
rect 4956 125088 5020 125092
rect 5036 125148 5100 125152
rect 5036 125092 5040 125148
rect 5040 125092 5096 125148
rect 5096 125092 5100 125148
rect 5036 125088 5100 125092
rect 5116 125148 5180 125152
rect 5116 125092 5120 125148
rect 5120 125092 5176 125148
rect 5176 125092 5180 125148
rect 5116 125088 5180 125092
rect 106660 125148 106724 125152
rect 106660 125092 106664 125148
rect 106664 125092 106720 125148
rect 106720 125092 106724 125148
rect 106660 125088 106724 125092
rect 106740 125148 106804 125152
rect 106740 125092 106744 125148
rect 106744 125092 106800 125148
rect 106800 125092 106804 125148
rect 106740 125088 106804 125092
rect 106820 125148 106884 125152
rect 106820 125092 106824 125148
rect 106824 125092 106880 125148
rect 106880 125092 106884 125148
rect 106820 125088 106884 125092
rect 106900 125148 106964 125152
rect 106900 125092 106904 125148
rect 106904 125092 106960 125148
rect 106960 125092 106964 125148
rect 106900 125088 106964 125092
rect 4216 124604 4280 124608
rect 4216 124548 4220 124604
rect 4220 124548 4276 124604
rect 4276 124548 4280 124604
rect 4216 124544 4280 124548
rect 4296 124604 4360 124608
rect 4296 124548 4300 124604
rect 4300 124548 4356 124604
rect 4356 124548 4360 124604
rect 4296 124544 4360 124548
rect 4376 124604 4440 124608
rect 4376 124548 4380 124604
rect 4380 124548 4436 124604
rect 4436 124548 4440 124604
rect 4376 124544 4440 124548
rect 4456 124604 4520 124608
rect 4456 124548 4460 124604
rect 4460 124548 4516 124604
rect 4516 124548 4520 124604
rect 4456 124544 4520 124548
rect 105924 124604 105988 124608
rect 105924 124548 105928 124604
rect 105928 124548 105984 124604
rect 105984 124548 105988 124604
rect 105924 124544 105988 124548
rect 106004 124604 106068 124608
rect 106004 124548 106008 124604
rect 106008 124548 106064 124604
rect 106064 124548 106068 124604
rect 106004 124544 106068 124548
rect 106084 124604 106148 124608
rect 106084 124548 106088 124604
rect 106088 124548 106144 124604
rect 106144 124548 106148 124604
rect 106084 124544 106148 124548
rect 106164 124604 106228 124608
rect 106164 124548 106168 124604
rect 106168 124548 106224 124604
rect 106224 124548 106228 124604
rect 106164 124544 106228 124548
rect 4876 124060 4940 124064
rect 4876 124004 4880 124060
rect 4880 124004 4936 124060
rect 4936 124004 4940 124060
rect 4876 124000 4940 124004
rect 4956 124060 5020 124064
rect 4956 124004 4960 124060
rect 4960 124004 5016 124060
rect 5016 124004 5020 124060
rect 4956 124000 5020 124004
rect 5036 124060 5100 124064
rect 5036 124004 5040 124060
rect 5040 124004 5096 124060
rect 5096 124004 5100 124060
rect 5036 124000 5100 124004
rect 5116 124060 5180 124064
rect 5116 124004 5120 124060
rect 5120 124004 5176 124060
rect 5176 124004 5180 124060
rect 5116 124000 5180 124004
rect 106660 124060 106724 124064
rect 106660 124004 106664 124060
rect 106664 124004 106720 124060
rect 106720 124004 106724 124060
rect 106660 124000 106724 124004
rect 106740 124060 106804 124064
rect 106740 124004 106744 124060
rect 106744 124004 106800 124060
rect 106800 124004 106804 124060
rect 106740 124000 106804 124004
rect 106820 124060 106884 124064
rect 106820 124004 106824 124060
rect 106824 124004 106880 124060
rect 106880 124004 106884 124060
rect 106820 124000 106884 124004
rect 106900 124060 106964 124064
rect 106900 124004 106904 124060
rect 106904 124004 106960 124060
rect 106960 124004 106964 124060
rect 106900 124000 106964 124004
rect 4216 123516 4280 123520
rect 4216 123460 4220 123516
rect 4220 123460 4276 123516
rect 4276 123460 4280 123516
rect 4216 123456 4280 123460
rect 4296 123516 4360 123520
rect 4296 123460 4300 123516
rect 4300 123460 4356 123516
rect 4356 123460 4360 123516
rect 4296 123456 4360 123460
rect 4376 123516 4440 123520
rect 4376 123460 4380 123516
rect 4380 123460 4436 123516
rect 4436 123460 4440 123516
rect 4376 123456 4440 123460
rect 4456 123516 4520 123520
rect 4456 123460 4460 123516
rect 4460 123460 4516 123516
rect 4516 123460 4520 123516
rect 4456 123456 4520 123460
rect 105924 123516 105988 123520
rect 105924 123460 105928 123516
rect 105928 123460 105984 123516
rect 105984 123460 105988 123516
rect 105924 123456 105988 123460
rect 106004 123516 106068 123520
rect 106004 123460 106008 123516
rect 106008 123460 106064 123516
rect 106064 123460 106068 123516
rect 106004 123456 106068 123460
rect 106084 123516 106148 123520
rect 106084 123460 106088 123516
rect 106088 123460 106144 123516
rect 106144 123460 106148 123516
rect 106084 123456 106148 123460
rect 106164 123516 106228 123520
rect 106164 123460 106168 123516
rect 106168 123460 106224 123516
rect 106224 123460 106228 123516
rect 106164 123456 106228 123460
rect 4876 122972 4940 122976
rect 4876 122916 4880 122972
rect 4880 122916 4936 122972
rect 4936 122916 4940 122972
rect 4876 122912 4940 122916
rect 4956 122972 5020 122976
rect 4956 122916 4960 122972
rect 4960 122916 5016 122972
rect 5016 122916 5020 122972
rect 4956 122912 5020 122916
rect 5036 122972 5100 122976
rect 5036 122916 5040 122972
rect 5040 122916 5096 122972
rect 5096 122916 5100 122972
rect 5036 122912 5100 122916
rect 5116 122972 5180 122976
rect 5116 122916 5120 122972
rect 5120 122916 5176 122972
rect 5176 122916 5180 122972
rect 5116 122912 5180 122916
rect 106660 122972 106724 122976
rect 106660 122916 106664 122972
rect 106664 122916 106720 122972
rect 106720 122916 106724 122972
rect 106660 122912 106724 122916
rect 106740 122972 106804 122976
rect 106740 122916 106744 122972
rect 106744 122916 106800 122972
rect 106800 122916 106804 122972
rect 106740 122912 106804 122916
rect 106820 122972 106884 122976
rect 106820 122916 106824 122972
rect 106824 122916 106880 122972
rect 106880 122916 106884 122972
rect 106820 122912 106884 122916
rect 106900 122972 106964 122976
rect 106900 122916 106904 122972
rect 106904 122916 106960 122972
rect 106960 122916 106964 122972
rect 106900 122912 106964 122916
rect 4216 122428 4280 122432
rect 4216 122372 4220 122428
rect 4220 122372 4276 122428
rect 4276 122372 4280 122428
rect 4216 122368 4280 122372
rect 4296 122428 4360 122432
rect 4296 122372 4300 122428
rect 4300 122372 4356 122428
rect 4356 122372 4360 122428
rect 4296 122368 4360 122372
rect 4376 122428 4440 122432
rect 4376 122372 4380 122428
rect 4380 122372 4436 122428
rect 4436 122372 4440 122428
rect 4376 122368 4440 122372
rect 4456 122428 4520 122432
rect 4456 122372 4460 122428
rect 4460 122372 4516 122428
rect 4516 122372 4520 122428
rect 4456 122368 4520 122372
rect 105924 122428 105988 122432
rect 105924 122372 105928 122428
rect 105928 122372 105984 122428
rect 105984 122372 105988 122428
rect 105924 122368 105988 122372
rect 106004 122428 106068 122432
rect 106004 122372 106008 122428
rect 106008 122372 106064 122428
rect 106064 122372 106068 122428
rect 106004 122368 106068 122372
rect 106084 122428 106148 122432
rect 106084 122372 106088 122428
rect 106088 122372 106144 122428
rect 106144 122372 106148 122428
rect 106084 122368 106148 122372
rect 106164 122428 106228 122432
rect 106164 122372 106168 122428
rect 106168 122372 106224 122428
rect 106224 122372 106228 122428
rect 106164 122368 106228 122372
rect 4876 121884 4940 121888
rect 4876 121828 4880 121884
rect 4880 121828 4936 121884
rect 4936 121828 4940 121884
rect 4876 121824 4940 121828
rect 4956 121884 5020 121888
rect 4956 121828 4960 121884
rect 4960 121828 5016 121884
rect 5016 121828 5020 121884
rect 4956 121824 5020 121828
rect 5036 121884 5100 121888
rect 5036 121828 5040 121884
rect 5040 121828 5096 121884
rect 5096 121828 5100 121884
rect 5036 121824 5100 121828
rect 5116 121884 5180 121888
rect 5116 121828 5120 121884
rect 5120 121828 5176 121884
rect 5176 121828 5180 121884
rect 5116 121824 5180 121828
rect 106660 121884 106724 121888
rect 106660 121828 106664 121884
rect 106664 121828 106720 121884
rect 106720 121828 106724 121884
rect 106660 121824 106724 121828
rect 106740 121884 106804 121888
rect 106740 121828 106744 121884
rect 106744 121828 106800 121884
rect 106800 121828 106804 121884
rect 106740 121824 106804 121828
rect 106820 121884 106884 121888
rect 106820 121828 106824 121884
rect 106824 121828 106880 121884
rect 106880 121828 106884 121884
rect 106820 121824 106884 121828
rect 106900 121884 106964 121888
rect 106900 121828 106904 121884
rect 106904 121828 106960 121884
rect 106960 121828 106964 121884
rect 106900 121824 106964 121828
rect 4216 121340 4280 121344
rect 4216 121284 4220 121340
rect 4220 121284 4276 121340
rect 4276 121284 4280 121340
rect 4216 121280 4280 121284
rect 4296 121340 4360 121344
rect 4296 121284 4300 121340
rect 4300 121284 4356 121340
rect 4356 121284 4360 121340
rect 4296 121280 4360 121284
rect 4376 121340 4440 121344
rect 4376 121284 4380 121340
rect 4380 121284 4436 121340
rect 4436 121284 4440 121340
rect 4376 121280 4440 121284
rect 4456 121340 4520 121344
rect 4456 121284 4460 121340
rect 4460 121284 4516 121340
rect 4516 121284 4520 121340
rect 4456 121280 4520 121284
rect 105924 121340 105988 121344
rect 105924 121284 105928 121340
rect 105928 121284 105984 121340
rect 105984 121284 105988 121340
rect 105924 121280 105988 121284
rect 106004 121340 106068 121344
rect 106004 121284 106008 121340
rect 106008 121284 106064 121340
rect 106064 121284 106068 121340
rect 106004 121280 106068 121284
rect 106084 121340 106148 121344
rect 106084 121284 106088 121340
rect 106088 121284 106144 121340
rect 106144 121284 106148 121340
rect 106084 121280 106148 121284
rect 106164 121340 106228 121344
rect 106164 121284 106168 121340
rect 106168 121284 106224 121340
rect 106224 121284 106228 121340
rect 106164 121280 106228 121284
rect 4876 120796 4940 120800
rect 4876 120740 4880 120796
rect 4880 120740 4936 120796
rect 4936 120740 4940 120796
rect 4876 120736 4940 120740
rect 4956 120796 5020 120800
rect 4956 120740 4960 120796
rect 4960 120740 5016 120796
rect 5016 120740 5020 120796
rect 4956 120736 5020 120740
rect 5036 120796 5100 120800
rect 5036 120740 5040 120796
rect 5040 120740 5096 120796
rect 5096 120740 5100 120796
rect 5036 120736 5100 120740
rect 5116 120796 5180 120800
rect 5116 120740 5120 120796
rect 5120 120740 5176 120796
rect 5176 120740 5180 120796
rect 5116 120736 5180 120740
rect 106660 120796 106724 120800
rect 106660 120740 106664 120796
rect 106664 120740 106720 120796
rect 106720 120740 106724 120796
rect 106660 120736 106724 120740
rect 106740 120796 106804 120800
rect 106740 120740 106744 120796
rect 106744 120740 106800 120796
rect 106800 120740 106804 120796
rect 106740 120736 106804 120740
rect 106820 120796 106884 120800
rect 106820 120740 106824 120796
rect 106824 120740 106880 120796
rect 106880 120740 106884 120796
rect 106820 120736 106884 120740
rect 106900 120796 106964 120800
rect 106900 120740 106904 120796
rect 106904 120740 106960 120796
rect 106960 120740 106964 120796
rect 106900 120736 106964 120740
rect 4216 120252 4280 120256
rect 4216 120196 4220 120252
rect 4220 120196 4276 120252
rect 4276 120196 4280 120252
rect 4216 120192 4280 120196
rect 4296 120252 4360 120256
rect 4296 120196 4300 120252
rect 4300 120196 4356 120252
rect 4356 120196 4360 120252
rect 4296 120192 4360 120196
rect 4376 120252 4440 120256
rect 4376 120196 4380 120252
rect 4380 120196 4436 120252
rect 4436 120196 4440 120252
rect 4376 120192 4440 120196
rect 4456 120252 4520 120256
rect 4456 120196 4460 120252
rect 4460 120196 4516 120252
rect 4516 120196 4520 120252
rect 4456 120192 4520 120196
rect 105924 120252 105988 120256
rect 105924 120196 105928 120252
rect 105928 120196 105984 120252
rect 105984 120196 105988 120252
rect 105924 120192 105988 120196
rect 106004 120252 106068 120256
rect 106004 120196 106008 120252
rect 106008 120196 106064 120252
rect 106064 120196 106068 120252
rect 106004 120192 106068 120196
rect 106084 120252 106148 120256
rect 106084 120196 106088 120252
rect 106088 120196 106144 120252
rect 106144 120196 106148 120252
rect 106084 120192 106148 120196
rect 106164 120252 106228 120256
rect 106164 120196 106168 120252
rect 106168 120196 106224 120252
rect 106224 120196 106228 120252
rect 106164 120192 106228 120196
rect 4876 119708 4940 119712
rect 4876 119652 4880 119708
rect 4880 119652 4936 119708
rect 4936 119652 4940 119708
rect 4876 119648 4940 119652
rect 4956 119708 5020 119712
rect 4956 119652 4960 119708
rect 4960 119652 5016 119708
rect 5016 119652 5020 119708
rect 4956 119648 5020 119652
rect 5036 119708 5100 119712
rect 5036 119652 5040 119708
rect 5040 119652 5096 119708
rect 5096 119652 5100 119708
rect 5036 119648 5100 119652
rect 5116 119708 5180 119712
rect 5116 119652 5120 119708
rect 5120 119652 5176 119708
rect 5176 119652 5180 119708
rect 5116 119648 5180 119652
rect 106660 119708 106724 119712
rect 106660 119652 106664 119708
rect 106664 119652 106720 119708
rect 106720 119652 106724 119708
rect 106660 119648 106724 119652
rect 106740 119708 106804 119712
rect 106740 119652 106744 119708
rect 106744 119652 106800 119708
rect 106800 119652 106804 119708
rect 106740 119648 106804 119652
rect 106820 119708 106884 119712
rect 106820 119652 106824 119708
rect 106824 119652 106880 119708
rect 106880 119652 106884 119708
rect 106820 119648 106884 119652
rect 106900 119708 106964 119712
rect 106900 119652 106904 119708
rect 106904 119652 106960 119708
rect 106960 119652 106964 119708
rect 106900 119648 106964 119652
rect 4216 119164 4280 119168
rect 4216 119108 4220 119164
rect 4220 119108 4276 119164
rect 4276 119108 4280 119164
rect 4216 119104 4280 119108
rect 4296 119164 4360 119168
rect 4296 119108 4300 119164
rect 4300 119108 4356 119164
rect 4356 119108 4360 119164
rect 4296 119104 4360 119108
rect 4376 119164 4440 119168
rect 4376 119108 4380 119164
rect 4380 119108 4436 119164
rect 4436 119108 4440 119164
rect 4376 119104 4440 119108
rect 4456 119164 4520 119168
rect 4456 119108 4460 119164
rect 4460 119108 4516 119164
rect 4516 119108 4520 119164
rect 4456 119104 4520 119108
rect 105924 119164 105988 119168
rect 105924 119108 105928 119164
rect 105928 119108 105984 119164
rect 105984 119108 105988 119164
rect 105924 119104 105988 119108
rect 106004 119164 106068 119168
rect 106004 119108 106008 119164
rect 106008 119108 106064 119164
rect 106064 119108 106068 119164
rect 106004 119104 106068 119108
rect 106084 119164 106148 119168
rect 106084 119108 106088 119164
rect 106088 119108 106144 119164
rect 106144 119108 106148 119164
rect 106084 119104 106148 119108
rect 106164 119164 106228 119168
rect 106164 119108 106168 119164
rect 106168 119108 106224 119164
rect 106224 119108 106228 119164
rect 106164 119104 106228 119108
rect 4876 118620 4940 118624
rect 4876 118564 4880 118620
rect 4880 118564 4936 118620
rect 4936 118564 4940 118620
rect 4876 118560 4940 118564
rect 4956 118620 5020 118624
rect 4956 118564 4960 118620
rect 4960 118564 5016 118620
rect 5016 118564 5020 118620
rect 4956 118560 5020 118564
rect 5036 118620 5100 118624
rect 5036 118564 5040 118620
rect 5040 118564 5096 118620
rect 5096 118564 5100 118620
rect 5036 118560 5100 118564
rect 5116 118620 5180 118624
rect 5116 118564 5120 118620
rect 5120 118564 5176 118620
rect 5176 118564 5180 118620
rect 5116 118560 5180 118564
rect 106660 118620 106724 118624
rect 106660 118564 106664 118620
rect 106664 118564 106720 118620
rect 106720 118564 106724 118620
rect 106660 118560 106724 118564
rect 106740 118620 106804 118624
rect 106740 118564 106744 118620
rect 106744 118564 106800 118620
rect 106800 118564 106804 118620
rect 106740 118560 106804 118564
rect 106820 118620 106884 118624
rect 106820 118564 106824 118620
rect 106824 118564 106880 118620
rect 106880 118564 106884 118620
rect 106820 118560 106884 118564
rect 106900 118620 106964 118624
rect 106900 118564 106904 118620
rect 106904 118564 106960 118620
rect 106960 118564 106964 118620
rect 106900 118560 106964 118564
rect 4216 118076 4280 118080
rect 4216 118020 4220 118076
rect 4220 118020 4276 118076
rect 4276 118020 4280 118076
rect 4216 118016 4280 118020
rect 4296 118076 4360 118080
rect 4296 118020 4300 118076
rect 4300 118020 4356 118076
rect 4356 118020 4360 118076
rect 4296 118016 4360 118020
rect 4376 118076 4440 118080
rect 4376 118020 4380 118076
rect 4380 118020 4436 118076
rect 4436 118020 4440 118076
rect 4376 118016 4440 118020
rect 4456 118076 4520 118080
rect 4456 118020 4460 118076
rect 4460 118020 4516 118076
rect 4516 118020 4520 118076
rect 4456 118016 4520 118020
rect 105924 118076 105988 118080
rect 105924 118020 105928 118076
rect 105928 118020 105984 118076
rect 105984 118020 105988 118076
rect 105924 118016 105988 118020
rect 106004 118076 106068 118080
rect 106004 118020 106008 118076
rect 106008 118020 106064 118076
rect 106064 118020 106068 118076
rect 106004 118016 106068 118020
rect 106084 118076 106148 118080
rect 106084 118020 106088 118076
rect 106088 118020 106144 118076
rect 106144 118020 106148 118076
rect 106084 118016 106148 118020
rect 106164 118076 106228 118080
rect 106164 118020 106168 118076
rect 106168 118020 106224 118076
rect 106224 118020 106228 118076
rect 106164 118016 106228 118020
rect 4876 117532 4940 117536
rect 4876 117476 4880 117532
rect 4880 117476 4936 117532
rect 4936 117476 4940 117532
rect 4876 117472 4940 117476
rect 4956 117532 5020 117536
rect 4956 117476 4960 117532
rect 4960 117476 5016 117532
rect 5016 117476 5020 117532
rect 4956 117472 5020 117476
rect 5036 117532 5100 117536
rect 5036 117476 5040 117532
rect 5040 117476 5096 117532
rect 5096 117476 5100 117532
rect 5036 117472 5100 117476
rect 5116 117532 5180 117536
rect 5116 117476 5120 117532
rect 5120 117476 5176 117532
rect 5176 117476 5180 117532
rect 5116 117472 5180 117476
rect 106660 117532 106724 117536
rect 106660 117476 106664 117532
rect 106664 117476 106720 117532
rect 106720 117476 106724 117532
rect 106660 117472 106724 117476
rect 106740 117532 106804 117536
rect 106740 117476 106744 117532
rect 106744 117476 106800 117532
rect 106800 117476 106804 117532
rect 106740 117472 106804 117476
rect 106820 117532 106884 117536
rect 106820 117476 106824 117532
rect 106824 117476 106880 117532
rect 106880 117476 106884 117532
rect 106820 117472 106884 117476
rect 106900 117532 106964 117536
rect 106900 117476 106904 117532
rect 106904 117476 106960 117532
rect 106960 117476 106964 117532
rect 106900 117472 106964 117476
rect 4216 116988 4280 116992
rect 4216 116932 4220 116988
rect 4220 116932 4276 116988
rect 4276 116932 4280 116988
rect 4216 116928 4280 116932
rect 4296 116988 4360 116992
rect 4296 116932 4300 116988
rect 4300 116932 4356 116988
rect 4356 116932 4360 116988
rect 4296 116928 4360 116932
rect 4376 116988 4440 116992
rect 4376 116932 4380 116988
rect 4380 116932 4436 116988
rect 4436 116932 4440 116988
rect 4376 116928 4440 116932
rect 4456 116988 4520 116992
rect 4456 116932 4460 116988
rect 4460 116932 4516 116988
rect 4516 116932 4520 116988
rect 4456 116928 4520 116932
rect 105924 116988 105988 116992
rect 105924 116932 105928 116988
rect 105928 116932 105984 116988
rect 105984 116932 105988 116988
rect 105924 116928 105988 116932
rect 106004 116988 106068 116992
rect 106004 116932 106008 116988
rect 106008 116932 106064 116988
rect 106064 116932 106068 116988
rect 106004 116928 106068 116932
rect 106084 116988 106148 116992
rect 106084 116932 106088 116988
rect 106088 116932 106144 116988
rect 106144 116932 106148 116988
rect 106084 116928 106148 116932
rect 106164 116988 106228 116992
rect 106164 116932 106168 116988
rect 106168 116932 106224 116988
rect 106224 116932 106228 116988
rect 106164 116928 106228 116932
rect 4876 116444 4940 116448
rect 4876 116388 4880 116444
rect 4880 116388 4936 116444
rect 4936 116388 4940 116444
rect 4876 116384 4940 116388
rect 4956 116444 5020 116448
rect 4956 116388 4960 116444
rect 4960 116388 5016 116444
rect 5016 116388 5020 116444
rect 4956 116384 5020 116388
rect 5036 116444 5100 116448
rect 5036 116388 5040 116444
rect 5040 116388 5096 116444
rect 5096 116388 5100 116444
rect 5036 116384 5100 116388
rect 5116 116444 5180 116448
rect 5116 116388 5120 116444
rect 5120 116388 5176 116444
rect 5176 116388 5180 116444
rect 5116 116384 5180 116388
rect 106660 116444 106724 116448
rect 106660 116388 106664 116444
rect 106664 116388 106720 116444
rect 106720 116388 106724 116444
rect 106660 116384 106724 116388
rect 106740 116444 106804 116448
rect 106740 116388 106744 116444
rect 106744 116388 106800 116444
rect 106800 116388 106804 116444
rect 106740 116384 106804 116388
rect 106820 116444 106884 116448
rect 106820 116388 106824 116444
rect 106824 116388 106880 116444
rect 106880 116388 106884 116444
rect 106820 116384 106884 116388
rect 106900 116444 106964 116448
rect 106900 116388 106904 116444
rect 106904 116388 106960 116444
rect 106960 116388 106964 116444
rect 106900 116384 106964 116388
rect 4216 115900 4280 115904
rect 4216 115844 4220 115900
rect 4220 115844 4276 115900
rect 4276 115844 4280 115900
rect 4216 115840 4280 115844
rect 4296 115900 4360 115904
rect 4296 115844 4300 115900
rect 4300 115844 4356 115900
rect 4356 115844 4360 115900
rect 4296 115840 4360 115844
rect 4376 115900 4440 115904
rect 4376 115844 4380 115900
rect 4380 115844 4436 115900
rect 4436 115844 4440 115900
rect 4376 115840 4440 115844
rect 4456 115900 4520 115904
rect 4456 115844 4460 115900
rect 4460 115844 4516 115900
rect 4516 115844 4520 115900
rect 4456 115840 4520 115844
rect 105924 115900 105988 115904
rect 105924 115844 105928 115900
rect 105928 115844 105984 115900
rect 105984 115844 105988 115900
rect 105924 115840 105988 115844
rect 106004 115900 106068 115904
rect 106004 115844 106008 115900
rect 106008 115844 106064 115900
rect 106064 115844 106068 115900
rect 106004 115840 106068 115844
rect 106084 115900 106148 115904
rect 106084 115844 106088 115900
rect 106088 115844 106144 115900
rect 106144 115844 106148 115900
rect 106084 115840 106148 115844
rect 106164 115900 106228 115904
rect 106164 115844 106168 115900
rect 106168 115844 106224 115900
rect 106224 115844 106228 115900
rect 106164 115840 106228 115844
rect 4876 115356 4940 115360
rect 4876 115300 4880 115356
rect 4880 115300 4936 115356
rect 4936 115300 4940 115356
rect 4876 115296 4940 115300
rect 4956 115356 5020 115360
rect 4956 115300 4960 115356
rect 4960 115300 5016 115356
rect 5016 115300 5020 115356
rect 4956 115296 5020 115300
rect 5036 115356 5100 115360
rect 5036 115300 5040 115356
rect 5040 115300 5096 115356
rect 5096 115300 5100 115356
rect 5036 115296 5100 115300
rect 5116 115356 5180 115360
rect 5116 115300 5120 115356
rect 5120 115300 5176 115356
rect 5176 115300 5180 115356
rect 5116 115296 5180 115300
rect 106660 115356 106724 115360
rect 106660 115300 106664 115356
rect 106664 115300 106720 115356
rect 106720 115300 106724 115356
rect 106660 115296 106724 115300
rect 106740 115356 106804 115360
rect 106740 115300 106744 115356
rect 106744 115300 106800 115356
rect 106800 115300 106804 115356
rect 106740 115296 106804 115300
rect 106820 115356 106884 115360
rect 106820 115300 106824 115356
rect 106824 115300 106880 115356
rect 106880 115300 106884 115356
rect 106820 115296 106884 115300
rect 106900 115356 106964 115360
rect 106900 115300 106904 115356
rect 106904 115300 106960 115356
rect 106960 115300 106964 115356
rect 106900 115296 106964 115300
rect 4216 114812 4280 114816
rect 4216 114756 4220 114812
rect 4220 114756 4276 114812
rect 4276 114756 4280 114812
rect 4216 114752 4280 114756
rect 4296 114812 4360 114816
rect 4296 114756 4300 114812
rect 4300 114756 4356 114812
rect 4356 114756 4360 114812
rect 4296 114752 4360 114756
rect 4376 114812 4440 114816
rect 4376 114756 4380 114812
rect 4380 114756 4436 114812
rect 4436 114756 4440 114812
rect 4376 114752 4440 114756
rect 4456 114812 4520 114816
rect 4456 114756 4460 114812
rect 4460 114756 4516 114812
rect 4516 114756 4520 114812
rect 4456 114752 4520 114756
rect 105924 114812 105988 114816
rect 105924 114756 105928 114812
rect 105928 114756 105984 114812
rect 105984 114756 105988 114812
rect 105924 114752 105988 114756
rect 106004 114812 106068 114816
rect 106004 114756 106008 114812
rect 106008 114756 106064 114812
rect 106064 114756 106068 114812
rect 106004 114752 106068 114756
rect 106084 114812 106148 114816
rect 106084 114756 106088 114812
rect 106088 114756 106144 114812
rect 106144 114756 106148 114812
rect 106084 114752 106148 114756
rect 106164 114812 106228 114816
rect 106164 114756 106168 114812
rect 106168 114756 106224 114812
rect 106224 114756 106228 114812
rect 106164 114752 106228 114756
rect 4876 114268 4940 114272
rect 4876 114212 4880 114268
rect 4880 114212 4936 114268
rect 4936 114212 4940 114268
rect 4876 114208 4940 114212
rect 4956 114268 5020 114272
rect 4956 114212 4960 114268
rect 4960 114212 5016 114268
rect 5016 114212 5020 114268
rect 4956 114208 5020 114212
rect 5036 114268 5100 114272
rect 5036 114212 5040 114268
rect 5040 114212 5096 114268
rect 5096 114212 5100 114268
rect 5036 114208 5100 114212
rect 5116 114268 5180 114272
rect 5116 114212 5120 114268
rect 5120 114212 5176 114268
rect 5176 114212 5180 114268
rect 5116 114208 5180 114212
rect 106660 114268 106724 114272
rect 106660 114212 106664 114268
rect 106664 114212 106720 114268
rect 106720 114212 106724 114268
rect 106660 114208 106724 114212
rect 106740 114268 106804 114272
rect 106740 114212 106744 114268
rect 106744 114212 106800 114268
rect 106800 114212 106804 114268
rect 106740 114208 106804 114212
rect 106820 114268 106884 114272
rect 106820 114212 106824 114268
rect 106824 114212 106880 114268
rect 106880 114212 106884 114268
rect 106820 114208 106884 114212
rect 106900 114268 106964 114272
rect 106900 114212 106904 114268
rect 106904 114212 106960 114268
rect 106960 114212 106964 114268
rect 106900 114208 106964 114212
rect 4216 113724 4280 113728
rect 4216 113668 4220 113724
rect 4220 113668 4276 113724
rect 4276 113668 4280 113724
rect 4216 113664 4280 113668
rect 4296 113724 4360 113728
rect 4296 113668 4300 113724
rect 4300 113668 4356 113724
rect 4356 113668 4360 113724
rect 4296 113664 4360 113668
rect 4376 113724 4440 113728
rect 4376 113668 4380 113724
rect 4380 113668 4436 113724
rect 4436 113668 4440 113724
rect 4376 113664 4440 113668
rect 4456 113724 4520 113728
rect 4456 113668 4460 113724
rect 4460 113668 4516 113724
rect 4516 113668 4520 113724
rect 4456 113664 4520 113668
rect 105924 113724 105988 113728
rect 105924 113668 105928 113724
rect 105928 113668 105984 113724
rect 105984 113668 105988 113724
rect 105924 113664 105988 113668
rect 106004 113724 106068 113728
rect 106004 113668 106008 113724
rect 106008 113668 106064 113724
rect 106064 113668 106068 113724
rect 106004 113664 106068 113668
rect 106084 113724 106148 113728
rect 106084 113668 106088 113724
rect 106088 113668 106144 113724
rect 106144 113668 106148 113724
rect 106084 113664 106148 113668
rect 106164 113724 106228 113728
rect 106164 113668 106168 113724
rect 106168 113668 106224 113724
rect 106224 113668 106228 113724
rect 106164 113664 106228 113668
rect 4876 113180 4940 113184
rect 4876 113124 4880 113180
rect 4880 113124 4936 113180
rect 4936 113124 4940 113180
rect 4876 113120 4940 113124
rect 4956 113180 5020 113184
rect 4956 113124 4960 113180
rect 4960 113124 5016 113180
rect 5016 113124 5020 113180
rect 4956 113120 5020 113124
rect 5036 113180 5100 113184
rect 5036 113124 5040 113180
rect 5040 113124 5096 113180
rect 5096 113124 5100 113180
rect 5036 113120 5100 113124
rect 5116 113180 5180 113184
rect 5116 113124 5120 113180
rect 5120 113124 5176 113180
rect 5176 113124 5180 113180
rect 5116 113120 5180 113124
rect 106660 113180 106724 113184
rect 106660 113124 106664 113180
rect 106664 113124 106720 113180
rect 106720 113124 106724 113180
rect 106660 113120 106724 113124
rect 106740 113180 106804 113184
rect 106740 113124 106744 113180
rect 106744 113124 106800 113180
rect 106800 113124 106804 113180
rect 106740 113120 106804 113124
rect 106820 113180 106884 113184
rect 106820 113124 106824 113180
rect 106824 113124 106880 113180
rect 106880 113124 106884 113180
rect 106820 113120 106884 113124
rect 106900 113180 106964 113184
rect 106900 113124 106904 113180
rect 106904 113124 106960 113180
rect 106960 113124 106964 113180
rect 106900 113120 106964 113124
rect 4216 112636 4280 112640
rect 4216 112580 4220 112636
rect 4220 112580 4276 112636
rect 4276 112580 4280 112636
rect 4216 112576 4280 112580
rect 4296 112636 4360 112640
rect 4296 112580 4300 112636
rect 4300 112580 4356 112636
rect 4356 112580 4360 112636
rect 4296 112576 4360 112580
rect 4376 112636 4440 112640
rect 4376 112580 4380 112636
rect 4380 112580 4436 112636
rect 4436 112580 4440 112636
rect 4376 112576 4440 112580
rect 4456 112636 4520 112640
rect 4456 112580 4460 112636
rect 4460 112580 4516 112636
rect 4516 112580 4520 112636
rect 4456 112576 4520 112580
rect 105924 112636 105988 112640
rect 105924 112580 105928 112636
rect 105928 112580 105984 112636
rect 105984 112580 105988 112636
rect 105924 112576 105988 112580
rect 106004 112636 106068 112640
rect 106004 112580 106008 112636
rect 106008 112580 106064 112636
rect 106064 112580 106068 112636
rect 106004 112576 106068 112580
rect 106084 112636 106148 112640
rect 106084 112580 106088 112636
rect 106088 112580 106144 112636
rect 106144 112580 106148 112636
rect 106084 112576 106148 112580
rect 106164 112636 106228 112640
rect 106164 112580 106168 112636
rect 106168 112580 106224 112636
rect 106224 112580 106228 112636
rect 106164 112576 106228 112580
rect 4876 112092 4940 112096
rect 4876 112036 4880 112092
rect 4880 112036 4936 112092
rect 4936 112036 4940 112092
rect 4876 112032 4940 112036
rect 4956 112092 5020 112096
rect 4956 112036 4960 112092
rect 4960 112036 5016 112092
rect 5016 112036 5020 112092
rect 4956 112032 5020 112036
rect 5036 112092 5100 112096
rect 5036 112036 5040 112092
rect 5040 112036 5096 112092
rect 5096 112036 5100 112092
rect 5036 112032 5100 112036
rect 5116 112092 5180 112096
rect 5116 112036 5120 112092
rect 5120 112036 5176 112092
rect 5176 112036 5180 112092
rect 5116 112032 5180 112036
rect 106660 112092 106724 112096
rect 106660 112036 106664 112092
rect 106664 112036 106720 112092
rect 106720 112036 106724 112092
rect 106660 112032 106724 112036
rect 106740 112092 106804 112096
rect 106740 112036 106744 112092
rect 106744 112036 106800 112092
rect 106800 112036 106804 112092
rect 106740 112032 106804 112036
rect 106820 112092 106884 112096
rect 106820 112036 106824 112092
rect 106824 112036 106880 112092
rect 106880 112036 106884 112092
rect 106820 112032 106884 112036
rect 106900 112092 106964 112096
rect 106900 112036 106904 112092
rect 106904 112036 106960 112092
rect 106960 112036 106964 112092
rect 106900 112032 106964 112036
rect 4216 111548 4280 111552
rect 4216 111492 4220 111548
rect 4220 111492 4276 111548
rect 4276 111492 4280 111548
rect 4216 111488 4280 111492
rect 4296 111548 4360 111552
rect 4296 111492 4300 111548
rect 4300 111492 4356 111548
rect 4356 111492 4360 111548
rect 4296 111488 4360 111492
rect 4376 111548 4440 111552
rect 4376 111492 4380 111548
rect 4380 111492 4436 111548
rect 4436 111492 4440 111548
rect 4376 111488 4440 111492
rect 4456 111548 4520 111552
rect 4456 111492 4460 111548
rect 4460 111492 4516 111548
rect 4516 111492 4520 111548
rect 4456 111488 4520 111492
rect 105924 111548 105988 111552
rect 105924 111492 105928 111548
rect 105928 111492 105984 111548
rect 105984 111492 105988 111548
rect 105924 111488 105988 111492
rect 106004 111548 106068 111552
rect 106004 111492 106008 111548
rect 106008 111492 106064 111548
rect 106064 111492 106068 111548
rect 106004 111488 106068 111492
rect 106084 111548 106148 111552
rect 106084 111492 106088 111548
rect 106088 111492 106144 111548
rect 106144 111492 106148 111548
rect 106084 111488 106148 111492
rect 106164 111548 106228 111552
rect 106164 111492 106168 111548
rect 106168 111492 106224 111548
rect 106224 111492 106228 111548
rect 106164 111488 106228 111492
rect 4876 111004 4940 111008
rect 4876 110948 4880 111004
rect 4880 110948 4936 111004
rect 4936 110948 4940 111004
rect 4876 110944 4940 110948
rect 4956 111004 5020 111008
rect 4956 110948 4960 111004
rect 4960 110948 5016 111004
rect 5016 110948 5020 111004
rect 4956 110944 5020 110948
rect 5036 111004 5100 111008
rect 5036 110948 5040 111004
rect 5040 110948 5096 111004
rect 5096 110948 5100 111004
rect 5036 110944 5100 110948
rect 5116 111004 5180 111008
rect 5116 110948 5120 111004
rect 5120 110948 5176 111004
rect 5176 110948 5180 111004
rect 5116 110944 5180 110948
rect 106660 111004 106724 111008
rect 106660 110948 106664 111004
rect 106664 110948 106720 111004
rect 106720 110948 106724 111004
rect 106660 110944 106724 110948
rect 106740 111004 106804 111008
rect 106740 110948 106744 111004
rect 106744 110948 106800 111004
rect 106800 110948 106804 111004
rect 106740 110944 106804 110948
rect 106820 111004 106884 111008
rect 106820 110948 106824 111004
rect 106824 110948 106880 111004
rect 106880 110948 106884 111004
rect 106820 110944 106884 110948
rect 106900 111004 106964 111008
rect 106900 110948 106904 111004
rect 106904 110948 106960 111004
rect 106960 110948 106964 111004
rect 106900 110944 106964 110948
rect 4216 110460 4280 110464
rect 4216 110404 4220 110460
rect 4220 110404 4276 110460
rect 4276 110404 4280 110460
rect 4216 110400 4280 110404
rect 4296 110460 4360 110464
rect 4296 110404 4300 110460
rect 4300 110404 4356 110460
rect 4356 110404 4360 110460
rect 4296 110400 4360 110404
rect 4376 110460 4440 110464
rect 4376 110404 4380 110460
rect 4380 110404 4436 110460
rect 4436 110404 4440 110460
rect 4376 110400 4440 110404
rect 4456 110460 4520 110464
rect 4456 110404 4460 110460
rect 4460 110404 4516 110460
rect 4516 110404 4520 110460
rect 4456 110400 4520 110404
rect 105924 110460 105988 110464
rect 105924 110404 105928 110460
rect 105928 110404 105984 110460
rect 105984 110404 105988 110460
rect 105924 110400 105988 110404
rect 106004 110460 106068 110464
rect 106004 110404 106008 110460
rect 106008 110404 106064 110460
rect 106064 110404 106068 110460
rect 106004 110400 106068 110404
rect 106084 110460 106148 110464
rect 106084 110404 106088 110460
rect 106088 110404 106144 110460
rect 106144 110404 106148 110460
rect 106084 110400 106148 110404
rect 106164 110460 106228 110464
rect 106164 110404 106168 110460
rect 106168 110404 106224 110460
rect 106224 110404 106228 110460
rect 106164 110400 106228 110404
rect 4876 109916 4940 109920
rect 4876 109860 4880 109916
rect 4880 109860 4936 109916
rect 4936 109860 4940 109916
rect 4876 109856 4940 109860
rect 4956 109916 5020 109920
rect 4956 109860 4960 109916
rect 4960 109860 5016 109916
rect 5016 109860 5020 109916
rect 4956 109856 5020 109860
rect 5036 109916 5100 109920
rect 5036 109860 5040 109916
rect 5040 109860 5096 109916
rect 5096 109860 5100 109916
rect 5036 109856 5100 109860
rect 5116 109916 5180 109920
rect 5116 109860 5120 109916
rect 5120 109860 5176 109916
rect 5176 109860 5180 109916
rect 5116 109856 5180 109860
rect 106660 109916 106724 109920
rect 106660 109860 106664 109916
rect 106664 109860 106720 109916
rect 106720 109860 106724 109916
rect 106660 109856 106724 109860
rect 106740 109916 106804 109920
rect 106740 109860 106744 109916
rect 106744 109860 106800 109916
rect 106800 109860 106804 109916
rect 106740 109856 106804 109860
rect 106820 109916 106884 109920
rect 106820 109860 106824 109916
rect 106824 109860 106880 109916
rect 106880 109860 106884 109916
rect 106820 109856 106884 109860
rect 106900 109916 106964 109920
rect 106900 109860 106904 109916
rect 106904 109860 106960 109916
rect 106960 109860 106964 109916
rect 106900 109856 106964 109860
rect 4216 109372 4280 109376
rect 4216 109316 4220 109372
rect 4220 109316 4276 109372
rect 4276 109316 4280 109372
rect 4216 109312 4280 109316
rect 4296 109372 4360 109376
rect 4296 109316 4300 109372
rect 4300 109316 4356 109372
rect 4356 109316 4360 109372
rect 4296 109312 4360 109316
rect 4376 109372 4440 109376
rect 4376 109316 4380 109372
rect 4380 109316 4436 109372
rect 4436 109316 4440 109372
rect 4376 109312 4440 109316
rect 4456 109372 4520 109376
rect 4456 109316 4460 109372
rect 4460 109316 4516 109372
rect 4516 109316 4520 109372
rect 4456 109312 4520 109316
rect 105924 109372 105988 109376
rect 105924 109316 105928 109372
rect 105928 109316 105984 109372
rect 105984 109316 105988 109372
rect 105924 109312 105988 109316
rect 106004 109372 106068 109376
rect 106004 109316 106008 109372
rect 106008 109316 106064 109372
rect 106064 109316 106068 109372
rect 106004 109312 106068 109316
rect 106084 109372 106148 109376
rect 106084 109316 106088 109372
rect 106088 109316 106144 109372
rect 106144 109316 106148 109372
rect 106084 109312 106148 109316
rect 106164 109372 106228 109376
rect 106164 109316 106168 109372
rect 106168 109316 106224 109372
rect 106224 109316 106228 109372
rect 106164 109312 106228 109316
rect 4876 108828 4940 108832
rect 4876 108772 4880 108828
rect 4880 108772 4936 108828
rect 4936 108772 4940 108828
rect 4876 108768 4940 108772
rect 4956 108828 5020 108832
rect 4956 108772 4960 108828
rect 4960 108772 5016 108828
rect 5016 108772 5020 108828
rect 4956 108768 5020 108772
rect 5036 108828 5100 108832
rect 5036 108772 5040 108828
rect 5040 108772 5096 108828
rect 5096 108772 5100 108828
rect 5036 108768 5100 108772
rect 5116 108828 5180 108832
rect 5116 108772 5120 108828
rect 5120 108772 5176 108828
rect 5176 108772 5180 108828
rect 5116 108768 5180 108772
rect 106660 108828 106724 108832
rect 106660 108772 106664 108828
rect 106664 108772 106720 108828
rect 106720 108772 106724 108828
rect 106660 108768 106724 108772
rect 106740 108828 106804 108832
rect 106740 108772 106744 108828
rect 106744 108772 106800 108828
rect 106800 108772 106804 108828
rect 106740 108768 106804 108772
rect 106820 108828 106884 108832
rect 106820 108772 106824 108828
rect 106824 108772 106880 108828
rect 106880 108772 106884 108828
rect 106820 108768 106884 108772
rect 106900 108828 106964 108832
rect 106900 108772 106904 108828
rect 106904 108772 106960 108828
rect 106960 108772 106964 108828
rect 106900 108768 106964 108772
rect 4216 108284 4280 108288
rect 4216 108228 4220 108284
rect 4220 108228 4276 108284
rect 4276 108228 4280 108284
rect 4216 108224 4280 108228
rect 4296 108284 4360 108288
rect 4296 108228 4300 108284
rect 4300 108228 4356 108284
rect 4356 108228 4360 108284
rect 4296 108224 4360 108228
rect 4376 108284 4440 108288
rect 4376 108228 4380 108284
rect 4380 108228 4436 108284
rect 4436 108228 4440 108284
rect 4376 108224 4440 108228
rect 4456 108284 4520 108288
rect 4456 108228 4460 108284
rect 4460 108228 4516 108284
rect 4516 108228 4520 108284
rect 4456 108224 4520 108228
rect 105924 108284 105988 108288
rect 105924 108228 105928 108284
rect 105928 108228 105984 108284
rect 105984 108228 105988 108284
rect 105924 108224 105988 108228
rect 106004 108284 106068 108288
rect 106004 108228 106008 108284
rect 106008 108228 106064 108284
rect 106064 108228 106068 108284
rect 106004 108224 106068 108228
rect 106084 108284 106148 108288
rect 106084 108228 106088 108284
rect 106088 108228 106144 108284
rect 106144 108228 106148 108284
rect 106084 108224 106148 108228
rect 106164 108284 106228 108288
rect 106164 108228 106168 108284
rect 106168 108228 106224 108284
rect 106224 108228 106228 108284
rect 106164 108224 106228 108228
rect 4876 107740 4940 107744
rect 4876 107684 4880 107740
rect 4880 107684 4936 107740
rect 4936 107684 4940 107740
rect 4876 107680 4940 107684
rect 4956 107740 5020 107744
rect 4956 107684 4960 107740
rect 4960 107684 5016 107740
rect 5016 107684 5020 107740
rect 4956 107680 5020 107684
rect 5036 107740 5100 107744
rect 5036 107684 5040 107740
rect 5040 107684 5096 107740
rect 5096 107684 5100 107740
rect 5036 107680 5100 107684
rect 5116 107740 5180 107744
rect 5116 107684 5120 107740
rect 5120 107684 5176 107740
rect 5176 107684 5180 107740
rect 5116 107680 5180 107684
rect 106660 107740 106724 107744
rect 106660 107684 106664 107740
rect 106664 107684 106720 107740
rect 106720 107684 106724 107740
rect 106660 107680 106724 107684
rect 106740 107740 106804 107744
rect 106740 107684 106744 107740
rect 106744 107684 106800 107740
rect 106800 107684 106804 107740
rect 106740 107680 106804 107684
rect 106820 107740 106884 107744
rect 106820 107684 106824 107740
rect 106824 107684 106880 107740
rect 106880 107684 106884 107740
rect 106820 107680 106884 107684
rect 106900 107740 106964 107744
rect 106900 107684 106904 107740
rect 106904 107684 106960 107740
rect 106960 107684 106964 107740
rect 106900 107680 106964 107684
rect 4216 107196 4280 107200
rect 4216 107140 4220 107196
rect 4220 107140 4276 107196
rect 4276 107140 4280 107196
rect 4216 107136 4280 107140
rect 4296 107196 4360 107200
rect 4296 107140 4300 107196
rect 4300 107140 4356 107196
rect 4356 107140 4360 107196
rect 4296 107136 4360 107140
rect 4376 107196 4440 107200
rect 4376 107140 4380 107196
rect 4380 107140 4436 107196
rect 4436 107140 4440 107196
rect 4376 107136 4440 107140
rect 4456 107196 4520 107200
rect 4456 107140 4460 107196
rect 4460 107140 4516 107196
rect 4516 107140 4520 107196
rect 4456 107136 4520 107140
rect 105924 107196 105988 107200
rect 105924 107140 105928 107196
rect 105928 107140 105984 107196
rect 105984 107140 105988 107196
rect 105924 107136 105988 107140
rect 106004 107196 106068 107200
rect 106004 107140 106008 107196
rect 106008 107140 106064 107196
rect 106064 107140 106068 107196
rect 106004 107136 106068 107140
rect 106084 107196 106148 107200
rect 106084 107140 106088 107196
rect 106088 107140 106144 107196
rect 106144 107140 106148 107196
rect 106084 107136 106148 107140
rect 106164 107196 106228 107200
rect 106164 107140 106168 107196
rect 106168 107140 106224 107196
rect 106224 107140 106228 107196
rect 106164 107136 106228 107140
rect 4876 106652 4940 106656
rect 4876 106596 4880 106652
rect 4880 106596 4936 106652
rect 4936 106596 4940 106652
rect 4876 106592 4940 106596
rect 4956 106652 5020 106656
rect 4956 106596 4960 106652
rect 4960 106596 5016 106652
rect 5016 106596 5020 106652
rect 4956 106592 5020 106596
rect 5036 106652 5100 106656
rect 5036 106596 5040 106652
rect 5040 106596 5096 106652
rect 5096 106596 5100 106652
rect 5036 106592 5100 106596
rect 5116 106652 5180 106656
rect 5116 106596 5120 106652
rect 5120 106596 5176 106652
rect 5176 106596 5180 106652
rect 5116 106592 5180 106596
rect 106660 106652 106724 106656
rect 106660 106596 106664 106652
rect 106664 106596 106720 106652
rect 106720 106596 106724 106652
rect 106660 106592 106724 106596
rect 106740 106652 106804 106656
rect 106740 106596 106744 106652
rect 106744 106596 106800 106652
rect 106800 106596 106804 106652
rect 106740 106592 106804 106596
rect 106820 106652 106884 106656
rect 106820 106596 106824 106652
rect 106824 106596 106880 106652
rect 106880 106596 106884 106652
rect 106820 106592 106884 106596
rect 106900 106652 106964 106656
rect 106900 106596 106904 106652
rect 106904 106596 106960 106652
rect 106960 106596 106964 106652
rect 106900 106592 106964 106596
rect 4216 106108 4280 106112
rect 4216 106052 4220 106108
rect 4220 106052 4276 106108
rect 4276 106052 4280 106108
rect 4216 106048 4280 106052
rect 4296 106108 4360 106112
rect 4296 106052 4300 106108
rect 4300 106052 4356 106108
rect 4356 106052 4360 106108
rect 4296 106048 4360 106052
rect 4376 106108 4440 106112
rect 4376 106052 4380 106108
rect 4380 106052 4436 106108
rect 4436 106052 4440 106108
rect 4376 106048 4440 106052
rect 4456 106108 4520 106112
rect 4456 106052 4460 106108
rect 4460 106052 4516 106108
rect 4516 106052 4520 106108
rect 4456 106048 4520 106052
rect 105924 106108 105988 106112
rect 105924 106052 105928 106108
rect 105928 106052 105984 106108
rect 105984 106052 105988 106108
rect 105924 106048 105988 106052
rect 106004 106108 106068 106112
rect 106004 106052 106008 106108
rect 106008 106052 106064 106108
rect 106064 106052 106068 106108
rect 106004 106048 106068 106052
rect 106084 106108 106148 106112
rect 106084 106052 106088 106108
rect 106088 106052 106144 106108
rect 106144 106052 106148 106108
rect 106084 106048 106148 106052
rect 106164 106108 106228 106112
rect 106164 106052 106168 106108
rect 106168 106052 106224 106108
rect 106224 106052 106228 106108
rect 106164 106048 106228 106052
rect 4876 105564 4940 105568
rect 4876 105508 4880 105564
rect 4880 105508 4936 105564
rect 4936 105508 4940 105564
rect 4876 105504 4940 105508
rect 4956 105564 5020 105568
rect 4956 105508 4960 105564
rect 4960 105508 5016 105564
rect 5016 105508 5020 105564
rect 4956 105504 5020 105508
rect 5036 105564 5100 105568
rect 5036 105508 5040 105564
rect 5040 105508 5096 105564
rect 5096 105508 5100 105564
rect 5036 105504 5100 105508
rect 5116 105564 5180 105568
rect 5116 105508 5120 105564
rect 5120 105508 5176 105564
rect 5176 105508 5180 105564
rect 5116 105504 5180 105508
rect 106660 105564 106724 105568
rect 106660 105508 106664 105564
rect 106664 105508 106720 105564
rect 106720 105508 106724 105564
rect 106660 105504 106724 105508
rect 106740 105564 106804 105568
rect 106740 105508 106744 105564
rect 106744 105508 106800 105564
rect 106800 105508 106804 105564
rect 106740 105504 106804 105508
rect 106820 105564 106884 105568
rect 106820 105508 106824 105564
rect 106824 105508 106880 105564
rect 106880 105508 106884 105564
rect 106820 105504 106884 105508
rect 106900 105564 106964 105568
rect 106900 105508 106904 105564
rect 106904 105508 106960 105564
rect 106960 105508 106964 105564
rect 106900 105504 106964 105508
rect 4216 105020 4280 105024
rect 4216 104964 4220 105020
rect 4220 104964 4276 105020
rect 4276 104964 4280 105020
rect 4216 104960 4280 104964
rect 4296 105020 4360 105024
rect 4296 104964 4300 105020
rect 4300 104964 4356 105020
rect 4356 104964 4360 105020
rect 4296 104960 4360 104964
rect 4376 105020 4440 105024
rect 4376 104964 4380 105020
rect 4380 104964 4436 105020
rect 4436 104964 4440 105020
rect 4376 104960 4440 104964
rect 4456 105020 4520 105024
rect 4456 104964 4460 105020
rect 4460 104964 4516 105020
rect 4516 104964 4520 105020
rect 4456 104960 4520 104964
rect 105924 105020 105988 105024
rect 105924 104964 105928 105020
rect 105928 104964 105984 105020
rect 105984 104964 105988 105020
rect 105924 104960 105988 104964
rect 106004 105020 106068 105024
rect 106004 104964 106008 105020
rect 106008 104964 106064 105020
rect 106064 104964 106068 105020
rect 106004 104960 106068 104964
rect 106084 105020 106148 105024
rect 106084 104964 106088 105020
rect 106088 104964 106144 105020
rect 106144 104964 106148 105020
rect 106084 104960 106148 104964
rect 106164 105020 106228 105024
rect 106164 104964 106168 105020
rect 106168 104964 106224 105020
rect 106224 104964 106228 105020
rect 106164 104960 106228 104964
rect 4876 104476 4940 104480
rect 4876 104420 4880 104476
rect 4880 104420 4936 104476
rect 4936 104420 4940 104476
rect 4876 104416 4940 104420
rect 4956 104476 5020 104480
rect 4956 104420 4960 104476
rect 4960 104420 5016 104476
rect 5016 104420 5020 104476
rect 4956 104416 5020 104420
rect 5036 104476 5100 104480
rect 5036 104420 5040 104476
rect 5040 104420 5096 104476
rect 5096 104420 5100 104476
rect 5036 104416 5100 104420
rect 5116 104476 5180 104480
rect 5116 104420 5120 104476
rect 5120 104420 5176 104476
rect 5176 104420 5180 104476
rect 5116 104416 5180 104420
rect 106660 104476 106724 104480
rect 106660 104420 106664 104476
rect 106664 104420 106720 104476
rect 106720 104420 106724 104476
rect 106660 104416 106724 104420
rect 106740 104476 106804 104480
rect 106740 104420 106744 104476
rect 106744 104420 106800 104476
rect 106800 104420 106804 104476
rect 106740 104416 106804 104420
rect 106820 104476 106884 104480
rect 106820 104420 106824 104476
rect 106824 104420 106880 104476
rect 106880 104420 106884 104476
rect 106820 104416 106884 104420
rect 106900 104476 106964 104480
rect 106900 104420 106904 104476
rect 106904 104420 106960 104476
rect 106960 104420 106964 104476
rect 106900 104416 106964 104420
rect 4216 103932 4280 103936
rect 4216 103876 4220 103932
rect 4220 103876 4276 103932
rect 4276 103876 4280 103932
rect 4216 103872 4280 103876
rect 4296 103932 4360 103936
rect 4296 103876 4300 103932
rect 4300 103876 4356 103932
rect 4356 103876 4360 103932
rect 4296 103872 4360 103876
rect 4376 103932 4440 103936
rect 4376 103876 4380 103932
rect 4380 103876 4436 103932
rect 4436 103876 4440 103932
rect 4376 103872 4440 103876
rect 4456 103932 4520 103936
rect 4456 103876 4460 103932
rect 4460 103876 4516 103932
rect 4516 103876 4520 103932
rect 4456 103872 4520 103876
rect 105924 103932 105988 103936
rect 105924 103876 105928 103932
rect 105928 103876 105984 103932
rect 105984 103876 105988 103932
rect 105924 103872 105988 103876
rect 106004 103932 106068 103936
rect 106004 103876 106008 103932
rect 106008 103876 106064 103932
rect 106064 103876 106068 103932
rect 106004 103872 106068 103876
rect 106084 103932 106148 103936
rect 106084 103876 106088 103932
rect 106088 103876 106144 103932
rect 106144 103876 106148 103932
rect 106084 103872 106148 103876
rect 106164 103932 106228 103936
rect 106164 103876 106168 103932
rect 106168 103876 106224 103932
rect 106224 103876 106228 103932
rect 106164 103872 106228 103876
rect 4876 103388 4940 103392
rect 4876 103332 4880 103388
rect 4880 103332 4936 103388
rect 4936 103332 4940 103388
rect 4876 103328 4940 103332
rect 4956 103388 5020 103392
rect 4956 103332 4960 103388
rect 4960 103332 5016 103388
rect 5016 103332 5020 103388
rect 4956 103328 5020 103332
rect 5036 103388 5100 103392
rect 5036 103332 5040 103388
rect 5040 103332 5096 103388
rect 5096 103332 5100 103388
rect 5036 103328 5100 103332
rect 5116 103388 5180 103392
rect 5116 103332 5120 103388
rect 5120 103332 5176 103388
rect 5176 103332 5180 103388
rect 5116 103328 5180 103332
rect 106660 103388 106724 103392
rect 106660 103332 106664 103388
rect 106664 103332 106720 103388
rect 106720 103332 106724 103388
rect 106660 103328 106724 103332
rect 106740 103388 106804 103392
rect 106740 103332 106744 103388
rect 106744 103332 106800 103388
rect 106800 103332 106804 103388
rect 106740 103328 106804 103332
rect 106820 103388 106884 103392
rect 106820 103332 106824 103388
rect 106824 103332 106880 103388
rect 106880 103332 106884 103388
rect 106820 103328 106884 103332
rect 106900 103388 106964 103392
rect 106900 103332 106904 103388
rect 106904 103332 106960 103388
rect 106960 103332 106964 103388
rect 106900 103328 106964 103332
rect 4216 102844 4280 102848
rect 4216 102788 4220 102844
rect 4220 102788 4276 102844
rect 4276 102788 4280 102844
rect 4216 102784 4280 102788
rect 4296 102844 4360 102848
rect 4296 102788 4300 102844
rect 4300 102788 4356 102844
rect 4356 102788 4360 102844
rect 4296 102784 4360 102788
rect 4376 102844 4440 102848
rect 4376 102788 4380 102844
rect 4380 102788 4436 102844
rect 4436 102788 4440 102844
rect 4376 102784 4440 102788
rect 4456 102844 4520 102848
rect 4456 102788 4460 102844
rect 4460 102788 4516 102844
rect 4516 102788 4520 102844
rect 4456 102784 4520 102788
rect 105924 102844 105988 102848
rect 105924 102788 105928 102844
rect 105928 102788 105984 102844
rect 105984 102788 105988 102844
rect 105924 102784 105988 102788
rect 106004 102844 106068 102848
rect 106004 102788 106008 102844
rect 106008 102788 106064 102844
rect 106064 102788 106068 102844
rect 106004 102784 106068 102788
rect 106084 102844 106148 102848
rect 106084 102788 106088 102844
rect 106088 102788 106144 102844
rect 106144 102788 106148 102844
rect 106084 102784 106148 102788
rect 106164 102844 106228 102848
rect 106164 102788 106168 102844
rect 106168 102788 106224 102844
rect 106224 102788 106228 102844
rect 106164 102784 106228 102788
rect 4876 102300 4940 102304
rect 4876 102244 4880 102300
rect 4880 102244 4936 102300
rect 4936 102244 4940 102300
rect 4876 102240 4940 102244
rect 4956 102300 5020 102304
rect 4956 102244 4960 102300
rect 4960 102244 5016 102300
rect 5016 102244 5020 102300
rect 4956 102240 5020 102244
rect 5036 102300 5100 102304
rect 5036 102244 5040 102300
rect 5040 102244 5096 102300
rect 5096 102244 5100 102300
rect 5036 102240 5100 102244
rect 5116 102300 5180 102304
rect 5116 102244 5120 102300
rect 5120 102244 5176 102300
rect 5176 102244 5180 102300
rect 5116 102240 5180 102244
rect 106660 102300 106724 102304
rect 106660 102244 106664 102300
rect 106664 102244 106720 102300
rect 106720 102244 106724 102300
rect 106660 102240 106724 102244
rect 106740 102300 106804 102304
rect 106740 102244 106744 102300
rect 106744 102244 106800 102300
rect 106800 102244 106804 102300
rect 106740 102240 106804 102244
rect 106820 102300 106884 102304
rect 106820 102244 106824 102300
rect 106824 102244 106880 102300
rect 106880 102244 106884 102300
rect 106820 102240 106884 102244
rect 106900 102300 106964 102304
rect 106900 102244 106904 102300
rect 106904 102244 106960 102300
rect 106960 102244 106964 102300
rect 106900 102240 106964 102244
rect 4216 101756 4280 101760
rect 4216 101700 4220 101756
rect 4220 101700 4276 101756
rect 4276 101700 4280 101756
rect 4216 101696 4280 101700
rect 4296 101756 4360 101760
rect 4296 101700 4300 101756
rect 4300 101700 4356 101756
rect 4356 101700 4360 101756
rect 4296 101696 4360 101700
rect 4376 101756 4440 101760
rect 4376 101700 4380 101756
rect 4380 101700 4436 101756
rect 4436 101700 4440 101756
rect 4376 101696 4440 101700
rect 4456 101756 4520 101760
rect 4456 101700 4460 101756
rect 4460 101700 4516 101756
rect 4516 101700 4520 101756
rect 4456 101696 4520 101700
rect 105924 101756 105988 101760
rect 105924 101700 105928 101756
rect 105928 101700 105984 101756
rect 105984 101700 105988 101756
rect 105924 101696 105988 101700
rect 106004 101756 106068 101760
rect 106004 101700 106008 101756
rect 106008 101700 106064 101756
rect 106064 101700 106068 101756
rect 106004 101696 106068 101700
rect 106084 101756 106148 101760
rect 106084 101700 106088 101756
rect 106088 101700 106144 101756
rect 106144 101700 106148 101756
rect 106084 101696 106148 101700
rect 106164 101756 106228 101760
rect 106164 101700 106168 101756
rect 106168 101700 106224 101756
rect 106224 101700 106228 101756
rect 106164 101696 106228 101700
rect 4876 101212 4940 101216
rect 4876 101156 4880 101212
rect 4880 101156 4936 101212
rect 4936 101156 4940 101212
rect 4876 101152 4940 101156
rect 4956 101212 5020 101216
rect 4956 101156 4960 101212
rect 4960 101156 5016 101212
rect 5016 101156 5020 101212
rect 4956 101152 5020 101156
rect 5036 101212 5100 101216
rect 5036 101156 5040 101212
rect 5040 101156 5096 101212
rect 5096 101156 5100 101212
rect 5036 101152 5100 101156
rect 5116 101212 5180 101216
rect 5116 101156 5120 101212
rect 5120 101156 5176 101212
rect 5176 101156 5180 101212
rect 5116 101152 5180 101156
rect 106660 101212 106724 101216
rect 106660 101156 106664 101212
rect 106664 101156 106720 101212
rect 106720 101156 106724 101212
rect 106660 101152 106724 101156
rect 106740 101212 106804 101216
rect 106740 101156 106744 101212
rect 106744 101156 106800 101212
rect 106800 101156 106804 101212
rect 106740 101152 106804 101156
rect 106820 101212 106884 101216
rect 106820 101156 106824 101212
rect 106824 101156 106880 101212
rect 106880 101156 106884 101212
rect 106820 101152 106884 101156
rect 106900 101212 106964 101216
rect 106900 101156 106904 101212
rect 106904 101156 106960 101212
rect 106960 101156 106964 101212
rect 106900 101152 106964 101156
rect 4216 100668 4280 100672
rect 4216 100612 4220 100668
rect 4220 100612 4276 100668
rect 4276 100612 4280 100668
rect 4216 100608 4280 100612
rect 4296 100668 4360 100672
rect 4296 100612 4300 100668
rect 4300 100612 4356 100668
rect 4356 100612 4360 100668
rect 4296 100608 4360 100612
rect 4376 100668 4440 100672
rect 4376 100612 4380 100668
rect 4380 100612 4436 100668
rect 4436 100612 4440 100668
rect 4376 100608 4440 100612
rect 4456 100668 4520 100672
rect 4456 100612 4460 100668
rect 4460 100612 4516 100668
rect 4516 100612 4520 100668
rect 4456 100608 4520 100612
rect 105924 100668 105988 100672
rect 105924 100612 105928 100668
rect 105928 100612 105984 100668
rect 105984 100612 105988 100668
rect 105924 100608 105988 100612
rect 106004 100668 106068 100672
rect 106004 100612 106008 100668
rect 106008 100612 106064 100668
rect 106064 100612 106068 100668
rect 106004 100608 106068 100612
rect 106084 100668 106148 100672
rect 106084 100612 106088 100668
rect 106088 100612 106144 100668
rect 106144 100612 106148 100668
rect 106084 100608 106148 100612
rect 106164 100668 106228 100672
rect 106164 100612 106168 100668
rect 106168 100612 106224 100668
rect 106224 100612 106228 100668
rect 106164 100608 106228 100612
rect 4876 100124 4940 100128
rect 4876 100068 4880 100124
rect 4880 100068 4936 100124
rect 4936 100068 4940 100124
rect 4876 100064 4940 100068
rect 4956 100124 5020 100128
rect 4956 100068 4960 100124
rect 4960 100068 5016 100124
rect 5016 100068 5020 100124
rect 4956 100064 5020 100068
rect 5036 100124 5100 100128
rect 5036 100068 5040 100124
rect 5040 100068 5096 100124
rect 5096 100068 5100 100124
rect 5036 100064 5100 100068
rect 5116 100124 5180 100128
rect 5116 100068 5120 100124
rect 5120 100068 5176 100124
rect 5176 100068 5180 100124
rect 5116 100064 5180 100068
rect 106660 100124 106724 100128
rect 106660 100068 106664 100124
rect 106664 100068 106720 100124
rect 106720 100068 106724 100124
rect 106660 100064 106724 100068
rect 106740 100124 106804 100128
rect 106740 100068 106744 100124
rect 106744 100068 106800 100124
rect 106800 100068 106804 100124
rect 106740 100064 106804 100068
rect 106820 100124 106884 100128
rect 106820 100068 106824 100124
rect 106824 100068 106880 100124
rect 106880 100068 106884 100124
rect 106820 100064 106884 100068
rect 106900 100124 106964 100128
rect 106900 100068 106904 100124
rect 106904 100068 106960 100124
rect 106960 100068 106964 100124
rect 106900 100064 106964 100068
rect 4216 99580 4280 99584
rect 4216 99524 4220 99580
rect 4220 99524 4276 99580
rect 4276 99524 4280 99580
rect 4216 99520 4280 99524
rect 4296 99580 4360 99584
rect 4296 99524 4300 99580
rect 4300 99524 4356 99580
rect 4356 99524 4360 99580
rect 4296 99520 4360 99524
rect 4376 99580 4440 99584
rect 4376 99524 4380 99580
rect 4380 99524 4436 99580
rect 4436 99524 4440 99580
rect 4376 99520 4440 99524
rect 4456 99580 4520 99584
rect 4456 99524 4460 99580
rect 4460 99524 4516 99580
rect 4516 99524 4520 99580
rect 4456 99520 4520 99524
rect 105924 99580 105988 99584
rect 105924 99524 105928 99580
rect 105928 99524 105984 99580
rect 105984 99524 105988 99580
rect 105924 99520 105988 99524
rect 106004 99580 106068 99584
rect 106004 99524 106008 99580
rect 106008 99524 106064 99580
rect 106064 99524 106068 99580
rect 106004 99520 106068 99524
rect 106084 99580 106148 99584
rect 106084 99524 106088 99580
rect 106088 99524 106144 99580
rect 106144 99524 106148 99580
rect 106084 99520 106148 99524
rect 106164 99580 106228 99584
rect 106164 99524 106168 99580
rect 106168 99524 106224 99580
rect 106224 99524 106228 99580
rect 106164 99520 106228 99524
rect 4876 99036 4940 99040
rect 4876 98980 4880 99036
rect 4880 98980 4936 99036
rect 4936 98980 4940 99036
rect 4876 98976 4940 98980
rect 4956 99036 5020 99040
rect 4956 98980 4960 99036
rect 4960 98980 5016 99036
rect 5016 98980 5020 99036
rect 4956 98976 5020 98980
rect 5036 99036 5100 99040
rect 5036 98980 5040 99036
rect 5040 98980 5096 99036
rect 5096 98980 5100 99036
rect 5036 98976 5100 98980
rect 5116 99036 5180 99040
rect 5116 98980 5120 99036
rect 5120 98980 5176 99036
rect 5176 98980 5180 99036
rect 5116 98976 5180 98980
rect 106660 99036 106724 99040
rect 106660 98980 106664 99036
rect 106664 98980 106720 99036
rect 106720 98980 106724 99036
rect 106660 98976 106724 98980
rect 106740 99036 106804 99040
rect 106740 98980 106744 99036
rect 106744 98980 106800 99036
rect 106800 98980 106804 99036
rect 106740 98976 106804 98980
rect 106820 99036 106884 99040
rect 106820 98980 106824 99036
rect 106824 98980 106880 99036
rect 106880 98980 106884 99036
rect 106820 98976 106884 98980
rect 106900 99036 106964 99040
rect 106900 98980 106904 99036
rect 106904 98980 106960 99036
rect 106960 98980 106964 99036
rect 106900 98976 106964 98980
rect 4216 98492 4280 98496
rect 4216 98436 4220 98492
rect 4220 98436 4276 98492
rect 4276 98436 4280 98492
rect 4216 98432 4280 98436
rect 4296 98492 4360 98496
rect 4296 98436 4300 98492
rect 4300 98436 4356 98492
rect 4356 98436 4360 98492
rect 4296 98432 4360 98436
rect 4376 98492 4440 98496
rect 4376 98436 4380 98492
rect 4380 98436 4436 98492
rect 4436 98436 4440 98492
rect 4376 98432 4440 98436
rect 4456 98492 4520 98496
rect 4456 98436 4460 98492
rect 4460 98436 4516 98492
rect 4516 98436 4520 98492
rect 4456 98432 4520 98436
rect 105924 98492 105988 98496
rect 105924 98436 105928 98492
rect 105928 98436 105984 98492
rect 105984 98436 105988 98492
rect 105924 98432 105988 98436
rect 106004 98492 106068 98496
rect 106004 98436 106008 98492
rect 106008 98436 106064 98492
rect 106064 98436 106068 98492
rect 106004 98432 106068 98436
rect 106084 98492 106148 98496
rect 106084 98436 106088 98492
rect 106088 98436 106144 98492
rect 106144 98436 106148 98492
rect 106084 98432 106148 98436
rect 106164 98492 106228 98496
rect 106164 98436 106168 98492
rect 106168 98436 106224 98492
rect 106224 98436 106228 98492
rect 106164 98432 106228 98436
rect 4876 97948 4940 97952
rect 4876 97892 4880 97948
rect 4880 97892 4936 97948
rect 4936 97892 4940 97948
rect 4876 97888 4940 97892
rect 4956 97948 5020 97952
rect 4956 97892 4960 97948
rect 4960 97892 5016 97948
rect 5016 97892 5020 97948
rect 4956 97888 5020 97892
rect 5036 97948 5100 97952
rect 5036 97892 5040 97948
rect 5040 97892 5096 97948
rect 5096 97892 5100 97948
rect 5036 97888 5100 97892
rect 5116 97948 5180 97952
rect 5116 97892 5120 97948
rect 5120 97892 5176 97948
rect 5176 97892 5180 97948
rect 5116 97888 5180 97892
rect 106660 97948 106724 97952
rect 106660 97892 106664 97948
rect 106664 97892 106720 97948
rect 106720 97892 106724 97948
rect 106660 97888 106724 97892
rect 106740 97948 106804 97952
rect 106740 97892 106744 97948
rect 106744 97892 106800 97948
rect 106800 97892 106804 97948
rect 106740 97888 106804 97892
rect 106820 97948 106884 97952
rect 106820 97892 106824 97948
rect 106824 97892 106880 97948
rect 106880 97892 106884 97948
rect 106820 97888 106884 97892
rect 106900 97948 106964 97952
rect 106900 97892 106904 97948
rect 106904 97892 106960 97948
rect 106960 97892 106964 97948
rect 106900 97888 106964 97892
rect 4216 97404 4280 97408
rect 4216 97348 4220 97404
rect 4220 97348 4276 97404
rect 4276 97348 4280 97404
rect 4216 97344 4280 97348
rect 4296 97404 4360 97408
rect 4296 97348 4300 97404
rect 4300 97348 4356 97404
rect 4356 97348 4360 97404
rect 4296 97344 4360 97348
rect 4376 97404 4440 97408
rect 4376 97348 4380 97404
rect 4380 97348 4436 97404
rect 4436 97348 4440 97404
rect 4376 97344 4440 97348
rect 4456 97404 4520 97408
rect 4456 97348 4460 97404
rect 4460 97348 4516 97404
rect 4516 97348 4520 97404
rect 4456 97344 4520 97348
rect 105924 97404 105988 97408
rect 105924 97348 105928 97404
rect 105928 97348 105984 97404
rect 105984 97348 105988 97404
rect 105924 97344 105988 97348
rect 106004 97404 106068 97408
rect 106004 97348 106008 97404
rect 106008 97348 106064 97404
rect 106064 97348 106068 97404
rect 106004 97344 106068 97348
rect 106084 97404 106148 97408
rect 106084 97348 106088 97404
rect 106088 97348 106144 97404
rect 106144 97348 106148 97404
rect 106084 97344 106148 97348
rect 106164 97404 106228 97408
rect 106164 97348 106168 97404
rect 106168 97348 106224 97404
rect 106224 97348 106228 97404
rect 106164 97344 106228 97348
rect 4876 96860 4940 96864
rect 4876 96804 4880 96860
rect 4880 96804 4936 96860
rect 4936 96804 4940 96860
rect 4876 96800 4940 96804
rect 4956 96860 5020 96864
rect 4956 96804 4960 96860
rect 4960 96804 5016 96860
rect 5016 96804 5020 96860
rect 4956 96800 5020 96804
rect 5036 96860 5100 96864
rect 5036 96804 5040 96860
rect 5040 96804 5096 96860
rect 5096 96804 5100 96860
rect 5036 96800 5100 96804
rect 5116 96860 5180 96864
rect 5116 96804 5120 96860
rect 5120 96804 5176 96860
rect 5176 96804 5180 96860
rect 5116 96800 5180 96804
rect 106660 96860 106724 96864
rect 106660 96804 106664 96860
rect 106664 96804 106720 96860
rect 106720 96804 106724 96860
rect 106660 96800 106724 96804
rect 106740 96860 106804 96864
rect 106740 96804 106744 96860
rect 106744 96804 106800 96860
rect 106800 96804 106804 96860
rect 106740 96800 106804 96804
rect 106820 96860 106884 96864
rect 106820 96804 106824 96860
rect 106824 96804 106880 96860
rect 106880 96804 106884 96860
rect 106820 96800 106884 96804
rect 106900 96860 106964 96864
rect 106900 96804 106904 96860
rect 106904 96804 106960 96860
rect 106960 96804 106964 96860
rect 106900 96800 106964 96804
rect 4216 96316 4280 96320
rect 4216 96260 4220 96316
rect 4220 96260 4276 96316
rect 4276 96260 4280 96316
rect 4216 96256 4280 96260
rect 4296 96316 4360 96320
rect 4296 96260 4300 96316
rect 4300 96260 4356 96316
rect 4356 96260 4360 96316
rect 4296 96256 4360 96260
rect 4376 96316 4440 96320
rect 4376 96260 4380 96316
rect 4380 96260 4436 96316
rect 4436 96260 4440 96316
rect 4376 96256 4440 96260
rect 4456 96316 4520 96320
rect 4456 96260 4460 96316
rect 4460 96260 4516 96316
rect 4516 96260 4520 96316
rect 4456 96256 4520 96260
rect 105924 96316 105988 96320
rect 105924 96260 105928 96316
rect 105928 96260 105984 96316
rect 105984 96260 105988 96316
rect 105924 96256 105988 96260
rect 106004 96316 106068 96320
rect 106004 96260 106008 96316
rect 106008 96260 106064 96316
rect 106064 96260 106068 96316
rect 106004 96256 106068 96260
rect 106084 96316 106148 96320
rect 106084 96260 106088 96316
rect 106088 96260 106144 96316
rect 106144 96260 106148 96316
rect 106084 96256 106148 96260
rect 106164 96316 106228 96320
rect 106164 96260 106168 96316
rect 106168 96260 106224 96316
rect 106224 96260 106228 96316
rect 106164 96256 106228 96260
rect 4876 95772 4940 95776
rect 4876 95716 4880 95772
rect 4880 95716 4936 95772
rect 4936 95716 4940 95772
rect 4876 95712 4940 95716
rect 4956 95772 5020 95776
rect 4956 95716 4960 95772
rect 4960 95716 5016 95772
rect 5016 95716 5020 95772
rect 4956 95712 5020 95716
rect 5036 95772 5100 95776
rect 5036 95716 5040 95772
rect 5040 95716 5096 95772
rect 5096 95716 5100 95772
rect 5036 95712 5100 95716
rect 5116 95772 5180 95776
rect 5116 95716 5120 95772
rect 5120 95716 5176 95772
rect 5176 95716 5180 95772
rect 5116 95712 5180 95716
rect 106660 95772 106724 95776
rect 106660 95716 106664 95772
rect 106664 95716 106720 95772
rect 106720 95716 106724 95772
rect 106660 95712 106724 95716
rect 106740 95772 106804 95776
rect 106740 95716 106744 95772
rect 106744 95716 106800 95772
rect 106800 95716 106804 95772
rect 106740 95712 106804 95716
rect 106820 95772 106884 95776
rect 106820 95716 106824 95772
rect 106824 95716 106880 95772
rect 106880 95716 106884 95772
rect 106820 95712 106884 95716
rect 106900 95772 106964 95776
rect 106900 95716 106904 95772
rect 106904 95716 106960 95772
rect 106960 95716 106964 95772
rect 106900 95712 106964 95716
rect 4216 95228 4280 95232
rect 4216 95172 4220 95228
rect 4220 95172 4276 95228
rect 4276 95172 4280 95228
rect 4216 95168 4280 95172
rect 4296 95228 4360 95232
rect 4296 95172 4300 95228
rect 4300 95172 4356 95228
rect 4356 95172 4360 95228
rect 4296 95168 4360 95172
rect 4376 95228 4440 95232
rect 4376 95172 4380 95228
rect 4380 95172 4436 95228
rect 4436 95172 4440 95228
rect 4376 95168 4440 95172
rect 4456 95228 4520 95232
rect 4456 95172 4460 95228
rect 4460 95172 4516 95228
rect 4516 95172 4520 95228
rect 4456 95168 4520 95172
rect 105924 95228 105988 95232
rect 105924 95172 105928 95228
rect 105928 95172 105984 95228
rect 105984 95172 105988 95228
rect 105924 95168 105988 95172
rect 106004 95228 106068 95232
rect 106004 95172 106008 95228
rect 106008 95172 106064 95228
rect 106064 95172 106068 95228
rect 106004 95168 106068 95172
rect 106084 95228 106148 95232
rect 106084 95172 106088 95228
rect 106088 95172 106144 95228
rect 106144 95172 106148 95228
rect 106084 95168 106148 95172
rect 106164 95228 106228 95232
rect 106164 95172 106168 95228
rect 106168 95172 106224 95228
rect 106224 95172 106228 95228
rect 106164 95168 106228 95172
rect 4876 94684 4940 94688
rect 4876 94628 4880 94684
rect 4880 94628 4936 94684
rect 4936 94628 4940 94684
rect 4876 94624 4940 94628
rect 4956 94684 5020 94688
rect 4956 94628 4960 94684
rect 4960 94628 5016 94684
rect 5016 94628 5020 94684
rect 4956 94624 5020 94628
rect 5036 94684 5100 94688
rect 5036 94628 5040 94684
rect 5040 94628 5096 94684
rect 5096 94628 5100 94684
rect 5036 94624 5100 94628
rect 5116 94684 5180 94688
rect 5116 94628 5120 94684
rect 5120 94628 5176 94684
rect 5176 94628 5180 94684
rect 5116 94624 5180 94628
rect 106660 94684 106724 94688
rect 106660 94628 106664 94684
rect 106664 94628 106720 94684
rect 106720 94628 106724 94684
rect 106660 94624 106724 94628
rect 106740 94684 106804 94688
rect 106740 94628 106744 94684
rect 106744 94628 106800 94684
rect 106800 94628 106804 94684
rect 106740 94624 106804 94628
rect 106820 94684 106884 94688
rect 106820 94628 106824 94684
rect 106824 94628 106880 94684
rect 106880 94628 106884 94684
rect 106820 94624 106884 94628
rect 106900 94684 106964 94688
rect 106900 94628 106904 94684
rect 106904 94628 106960 94684
rect 106960 94628 106964 94684
rect 106900 94624 106964 94628
rect 4216 94140 4280 94144
rect 4216 94084 4220 94140
rect 4220 94084 4276 94140
rect 4276 94084 4280 94140
rect 4216 94080 4280 94084
rect 4296 94140 4360 94144
rect 4296 94084 4300 94140
rect 4300 94084 4356 94140
rect 4356 94084 4360 94140
rect 4296 94080 4360 94084
rect 4376 94140 4440 94144
rect 4376 94084 4380 94140
rect 4380 94084 4436 94140
rect 4436 94084 4440 94140
rect 4376 94080 4440 94084
rect 4456 94140 4520 94144
rect 4456 94084 4460 94140
rect 4460 94084 4516 94140
rect 4516 94084 4520 94140
rect 4456 94080 4520 94084
rect 105924 94140 105988 94144
rect 105924 94084 105928 94140
rect 105928 94084 105984 94140
rect 105984 94084 105988 94140
rect 105924 94080 105988 94084
rect 106004 94140 106068 94144
rect 106004 94084 106008 94140
rect 106008 94084 106064 94140
rect 106064 94084 106068 94140
rect 106004 94080 106068 94084
rect 106084 94140 106148 94144
rect 106084 94084 106088 94140
rect 106088 94084 106144 94140
rect 106144 94084 106148 94140
rect 106084 94080 106148 94084
rect 106164 94140 106228 94144
rect 106164 94084 106168 94140
rect 106168 94084 106224 94140
rect 106224 94084 106228 94140
rect 106164 94080 106228 94084
rect 4876 93596 4940 93600
rect 4876 93540 4880 93596
rect 4880 93540 4936 93596
rect 4936 93540 4940 93596
rect 4876 93536 4940 93540
rect 4956 93596 5020 93600
rect 4956 93540 4960 93596
rect 4960 93540 5016 93596
rect 5016 93540 5020 93596
rect 4956 93536 5020 93540
rect 5036 93596 5100 93600
rect 5036 93540 5040 93596
rect 5040 93540 5096 93596
rect 5096 93540 5100 93596
rect 5036 93536 5100 93540
rect 5116 93596 5180 93600
rect 5116 93540 5120 93596
rect 5120 93540 5176 93596
rect 5176 93540 5180 93596
rect 5116 93536 5180 93540
rect 106660 93596 106724 93600
rect 106660 93540 106664 93596
rect 106664 93540 106720 93596
rect 106720 93540 106724 93596
rect 106660 93536 106724 93540
rect 106740 93596 106804 93600
rect 106740 93540 106744 93596
rect 106744 93540 106800 93596
rect 106800 93540 106804 93596
rect 106740 93536 106804 93540
rect 106820 93596 106884 93600
rect 106820 93540 106824 93596
rect 106824 93540 106880 93596
rect 106880 93540 106884 93596
rect 106820 93536 106884 93540
rect 106900 93596 106964 93600
rect 106900 93540 106904 93596
rect 106904 93540 106960 93596
rect 106960 93540 106964 93596
rect 106900 93536 106964 93540
rect 4216 93052 4280 93056
rect 4216 92996 4220 93052
rect 4220 92996 4276 93052
rect 4276 92996 4280 93052
rect 4216 92992 4280 92996
rect 4296 93052 4360 93056
rect 4296 92996 4300 93052
rect 4300 92996 4356 93052
rect 4356 92996 4360 93052
rect 4296 92992 4360 92996
rect 4376 93052 4440 93056
rect 4376 92996 4380 93052
rect 4380 92996 4436 93052
rect 4436 92996 4440 93052
rect 4376 92992 4440 92996
rect 4456 93052 4520 93056
rect 4456 92996 4460 93052
rect 4460 92996 4516 93052
rect 4516 92996 4520 93052
rect 4456 92992 4520 92996
rect 105924 93052 105988 93056
rect 105924 92996 105928 93052
rect 105928 92996 105984 93052
rect 105984 92996 105988 93052
rect 105924 92992 105988 92996
rect 106004 93052 106068 93056
rect 106004 92996 106008 93052
rect 106008 92996 106064 93052
rect 106064 92996 106068 93052
rect 106004 92992 106068 92996
rect 106084 93052 106148 93056
rect 106084 92996 106088 93052
rect 106088 92996 106144 93052
rect 106144 92996 106148 93052
rect 106084 92992 106148 92996
rect 106164 93052 106228 93056
rect 106164 92996 106168 93052
rect 106168 92996 106224 93052
rect 106224 92996 106228 93052
rect 106164 92992 106228 92996
rect 4876 92508 4940 92512
rect 4876 92452 4880 92508
rect 4880 92452 4936 92508
rect 4936 92452 4940 92508
rect 4876 92448 4940 92452
rect 4956 92508 5020 92512
rect 4956 92452 4960 92508
rect 4960 92452 5016 92508
rect 5016 92452 5020 92508
rect 4956 92448 5020 92452
rect 5036 92508 5100 92512
rect 5036 92452 5040 92508
rect 5040 92452 5096 92508
rect 5096 92452 5100 92508
rect 5036 92448 5100 92452
rect 5116 92508 5180 92512
rect 5116 92452 5120 92508
rect 5120 92452 5176 92508
rect 5176 92452 5180 92508
rect 5116 92448 5180 92452
rect 106660 92508 106724 92512
rect 106660 92452 106664 92508
rect 106664 92452 106720 92508
rect 106720 92452 106724 92508
rect 106660 92448 106724 92452
rect 106740 92508 106804 92512
rect 106740 92452 106744 92508
rect 106744 92452 106800 92508
rect 106800 92452 106804 92508
rect 106740 92448 106804 92452
rect 106820 92508 106884 92512
rect 106820 92452 106824 92508
rect 106824 92452 106880 92508
rect 106880 92452 106884 92508
rect 106820 92448 106884 92452
rect 106900 92508 106964 92512
rect 106900 92452 106904 92508
rect 106904 92452 106960 92508
rect 106960 92452 106964 92508
rect 106900 92448 106964 92452
rect 4216 91964 4280 91968
rect 4216 91908 4220 91964
rect 4220 91908 4276 91964
rect 4276 91908 4280 91964
rect 4216 91904 4280 91908
rect 4296 91964 4360 91968
rect 4296 91908 4300 91964
rect 4300 91908 4356 91964
rect 4356 91908 4360 91964
rect 4296 91904 4360 91908
rect 4376 91964 4440 91968
rect 4376 91908 4380 91964
rect 4380 91908 4436 91964
rect 4436 91908 4440 91964
rect 4376 91904 4440 91908
rect 4456 91964 4520 91968
rect 4456 91908 4460 91964
rect 4460 91908 4516 91964
rect 4516 91908 4520 91964
rect 4456 91904 4520 91908
rect 105924 91964 105988 91968
rect 105924 91908 105928 91964
rect 105928 91908 105984 91964
rect 105984 91908 105988 91964
rect 105924 91904 105988 91908
rect 106004 91964 106068 91968
rect 106004 91908 106008 91964
rect 106008 91908 106064 91964
rect 106064 91908 106068 91964
rect 106004 91904 106068 91908
rect 106084 91964 106148 91968
rect 106084 91908 106088 91964
rect 106088 91908 106144 91964
rect 106144 91908 106148 91964
rect 106084 91904 106148 91908
rect 106164 91964 106228 91968
rect 106164 91908 106168 91964
rect 106168 91908 106224 91964
rect 106224 91908 106228 91964
rect 106164 91904 106228 91908
rect 4876 91420 4940 91424
rect 4876 91364 4880 91420
rect 4880 91364 4936 91420
rect 4936 91364 4940 91420
rect 4876 91360 4940 91364
rect 4956 91420 5020 91424
rect 4956 91364 4960 91420
rect 4960 91364 5016 91420
rect 5016 91364 5020 91420
rect 4956 91360 5020 91364
rect 5036 91420 5100 91424
rect 5036 91364 5040 91420
rect 5040 91364 5096 91420
rect 5096 91364 5100 91420
rect 5036 91360 5100 91364
rect 5116 91420 5180 91424
rect 5116 91364 5120 91420
rect 5120 91364 5176 91420
rect 5176 91364 5180 91420
rect 5116 91360 5180 91364
rect 106660 91420 106724 91424
rect 106660 91364 106664 91420
rect 106664 91364 106720 91420
rect 106720 91364 106724 91420
rect 106660 91360 106724 91364
rect 106740 91420 106804 91424
rect 106740 91364 106744 91420
rect 106744 91364 106800 91420
rect 106800 91364 106804 91420
rect 106740 91360 106804 91364
rect 106820 91420 106884 91424
rect 106820 91364 106824 91420
rect 106824 91364 106880 91420
rect 106880 91364 106884 91420
rect 106820 91360 106884 91364
rect 106900 91420 106964 91424
rect 106900 91364 106904 91420
rect 106904 91364 106960 91420
rect 106960 91364 106964 91420
rect 106900 91360 106964 91364
rect 4216 90876 4280 90880
rect 4216 90820 4220 90876
rect 4220 90820 4276 90876
rect 4276 90820 4280 90876
rect 4216 90816 4280 90820
rect 4296 90876 4360 90880
rect 4296 90820 4300 90876
rect 4300 90820 4356 90876
rect 4356 90820 4360 90876
rect 4296 90816 4360 90820
rect 4376 90876 4440 90880
rect 4376 90820 4380 90876
rect 4380 90820 4436 90876
rect 4436 90820 4440 90876
rect 4376 90816 4440 90820
rect 4456 90876 4520 90880
rect 4456 90820 4460 90876
rect 4460 90820 4516 90876
rect 4516 90820 4520 90876
rect 4456 90816 4520 90820
rect 105924 90876 105988 90880
rect 105924 90820 105928 90876
rect 105928 90820 105984 90876
rect 105984 90820 105988 90876
rect 105924 90816 105988 90820
rect 106004 90876 106068 90880
rect 106004 90820 106008 90876
rect 106008 90820 106064 90876
rect 106064 90820 106068 90876
rect 106004 90816 106068 90820
rect 106084 90876 106148 90880
rect 106084 90820 106088 90876
rect 106088 90820 106144 90876
rect 106144 90820 106148 90876
rect 106084 90816 106148 90820
rect 106164 90876 106228 90880
rect 106164 90820 106168 90876
rect 106168 90820 106224 90876
rect 106224 90820 106228 90876
rect 106164 90816 106228 90820
rect 4876 90332 4940 90336
rect 4876 90276 4880 90332
rect 4880 90276 4936 90332
rect 4936 90276 4940 90332
rect 4876 90272 4940 90276
rect 4956 90332 5020 90336
rect 4956 90276 4960 90332
rect 4960 90276 5016 90332
rect 5016 90276 5020 90332
rect 4956 90272 5020 90276
rect 5036 90332 5100 90336
rect 5036 90276 5040 90332
rect 5040 90276 5096 90332
rect 5096 90276 5100 90332
rect 5036 90272 5100 90276
rect 5116 90332 5180 90336
rect 5116 90276 5120 90332
rect 5120 90276 5176 90332
rect 5176 90276 5180 90332
rect 5116 90272 5180 90276
rect 106660 90332 106724 90336
rect 106660 90276 106664 90332
rect 106664 90276 106720 90332
rect 106720 90276 106724 90332
rect 106660 90272 106724 90276
rect 106740 90332 106804 90336
rect 106740 90276 106744 90332
rect 106744 90276 106800 90332
rect 106800 90276 106804 90332
rect 106740 90272 106804 90276
rect 106820 90332 106884 90336
rect 106820 90276 106824 90332
rect 106824 90276 106880 90332
rect 106880 90276 106884 90332
rect 106820 90272 106884 90276
rect 106900 90332 106964 90336
rect 106900 90276 106904 90332
rect 106904 90276 106960 90332
rect 106960 90276 106964 90332
rect 106900 90272 106964 90276
rect 4216 89788 4280 89792
rect 4216 89732 4220 89788
rect 4220 89732 4276 89788
rect 4276 89732 4280 89788
rect 4216 89728 4280 89732
rect 4296 89788 4360 89792
rect 4296 89732 4300 89788
rect 4300 89732 4356 89788
rect 4356 89732 4360 89788
rect 4296 89728 4360 89732
rect 4376 89788 4440 89792
rect 4376 89732 4380 89788
rect 4380 89732 4436 89788
rect 4436 89732 4440 89788
rect 4376 89728 4440 89732
rect 4456 89788 4520 89792
rect 4456 89732 4460 89788
rect 4460 89732 4516 89788
rect 4516 89732 4520 89788
rect 4456 89728 4520 89732
rect 105924 89788 105988 89792
rect 105924 89732 105928 89788
rect 105928 89732 105984 89788
rect 105984 89732 105988 89788
rect 105924 89728 105988 89732
rect 106004 89788 106068 89792
rect 106004 89732 106008 89788
rect 106008 89732 106064 89788
rect 106064 89732 106068 89788
rect 106004 89728 106068 89732
rect 106084 89788 106148 89792
rect 106084 89732 106088 89788
rect 106088 89732 106144 89788
rect 106144 89732 106148 89788
rect 106084 89728 106148 89732
rect 106164 89788 106228 89792
rect 106164 89732 106168 89788
rect 106168 89732 106224 89788
rect 106224 89732 106228 89788
rect 106164 89728 106228 89732
rect 4876 89244 4940 89248
rect 4876 89188 4880 89244
rect 4880 89188 4936 89244
rect 4936 89188 4940 89244
rect 4876 89184 4940 89188
rect 4956 89244 5020 89248
rect 4956 89188 4960 89244
rect 4960 89188 5016 89244
rect 5016 89188 5020 89244
rect 4956 89184 5020 89188
rect 5036 89244 5100 89248
rect 5036 89188 5040 89244
rect 5040 89188 5096 89244
rect 5096 89188 5100 89244
rect 5036 89184 5100 89188
rect 5116 89244 5180 89248
rect 5116 89188 5120 89244
rect 5120 89188 5176 89244
rect 5176 89188 5180 89244
rect 5116 89184 5180 89188
rect 106660 89244 106724 89248
rect 106660 89188 106664 89244
rect 106664 89188 106720 89244
rect 106720 89188 106724 89244
rect 106660 89184 106724 89188
rect 106740 89244 106804 89248
rect 106740 89188 106744 89244
rect 106744 89188 106800 89244
rect 106800 89188 106804 89244
rect 106740 89184 106804 89188
rect 106820 89244 106884 89248
rect 106820 89188 106824 89244
rect 106824 89188 106880 89244
rect 106880 89188 106884 89244
rect 106820 89184 106884 89188
rect 106900 89244 106964 89248
rect 106900 89188 106904 89244
rect 106904 89188 106960 89244
rect 106960 89188 106964 89244
rect 106900 89184 106964 89188
rect 4216 88700 4280 88704
rect 4216 88644 4220 88700
rect 4220 88644 4276 88700
rect 4276 88644 4280 88700
rect 4216 88640 4280 88644
rect 4296 88700 4360 88704
rect 4296 88644 4300 88700
rect 4300 88644 4356 88700
rect 4356 88644 4360 88700
rect 4296 88640 4360 88644
rect 4376 88700 4440 88704
rect 4376 88644 4380 88700
rect 4380 88644 4436 88700
rect 4436 88644 4440 88700
rect 4376 88640 4440 88644
rect 4456 88700 4520 88704
rect 4456 88644 4460 88700
rect 4460 88644 4516 88700
rect 4516 88644 4520 88700
rect 4456 88640 4520 88644
rect 105924 88700 105988 88704
rect 105924 88644 105928 88700
rect 105928 88644 105984 88700
rect 105984 88644 105988 88700
rect 105924 88640 105988 88644
rect 106004 88700 106068 88704
rect 106004 88644 106008 88700
rect 106008 88644 106064 88700
rect 106064 88644 106068 88700
rect 106004 88640 106068 88644
rect 106084 88700 106148 88704
rect 106084 88644 106088 88700
rect 106088 88644 106144 88700
rect 106144 88644 106148 88700
rect 106084 88640 106148 88644
rect 106164 88700 106228 88704
rect 106164 88644 106168 88700
rect 106168 88644 106224 88700
rect 106224 88644 106228 88700
rect 106164 88640 106228 88644
rect 4876 88156 4940 88160
rect 4876 88100 4880 88156
rect 4880 88100 4936 88156
rect 4936 88100 4940 88156
rect 4876 88096 4940 88100
rect 4956 88156 5020 88160
rect 4956 88100 4960 88156
rect 4960 88100 5016 88156
rect 5016 88100 5020 88156
rect 4956 88096 5020 88100
rect 5036 88156 5100 88160
rect 5036 88100 5040 88156
rect 5040 88100 5096 88156
rect 5096 88100 5100 88156
rect 5036 88096 5100 88100
rect 5116 88156 5180 88160
rect 5116 88100 5120 88156
rect 5120 88100 5176 88156
rect 5176 88100 5180 88156
rect 5116 88096 5180 88100
rect 106660 88156 106724 88160
rect 106660 88100 106664 88156
rect 106664 88100 106720 88156
rect 106720 88100 106724 88156
rect 106660 88096 106724 88100
rect 106740 88156 106804 88160
rect 106740 88100 106744 88156
rect 106744 88100 106800 88156
rect 106800 88100 106804 88156
rect 106740 88096 106804 88100
rect 106820 88156 106884 88160
rect 106820 88100 106824 88156
rect 106824 88100 106880 88156
rect 106880 88100 106884 88156
rect 106820 88096 106884 88100
rect 106900 88156 106964 88160
rect 106900 88100 106904 88156
rect 106904 88100 106960 88156
rect 106960 88100 106964 88156
rect 106900 88096 106964 88100
rect 4216 87612 4280 87616
rect 4216 87556 4220 87612
rect 4220 87556 4276 87612
rect 4276 87556 4280 87612
rect 4216 87552 4280 87556
rect 4296 87612 4360 87616
rect 4296 87556 4300 87612
rect 4300 87556 4356 87612
rect 4356 87556 4360 87612
rect 4296 87552 4360 87556
rect 4376 87612 4440 87616
rect 4376 87556 4380 87612
rect 4380 87556 4436 87612
rect 4436 87556 4440 87612
rect 4376 87552 4440 87556
rect 4456 87612 4520 87616
rect 4456 87556 4460 87612
rect 4460 87556 4516 87612
rect 4516 87556 4520 87612
rect 4456 87552 4520 87556
rect 105924 87612 105988 87616
rect 105924 87556 105928 87612
rect 105928 87556 105984 87612
rect 105984 87556 105988 87612
rect 105924 87552 105988 87556
rect 106004 87612 106068 87616
rect 106004 87556 106008 87612
rect 106008 87556 106064 87612
rect 106064 87556 106068 87612
rect 106004 87552 106068 87556
rect 106084 87612 106148 87616
rect 106084 87556 106088 87612
rect 106088 87556 106144 87612
rect 106144 87556 106148 87612
rect 106084 87552 106148 87556
rect 106164 87612 106228 87616
rect 106164 87556 106168 87612
rect 106168 87556 106224 87612
rect 106224 87556 106228 87612
rect 106164 87552 106228 87556
rect 4876 87068 4940 87072
rect 4876 87012 4880 87068
rect 4880 87012 4936 87068
rect 4936 87012 4940 87068
rect 4876 87008 4940 87012
rect 4956 87068 5020 87072
rect 4956 87012 4960 87068
rect 4960 87012 5016 87068
rect 5016 87012 5020 87068
rect 4956 87008 5020 87012
rect 5036 87068 5100 87072
rect 5036 87012 5040 87068
rect 5040 87012 5096 87068
rect 5096 87012 5100 87068
rect 5036 87008 5100 87012
rect 5116 87068 5180 87072
rect 5116 87012 5120 87068
rect 5120 87012 5176 87068
rect 5176 87012 5180 87068
rect 5116 87008 5180 87012
rect 106660 87068 106724 87072
rect 106660 87012 106664 87068
rect 106664 87012 106720 87068
rect 106720 87012 106724 87068
rect 106660 87008 106724 87012
rect 106740 87068 106804 87072
rect 106740 87012 106744 87068
rect 106744 87012 106800 87068
rect 106800 87012 106804 87068
rect 106740 87008 106804 87012
rect 106820 87068 106884 87072
rect 106820 87012 106824 87068
rect 106824 87012 106880 87068
rect 106880 87012 106884 87068
rect 106820 87008 106884 87012
rect 106900 87068 106964 87072
rect 106900 87012 106904 87068
rect 106904 87012 106960 87068
rect 106960 87012 106964 87068
rect 106900 87008 106964 87012
rect 4216 86524 4280 86528
rect 4216 86468 4220 86524
rect 4220 86468 4276 86524
rect 4276 86468 4280 86524
rect 4216 86464 4280 86468
rect 4296 86524 4360 86528
rect 4296 86468 4300 86524
rect 4300 86468 4356 86524
rect 4356 86468 4360 86524
rect 4296 86464 4360 86468
rect 4376 86524 4440 86528
rect 4376 86468 4380 86524
rect 4380 86468 4436 86524
rect 4436 86468 4440 86524
rect 4376 86464 4440 86468
rect 4456 86524 4520 86528
rect 4456 86468 4460 86524
rect 4460 86468 4516 86524
rect 4516 86468 4520 86524
rect 4456 86464 4520 86468
rect 105924 86524 105988 86528
rect 105924 86468 105928 86524
rect 105928 86468 105984 86524
rect 105984 86468 105988 86524
rect 105924 86464 105988 86468
rect 106004 86524 106068 86528
rect 106004 86468 106008 86524
rect 106008 86468 106064 86524
rect 106064 86468 106068 86524
rect 106004 86464 106068 86468
rect 106084 86524 106148 86528
rect 106084 86468 106088 86524
rect 106088 86468 106144 86524
rect 106144 86468 106148 86524
rect 106084 86464 106148 86468
rect 106164 86524 106228 86528
rect 106164 86468 106168 86524
rect 106168 86468 106224 86524
rect 106224 86468 106228 86524
rect 106164 86464 106228 86468
rect 4876 85980 4940 85984
rect 4876 85924 4880 85980
rect 4880 85924 4936 85980
rect 4936 85924 4940 85980
rect 4876 85920 4940 85924
rect 4956 85980 5020 85984
rect 4956 85924 4960 85980
rect 4960 85924 5016 85980
rect 5016 85924 5020 85980
rect 4956 85920 5020 85924
rect 5036 85980 5100 85984
rect 5036 85924 5040 85980
rect 5040 85924 5096 85980
rect 5096 85924 5100 85980
rect 5036 85920 5100 85924
rect 5116 85980 5180 85984
rect 5116 85924 5120 85980
rect 5120 85924 5176 85980
rect 5176 85924 5180 85980
rect 5116 85920 5180 85924
rect 106660 85980 106724 85984
rect 106660 85924 106664 85980
rect 106664 85924 106720 85980
rect 106720 85924 106724 85980
rect 106660 85920 106724 85924
rect 106740 85980 106804 85984
rect 106740 85924 106744 85980
rect 106744 85924 106800 85980
rect 106800 85924 106804 85980
rect 106740 85920 106804 85924
rect 106820 85980 106884 85984
rect 106820 85924 106824 85980
rect 106824 85924 106880 85980
rect 106880 85924 106884 85980
rect 106820 85920 106884 85924
rect 106900 85980 106964 85984
rect 106900 85924 106904 85980
rect 106904 85924 106960 85980
rect 106960 85924 106964 85980
rect 106900 85920 106964 85924
rect 4216 85436 4280 85440
rect 4216 85380 4220 85436
rect 4220 85380 4276 85436
rect 4276 85380 4280 85436
rect 4216 85376 4280 85380
rect 4296 85436 4360 85440
rect 4296 85380 4300 85436
rect 4300 85380 4356 85436
rect 4356 85380 4360 85436
rect 4296 85376 4360 85380
rect 4376 85436 4440 85440
rect 4376 85380 4380 85436
rect 4380 85380 4436 85436
rect 4436 85380 4440 85436
rect 4376 85376 4440 85380
rect 4456 85436 4520 85440
rect 4456 85380 4460 85436
rect 4460 85380 4516 85436
rect 4516 85380 4520 85436
rect 4456 85376 4520 85380
rect 105924 85436 105988 85440
rect 105924 85380 105928 85436
rect 105928 85380 105984 85436
rect 105984 85380 105988 85436
rect 105924 85376 105988 85380
rect 106004 85436 106068 85440
rect 106004 85380 106008 85436
rect 106008 85380 106064 85436
rect 106064 85380 106068 85436
rect 106004 85376 106068 85380
rect 106084 85436 106148 85440
rect 106084 85380 106088 85436
rect 106088 85380 106144 85436
rect 106144 85380 106148 85436
rect 106084 85376 106148 85380
rect 106164 85436 106228 85440
rect 106164 85380 106168 85436
rect 106168 85380 106224 85436
rect 106224 85380 106228 85436
rect 106164 85376 106228 85380
rect 4876 84892 4940 84896
rect 4876 84836 4880 84892
rect 4880 84836 4936 84892
rect 4936 84836 4940 84892
rect 4876 84832 4940 84836
rect 4956 84892 5020 84896
rect 4956 84836 4960 84892
rect 4960 84836 5016 84892
rect 5016 84836 5020 84892
rect 4956 84832 5020 84836
rect 5036 84892 5100 84896
rect 5036 84836 5040 84892
rect 5040 84836 5096 84892
rect 5096 84836 5100 84892
rect 5036 84832 5100 84836
rect 5116 84892 5180 84896
rect 5116 84836 5120 84892
rect 5120 84836 5176 84892
rect 5176 84836 5180 84892
rect 5116 84832 5180 84836
rect 106660 84892 106724 84896
rect 106660 84836 106664 84892
rect 106664 84836 106720 84892
rect 106720 84836 106724 84892
rect 106660 84832 106724 84836
rect 106740 84892 106804 84896
rect 106740 84836 106744 84892
rect 106744 84836 106800 84892
rect 106800 84836 106804 84892
rect 106740 84832 106804 84836
rect 106820 84892 106884 84896
rect 106820 84836 106824 84892
rect 106824 84836 106880 84892
rect 106880 84836 106884 84892
rect 106820 84832 106884 84836
rect 106900 84892 106964 84896
rect 106900 84836 106904 84892
rect 106904 84836 106960 84892
rect 106960 84836 106964 84892
rect 106900 84832 106964 84836
rect 4216 84348 4280 84352
rect 4216 84292 4220 84348
rect 4220 84292 4276 84348
rect 4276 84292 4280 84348
rect 4216 84288 4280 84292
rect 4296 84348 4360 84352
rect 4296 84292 4300 84348
rect 4300 84292 4356 84348
rect 4356 84292 4360 84348
rect 4296 84288 4360 84292
rect 4376 84348 4440 84352
rect 4376 84292 4380 84348
rect 4380 84292 4436 84348
rect 4436 84292 4440 84348
rect 4376 84288 4440 84292
rect 4456 84348 4520 84352
rect 4456 84292 4460 84348
rect 4460 84292 4516 84348
rect 4516 84292 4520 84348
rect 4456 84288 4520 84292
rect 105924 84348 105988 84352
rect 105924 84292 105928 84348
rect 105928 84292 105984 84348
rect 105984 84292 105988 84348
rect 105924 84288 105988 84292
rect 106004 84348 106068 84352
rect 106004 84292 106008 84348
rect 106008 84292 106064 84348
rect 106064 84292 106068 84348
rect 106004 84288 106068 84292
rect 106084 84348 106148 84352
rect 106084 84292 106088 84348
rect 106088 84292 106144 84348
rect 106144 84292 106148 84348
rect 106084 84288 106148 84292
rect 106164 84348 106228 84352
rect 106164 84292 106168 84348
rect 106168 84292 106224 84348
rect 106224 84292 106228 84348
rect 106164 84288 106228 84292
rect 4876 83804 4940 83808
rect 4876 83748 4880 83804
rect 4880 83748 4936 83804
rect 4936 83748 4940 83804
rect 4876 83744 4940 83748
rect 4956 83804 5020 83808
rect 4956 83748 4960 83804
rect 4960 83748 5016 83804
rect 5016 83748 5020 83804
rect 4956 83744 5020 83748
rect 5036 83804 5100 83808
rect 5036 83748 5040 83804
rect 5040 83748 5096 83804
rect 5096 83748 5100 83804
rect 5036 83744 5100 83748
rect 5116 83804 5180 83808
rect 5116 83748 5120 83804
rect 5120 83748 5176 83804
rect 5176 83748 5180 83804
rect 5116 83744 5180 83748
rect 106660 83804 106724 83808
rect 106660 83748 106664 83804
rect 106664 83748 106720 83804
rect 106720 83748 106724 83804
rect 106660 83744 106724 83748
rect 106740 83804 106804 83808
rect 106740 83748 106744 83804
rect 106744 83748 106800 83804
rect 106800 83748 106804 83804
rect 106740 83744 106804 83748
rect 106820 83804 106884 83808
rect 106820 83748 106824 83804
rect 106824 83748 106880 83804
rect 106880 83748 106884 83804
rect 106820 83744 106884 83748
rect 106900 83804 106964 83808
rect 106900 83748 106904 83804
rect 106904 83748 106960 83804
rect 106960 83748 106964 83804
rect 106900 83744 106964 83748
rect 4216 83260 4280 83264
rect 4216 83204 4220 83260
rect 4220 83204 4276 83260
rect 4276 83204 4280 83260
rect 4216 83200 4280 83204
rect 4296 83260 4360 83264
rect 4296 83204 4300 83260
rect 4300 83204 4356 83260
rect 4356 83204 4360 83260
rect 4296 83200 4360 83204
rect 4376 83260 4440 83264
rect 4376 83204 4380 83260
rect 4380 83204 4436 83260
rect 4436 83204 4440 83260
rect 4376 83200 4440 83204
rect 4456 83260 4520 83264
rect 4456 83204 4460 83260
rect 4460 83204 4516 83260
rect 4516 83204 4520 83260
rect 4456 83200 4520 83204
rect 105924 83260 105988 83264
rect 105924 83204 105928 83260
rect 105928 83204 105984 83260
rect 105984 83204 105988 83260
rect 105924 83200 105988 83204
rect 106004 83260 106068 83264
rect 106004 83204 106008 83260
rect 106008 83204 106064 83260
rect 106064 83204 106068 83260
rect 106004 83200 106068 83204
rect 106084 83260 106148 83264
rect 106084 83204 106088 83260
rect 106088 83204 106144 83260
rect 106144 83204 106148 83260
rect 106084 83200 106148 83204
rect 106164 83260 106228 83264
rect 106164 83204 106168 83260
rect 106168 83204 106224 83260
rect 106224 83204 106228 83260
rect 106164 83200 106228 83204
rect 4876 82716 4940 82720
rect 4876 82660 4880 82716
rect 4880 82660 4936 82716
rect 4936 82660 4940 82716
rect 4876 82656 4940 82660
rect 4956 82716 5020 82720
rect 4956 82660 4960 82716
rect 4960 82660 5016 82716
rect 5016 82660 5020 82716
rect 4956 82656 5020 82660
rect 5036 82716 5100 82720
rect 5036 82660 5040 82716
rect 5040 82660 5096 82716
rect 5096 82660 5100 82716
rect 5036 82656 5100 82660
rect 5116 82716 5180 82720
rect 5116 82660 5120 82716
rect 5120 82660 5176 82716
rect 5176 82660 5180 82716
rect 5116 82656 5180 82660
rect 106660 82716 106724 82720
rect 106660 82660 106664 82716
rect 106664 82660 106720 82716
rect 106720 82660 106724 82716
rect 106660 82656 106724 82660
rect 106740 82716 106804 82720
rect 106740 82660 106744 82716
rect 106744 82660 106800 82716
rect 106800 82660 106804 82716
rect 106740 82656 106804 82660
rect 106820 82716 106884 82720
rect 106820 82660 106824 82716
rect 106824 82660 106880 82716
rect 106880 82660 106884 82716
rect 106820 82656 106884 82660
rect 106900 82716 106964 82720
rect 106900 82660 106904 82716
rect 106904 82660 106960 82716
rect 106960 82660 106964 82716
rect 106900 82656 106964 82660
rect 4216 82172 4280 82176
rect 4216 82116 4220 82172
rect 4220 82116 4276 82172
rect 4276 82116 4280 82172
rect 4216 82112 4280 82116
rect 4296 82172 4360 82176
rect 4296 82116 4300 82172
rect 4300 82116 4356 82172
rect 4356 82116 4360 82172
rect 4296 82112 4360 82116
rect 4376 82172 4440 82176
rect 4376 82116 4380 82172
rect 4380 82116 4436 82172
rect 4436 82116 4440 82172
rect 4376 82112 4440 82116
rect 4456 82172 4520 82176
rect 4456 82116 4460 82172
rect 4460 82116 4516 82172
rect 4516 82116 4520 82172
rect 4456 82112 4520 82116
rect 105924 82172 105988 82176
rect 105924 82116 105928 82172
rect 105928 82116 105984 82172
rect 105984 82116 105988 82172
rect 105924 82112 105988 82116
rect 106004 82172 106068 82176
rect 106004 82116 106008 82172
rect 106008 82116 106064 82172
rect 106064 82116 106068 82172
rect 106004 82112 106068 82116
rect 106084 82172 106148 82176
rect 106084 82116 106088 82172
rect 106088 82116 106144 82172
rect 106144 82116 106148 82172
rect 106084 82112 106148 82116
rect 106164 82172 106228 82176
rect 106164 82116 106168 82172
rect 106168 82116 106224 82172
rect 106224 82116 106228 82172
rect 106164 82112 106228 82116
rect 4876 81628 4940 81632
rect 4876 81572 4880 81628
rect 4880 81572 4936 81628
rect 4936 81572 4940 81628
rect 4876 81568 4940 81572
rect 4956 81628 5020 81632
rect 4956 81572 4960 81628
rect 4960 81572 5016 81628
rect 5016 81572 5020 81628
rect 4956 81568 5020 81572
rect 5036 81628 5100 81632
rect 5036 81572 5040 81628
rect 5040 81572 5096 81628
rect 5096 81572 5100 81628
rect 5036 81568 5100 81572
rect 5116 81628 5180 81632
rect 5116 81572 5120 81628
rect 5120 81572 5176 81628
rect 5176 81572 5180 81628
rect 5116 81568 5180 81572
rect 106660 81628 106724 81632
rect 106660 81572 106664 81628
rect 106664 81572 106720 81628
rect 106720 81572 106724 81628
rect 106660 81568 106724 81572
rect 106740 81628 106804 81632
rect 106740 81572 106744 81628
rect 106744 81572 106800 81628
rect 106800 81572 106804 81628
rect 106740 81568 106804 81572
rect 106820 81628 106884 81632
rect 106820 81572 106824 81628
rect 106824 81572 106880 81628
rect 106880 81572 106884 81628
rect 106820 81568 106884 81572
rect 106900 81628 106964 81632
rect 106900 81572 106904 81628
rect 106904 81572 106960 81628
rect 106960 81572 106964 81628
rect 106900 81568 106964 81572
rect 4216 81084 4280 81088
rect 4216 81028 4220 81084
rect 4220 81028 4276 81084
rect 4276 81028 4280 81084
rect 4216 81024 4280 81028
rect 4296 81084 4360 81088
rect 4296 81028 4300 81084
rect 4300 81028 4356 81084
rect 4356 81028 4360 81084
rect 4296 81024 4360 81028
rect 4376 81084 4440 81088
rect 4376 81028 4380 81084
rect 4380 81028 4436 81084
rect 4436 81028 4440 81084
rect 4376 81024 4440 81028
rect 4456 81084 4520 81088
rect 4456 81028 4460 81084
rect 4460 81028 4516 81084
rect 4516 81028 4520 81084
rect 4456 81024 4520 81028
rect 105924 81084 105988 81088
rect 105924 81028 105928 81084
rect 105928 81028 105984 81084
rect 105984 81028 105988 81084
rect 105924 81024 105988 81028
rect 106004 81084 106068 81088
rect 106004 81028 106008 81084
rect 106008 81028 106064 81084
rect 106064 81028 106068 81084
rect 106004 81024 106068 81028
rect 106084 81084 106148 81088
rect 106084 81028 106088 81084
rect 106088 81028 106144 81084
rect 106144 81028 106148 81084
rect 106084 81024 106148 81028
rect 106164 81084 106228 81088
rect 106164 81028 106168 81084
rect 106168 81028 106224 81084
rect 106224 81028 106228 81084
rect 106164 81024 106228 81028
rect 4876 80540 4940 80544
rect 4876 80484 4880 80540
rect 4880 80484 4936 80540
rect 4936 80484 4940 80540
rect 4876 80480 4940 80484
rect 4956 80540 5020 80544
rect 4956 80484 4960 80540
rect 4960 80484 5016 80540
rect 5016 80484 5020 80540
rect 4956 80480 5020 80484
rect 5036 80540 5100 80544
rect 5036 80484 5040 80540
rect 5040 80484 5096 80540
rect 5096 80484 5100 80540
rect 5036 80480 5100 80484
rect 5116 80540 5180 80544
rect 5116 80484 5120 80540
rect 5120 80484 5176 80540
rect 5176 80484 5180 80540
rect 5116 80480 5180 80484
rect 106660 80540 106724 80544
rect 106660 80484 106664 80540
rect 106664 80484 106720 80540
rect 106720 80484 106724 80540
rect 106660 80480 106724 80484
rect 106740 80540 106804 80544
rect 106740 80484 106744 80540
rect 106744 80484 106800 80540
rect 106800 80484 106804 80540
rect 106740 80480 106804 80484
rect 106820 80540 106884 80544
rect 106820 80484 106824 80540
rect 106824 80484 106880 80540
rect 106880 80484 106884 80540
rect 106820 80480 106884 80484
rect 106900 80540 106964 80544
rect 106900 80484 106904 80540
rect 106904 80484 106960 80540
rect 106960 80484 106964 80540
rect 106900 80480 106964 80484
rect 4216 79996 4280 80000
rect 4216 79940 4220 79996
rect 4220 79940 4276 79996
rect 4276 79940 4280 79996
rect 4216 79936 4280 79940
rect 4296 79996 4360 80000
rect 4296 79940 4300 79996
rect 4300 79940 4356 79996
rect 4356 79940 4360 79996
rect 4296 79936 4360 79940
rect 4376 79996 4440 80000
rect 4376 79940 4380 79996
rect 4380 79940 4436 79996
rect 4436 79940 4440 79996
rect 4376 79936 4440 79940
rect 4456 79996 4520 80000
rect 4456 79940 4460 79996
rect 4460 79940 4516 79996
rect 4516 79940 4520 79996
rect 4456 79936 4520 79940
rect 105924 79996 105988 80000
rect 105924 79940 105928 79996
rect 105928 79940 105984 79996
rect 105984 79940 105988 79996
rect 105924 79936 105988 79940
rect 106004 79996 106068 80000
rect 106004 79940 106008 79996
rect 106008 79940 106064 79996
rect 106064 79940 106068 79996
rect 106004 79936 106068 79940
rect 106084 79996 106148 80000
rect 106084 79940 106088 79996
rect 106088 79940 106144 79996
rect 106144 79940 106148 79996
rect 106084 79936 106148 79940
rect 106164 79996 106228 80000
rect 106164 79940 106168 79996
rect 106168 79940 106224 79996
rect 106224 79940 106228 79996
rect 106164 79936 106228 79940
rect 31614 79868 31678 79932
rect 36286 79928 36350 79932
rect 36286 79872 36322 79928
rect 36322 79872 36350 79928
rect 36286 79868 36350 79872
rect 38622 79928 38686 79932
rect 38622 79872 38658 79928
rect 38658 79872 38686 79928
rect 38622 79868 38686 79872
rect 39790 79928 39854 79932
rect 39790 79872 39818 79928
rect 39818 79872 39854 79928
rect 39790 79868 39854 79872
rect 40958 79928 41022 79932
rect 40958 79872 41014 79928
rect 41014 79872 41022 79928
rect 40958 79868 41022 79872
rect 90814 79868 90878 79932
rect 30446 79732 30510 79796
rect 32782 79732 32846 79796
rect 25774 79596 25838 79660
rect 37454 79596 37518 79660
rect 24606 79460 24670 79524
rect 29278 79460 29342 79524
rect 30446 79520 30510 79524
rect 30446 79464 30470 79520
rect 30470 79464 30510 79520
rect 30446 79460 30510 79464
rect 31614 79520 31678 79524
rect 31614 79464 31630 79520
rect 31630 79464 31678 79520
rect 31614 79460 31678 79464
rect 33950 79520 34014 79524
rect 33950 79464 33966 79520
rect 33966 79464 34014 79520
rect 33950 79460 34014 79464
rect 35112 79460 35176 79524
rect 42126 79520 42190 79524
rect 42126 79464 42154 79520
rect 42154 79464 42190 79520
rect 42126 79460 42190 79464
rect 43294 79520 43358 79524
rect 43294 79464 43314 79520
rect 43314 79464 43358 79520
rect 43294 79460 43358 79464
rect 90680 79460 90744 79524
rect 4876 79452 4940 79456
rect 4876 79396 4880 79452
rect 4880 79396 4936 79452
rect 4936 79396 4940 79452
rect 4876 79392 4940 79396
rect 4956 79452 5020 79456
rect 4956 79396 4960 79452
rect 4960 79396 5016 79452
rect 5016 79396 5020 79452
rect 4956 79392 5020 79396
rect 5036 79452 5100 79456
rect 5036 79396 5040 79452
rect 5040 79396 5096 79452
rect 5096 79396 5100 79452
rect 5036 79392 5100 79396
rect 5116 79452 5180 79456
rect 5116 79396 5120 79452
rect 5120 79396 5176 79452
rect 5176 79396 5180 79452
rect 5116 79392 5180 79396
rect 106660 79452 106724 79456
rect 106660 79396 106664 79452
rect 106664 79396 106720 79452
rect 106720 79396 106724 79452
rect 106660 79392 106724 79396
rect 106740 79452 106804 79456
rect 106740 79396 106744 79452
rect 106744 79396 106800 79452
rect 106800 79396 106804 79452
rect 106740 79392 106804 79396
rect 106820 79452 106884 79456
rect 106820 79396 106824 79452
rect 106824 79396 106880 79452
rect 106880 79396 106884 79452
rect 106820 79392 106884 79396
rect 106900 79452 106964 79456
rect 106900 79396 106904 79452
rect 106904 79396 106960 79452
rect 106960 79396 106964 79452
rect 106900 79392 106964 79396
rect 26924 79324 26988 79388
rect 23428 79188 23492 79252
rect 4216 78908 4280 78912
rect 4216 78852 4220 78908
rect 4220 78852 4276 78908
rect 4276 78852 4280 78908
rect 4216 78848 4280 78852
rect 4296 78908 4360 78912
rect 4296 78852 4300 78908
rect 4300 78852 4356 78908
rect 4356 78852 4360 78908
rect 4296 78848 4360 78852
rect 4376 78908 4440 78912
rect 4376 78852 4380 78908
rect 4380 78852 4436 78908
rect 4436 78852 4440 78908
rect 4376 78848 4440 78852
rect 4456 78908 4520 78912
rect 4456 78852 4460 78908
rect 4460 78852 4516 78908
rect 4516 78852 4520 78908
rect 4456 78848 4520 78852
rect 105924 78908 105988 78912
rect 105924 78852 105928 78908
rect 105928 78852 105984 78908
rect 105984 78852 105988 78908
rect 105924 78848 105988 78852
rect 106004 78908 106068 78912
rect 106004 78852 106008 78908
rect 106008 78852 106064 78908
rect 106064 78852 106068 78908
rect 106004 78848 106068 78852
rect 106084 78908 106148 78912
rect 106084 78852 106088 78908
rect 106088 78852 106144 78908
rect 106144 78852 106148 78908
rect 106084 78848 106148 78852
rect 106164 78908 106228 78912
rect 106164 78852 106168 78908
rect 106168 78852 106224 78908
rect 106224 78852 106228 78908
rect 106164 78848 106228 78852
rect 23428 78780 23492 78844
rect 4876 78364 4940 78368
rect 4876 78308 4880 78364
rect 4880 78308 4936 78364
rect 4936 78308 4940 78364
rect 4876 78304 4940 78308
rect 4956 78364 5020 78368
rect 4956 78308 4960 78364
rect 4960 78308 5016 78364
rect 5016 78308 5020 78364
rect 4956 78304 5020 78308
rect 5036 78364 5100 78368
rect 5036 78308 5040 78364
rect 5040 78308 5096 78364
rect 5096 78308 5100 78364
rect 5036 78304 5100 78308
rect 5116 78364 5180 78368
rect 5116 78308 5120 78364
rect 5120 78308 5176 78364
rect 5176 78308 5180 78364
rect 5116 78304 5180 78308
rect 106660 78364 106724 78368
rect 106660 78308 106664 78364
rect 106664 78308 106720 78364
rect 106720 78308 106724 78364
rect 106660 78304 106724 78308
rect 106740 78364 106804 78368
rect 106740 78308 106744 78364
rect 106744 78308 106800 78364
rect 106800 78308 106804 78364
rect 106740 78304 106804 78308
rect 106820 78364 106884 78368
rect 106820 78308 106824 78364
rect 106824 78308 106880 78364
rect 106880 78308 106884 78364
rect 106820 78304 106884 78308
rect 106900 78364 106964 78368
rect 106900 78308 106904 78364
rect 106904 78308 106960 78364
rect 106960 78308 106964 78364
rect 106900 78304 106964 78308
rect 16068 78024 16132 78028
rect 16068 77968 16082 78024
rect 16082 77968 16132 78024
rect 16068 77964 16132 77968
rect 4216 77820 4280 77824
rect 4216 77764 4220 77820
rect 4220 77764 4276 77820
rect 4276 77764 4280 77820
rect 4216 77760 4280 77764
rect 4296 77820 4360 77824
rect 4296 77764 4300 77820
rect 4300 77764 4356 77820
rect 4356 77764 4360 77820
rect 4296 77760 4360 77764
rect 4376 77820 4440 77824
rect 4376 77764 4380 77820
rect 4380 77764 4436 77820
rect 4436 77764 4440 77820
rect 4376 77760 4440 77764
rect 4456 77820 4520 77824
rect 4456 77764 4460 77820
rect 4460 77764 4516 77820
rect 4516 77764 4520 77820
rect 4456 77760 4520 77764
rect 34936 77820 35000 77824
rect 34936 77764 34940 77820
rect 34940 77764 34996 77820
rect 34996 77764 35000 77820
rect 34936 77760 35000 77764
rect 35016 77820 35080 77824
rect 35016 77764 35020 77820
rect 35020 77764 35076 77820
rect 35076 77764 35080 77820
rect 35016 77760 35080 77764
rect 35096 77820 35160 77824
rect 35096 77764 35100 77820
rect 35100 77764 35156 77820
rect 35156 77764 35160 77820
rect 35096 77760 35160 77764
rect 35176 77820 35240 77824
rect 35176 77764 35180 77820
rect 35180 77764 35236 77820
rect 35236 77764 35240 77820
rect 35176 77760 35240 77764
rect 65656 77820 65720 77824
rect 65656 77764 65660 77820
rect 65660 77764 65716 77820
rect 65716 77764 65720 77820
rect 65656 77760 65720 77764
rect 65736 77820 65800 77824
rect 65736 77764 65740 77820
rect 65740 77764 65796 77820
rect 65796 77764 65800 77820
rect 65736 77760 65800 77764
rect 65816 77820 65880 77824
rect 65816 77764 65820 77820
rect 65820 77764 65876 77820
rect 65876 77764 65880 77820
rect 65816 77760 65880 77764
rect 65896 77820 65960 77824
rect 65896 77764 65900 77820
rect 65900 77764 65956 77820
rect 65956 77764 65960 77820
rect 65896 77760 65960 77764
rect 96376 77820 96440 77824
rect 96376 77764 96380 77820
rect 96380 77764 96436 77820
rect 96436 77764 96440 77820
rect 96376 77760 96440 77764
rect 96456 77820 96520 77824
rect 96456 77764 96460 77820
rect 96460 77764 96516 77820
rect 96516 77764 96520 77820
rect 96456 77760 96520 77764
rect 96536 77820 96600 77824
rect 96536 77764 96540 77820
rect 96540 77764 96596 77820
rect 96596 77764 96600 77820
rect 96536 77760 96600 77764
rect 96616 77820 96680 77824
rect 96616 77764 96620 77820
rect 96620 77764 96676 77820
rect 96676 77764 96680 77820
rect 96616 77760 96680 77764
rect 105924 77820 105988 77824
rect 105924 77764 105928 77820
rect 105928 77764 105984 77820
rect 105984 77764 105988 77820
rect 105924 77760 105988 77764
rect 106004 77820 106068 77824
rect 106004 77764 106008 77820
rect 106008 77764 106064 77820
rect 106064 77764 106068 77820
rect 106004 77760 106068 77764
rect 106084 77820 106148 77824
rect 106084 77764 106088 77820
rect 106088 77764 106144 77820
rect 106144 77764 106148 77820
rect 106084 77760 106148 77764
rect 106164 77820 106228 77824
rect 106164 77764 106168 77820
rect 106168 77764 106224 77820
rect 106224 77764 106228 77820
rect 106164 77760 106228 77764
rect 28212 77752 28276 77756
rect 28212 77696 28226 77752
rect 28226 77696 28276 77752
rect 28212 77692 28276 77696
rect 4876 77276 4940 77280
rect 4876 77220 4880 77276
rect 4880 77220 4936 77276
rect 4936 77220 4940 77276
rect 4876 77216 4940 77220
rect 4956 77276 5020 77280
rect 4956 77220 4960 77276
rect 4960 77220 5016 77276
rect 5016 77220 5020 77276
rect 4956 77216 5020 77220
rect 5036 77276 5100 77280
rect 5036 77220 5040 77276
rect 5040 77220 5096 77276
rect 5096 77220 5100 77276
rect 5036 77216 5100 77220
rect 5116 77276 5180 77280
rect 5116 77220 5120 77276
rect 5120 77220 5176 77276
rect 5176 77220 5180 77276
rect 5116 77216 5180 77220
rect 35596 77276 35660 77280
rect 35596 77220 35600 77276
rect 35600 77220 35656 77276
rect 35656 77220 35660 77276
rect 35596 77216 35660 77220
rect 35676 77276 35740 77280
rect 35676 77220 35680 77276
rect 35680 77220 35736 77276
rect 35736 77220 35740 77276
rect 35676 77216 35740 77220
rect 35756 77276 35820 77280
rect 35756 77220 35760 77276
rect 35760 77220 35816 77276
rect 35816 77220 35820 77276
rect 35756 77216 35820 77220
rect 35836 77276 35900 77280
rect 35836 77220 35840 77276
rect 35840 77220 35896 77276
rect 35896 77220 35900 77276
rect 35836 77216 35900 77220
rect 66316 77276 66380 77280
rect 66316 77220 66320 77276
rect 66320 77220 66376 77276
rect 66376 77220 66380 77276
rect 66316 77216 66380 77220
rect 66396 77276 66460 77280
rect 66396 77220 66400 77276
rect 66400 77220 66456 77276
rect 66456 77220 66460 77276
rect 66396 77216 66460 77220
rect 66476 77276 66540 77280
rect 66476 77220 66480 77276
rect 66480 77220 66536 77276
rect 66536 77220 66540 77276
rect 66476 77216 66540 77220
rect 66556 77276 66620 77280
rect 66556 77220 66560 77276
rect 66560 77220 66616 77276
rect 66616 77220 66620 77276
rect 66556 77216 66620 77220
rect 97036 77276 97100 77280
rect 97036 77220 97040 77276
rect 97040 77220 97096 77276
rect 97096 77220 97100 77276
rect 97036 77216 97100 77220
rect 97116 77276 97180 77280
rect 97116 77220 97120 77276
rect 97120 77220 97176 77276
rect 97176 77220 97180 77276
rect 97116 77216 97180 77220
rect 97196 77276 97260 77280
rect 97196 77220 97200 77276
rect 97200 77220 97256 77276
rect 97256 77220 97260 77276
rect 97196 77216 97260 77220
rect 97276 77276 97340 77280
rect 97276 77220 97280 77276
rect 97280 77220 97336 77276
rect 97336 77220 97340 77276
rect 97276 77216 97340 77220
rect 106660 77276 106724 77280
rect 106660 77220 106664 77276
rect 106664 77220 106720 77276
rect 106720 77220 106724 77276
rect 106660 77216 106724 77220
rect 106740 77276 106804 77280
rect 106740 77220 106744 77276
rect 106744 77220 106800 77276
rect 106800 77220 106804 77276
rect 106740 77216 106804 77220
rect 106820 77276 106884 77280
rect 106820 77220 106824 77276
rect 106824 77220 106880 77276
rect 106880 77220 106884 77276
rect 106820 77216 106884 77220
rect 106900 77276 106964 77280
rect 106900 77220 106904 77276
rect 106904 77220 106960 77276
rect 106960 77220 106964 77276
rect 106900 77216 106964 77220
rect 90404 77148 90468 77212
rect 4216 76732 4280 76736
rect 4216 76676 4220 76732
rect 4220 76676 4276 76732
rect 4276 76676 4280 76732
rect 4216 76672 4280 76676
rect 4296 76732 4360 76736
rect 4296 76676 4300 76732
rect 4300 76676 4356 76732
rect 4356 76676 4360 76732
rect 4296 76672 4360 76676
rect 4376 76732 4440 76736
rect 4376 76676 4380 76732
rect 4380 76676 4436 76732
rect 4436 76676 4440 76732
rect 4376 76672 4440 76676
rect 4456 76732 4520 76736
rect 4456 76676 4460 76732
rect 4460 76676 4516 76732
rect 4516 76676 4520 76732
rect 4456 76672 4520 76676
rect 34936 76732 35000 76736
rect 34936 76676 34940 76732
rect 34940 76676 34996 76732
rect 34996 76676 35000 76732
rect 34936 76672 35000 76676
rect 35016 76732 35080 76736
rect 35016 76676 35020 76732
rect 35020 76676 35076 76732
rect 35076 76676 35080 76732
rect 35016 76672 35080 76676
rect 35096 76732 35160 76736
rect 35096 76676 35100 76732
rect 35100 76676 35156 76732
rect 35156 76676 35160 76732
rect 35096 76672 35160 76676
rect 35176 76732 35240 76736
rect 35176 76676 35180 76732
rect 35180 76676 35236 76732
rect 35236 76676 35240 76732
rect 35176 76672 35240 76676
rect 65656 76732 65720 76736
rect 65656 76676 65660 76732
rect 65660 76676 65716 76732
rect 65716 76676 65720 76732
rect 65656 76672 65720 76676
rect 65736 76732 65800 76736
rect 65736 76676 65740 76732
rect 65740 76676 65796 76732
rect 65796 76676 65800 76732
rect 65736 76672 65800 76676
rect 65816 76732 65880 76736
rect 65816 76676 65820 76732
rect 65820 76676 65876 76732
rect 65876 76676 65880 76732
rect 65816 76672 65880 76676
rect 65896 76732 65960 76736
rect 65896 76676 65900 76732
rect 65900 76676 65956 76732
rect 65956 76676 65960 76732
rect 65896 76672 65960 76676
rect 96376 76732 96440 76736
rect 96376 76676 96380 76732
rect 96380 76676 96436 76732
rect 96436 76676 96440 76732
rect 96376 76672 96440 76676
rect 96456 76732 96520 76736
rect 96456 76676 96460 76732
rect 96460 76676 96516 76732
rect 96516 76676 96520 76732
rect 96456 76672 96520 76676
rect 96536 76732 96600 76736
rect 96536 76676 96540 76732
rect 96540 76676 96596 76732
rect 96596 76676 96600 76732
rect 96536 76672 96600 76676
rect 96616 76732 96680 76736
rect 96616 76676 96620 76732
rect 96620 76676 96676 76732
rect 96676 76676 96680 76732
rect 96616 76672 96680 76676
rect 4876 76188 4940 76192
rect 4876 76132 4880 76188
rect 4880 76132 4936 76188
rect 4936 76132 4940 76188
rect 4876 76128 4940 76132
rect 4956 76188 5020 76192
rect 4956 76132 4960 76188
rect 4960 76132 5016 76188
rect 5016 76132 5020 76188
rect 4956 76128 5020 76132
rect 5036 76188 5100 76192
rect 5036 76132 5040 76188
rect 5040 76132 5096 76188
rect 5096 76132 5100 76188
rect 5036 76128 5100 76132
rect 5116 76188 5180 76192
rect 5116 76132 5120 76188
rect 5120 76132 5176 76188
rect 5176 76132 5180 76188
rect 5116 76128 5180 76132
rect 35596 76188 35660 76192
rect 35596 76132 35600 76188
rect 35600 76132 35656 76188
rect 35656 76132 35660 76188
rect 35596 76128 35660 76132
rect 35676 76188 35740 76192
rect 35676 76132 35680 76188
rect 35680 76132 35736 76188
rect 35736 76132 35740 76188
rect 35676 76128 35740 76132
rect 35756 76188 35820 76192
rect 35756 76132 35760 76188
rect 35760 76132 35816 76188
rect 35816 76132 35820 76188
rect 35756 76128 35820 76132
rect 35836 76188 35900 76192
rect 35836 76132 35840 76188
rect 35840 76132 35896 76188
rect 35896 76132 35900 76188
rect 35836 76128 35900 76132
rect 66316 76188 66380 76192
rect 66316 76132 66320 76188
rect 66320 76132 66376 76188
rect 66376 76132 66380 76188
rect 66316 76128 66380 76132
rect 66396 76188 66460 76192
rect 66396 76132 66400 76188
rect 66400 76132 66456 76188
rect 66456 76132 66460 76188
rect 66396 76128 66460 76132
rect 66476 76188 66540 76192
rect 66476 76132 66480 76188
rect 66480 76132 66536 76188
rect 66536 76132 66540 76188
rect 66476 76128 66540 76132
rect 66556 76188 66620 76192
rect 66556 76132 66560 76188
rect 66560 76132 66616 76188
rect 66616 76132 66620 76188
rect 66556 76128 66620 76132
rect 97036 76188 97100 76192
rect 97036 76132 97040 76188
rect 97040 76132 97096 76188
rect 97096 76132 97100 76188
rect 97036 76128 97100 76132
rect 97116 76188 97180 76192
rect 97116 76132 97120 76188
rect 97120 76132 97176 76188
rect 97176 76132 97180 76188
rect 97116 76128 97180 76132
rect 97196 76188 97260 76192
rect 97196 76132 97200 76188
rect 97200 76132 97256 76188
rect 97256 76132 97260 76188
rect 97196 76128 97260 76132
rect 97276 76188 97340 76192
rect 97276 76132 97280 76188
rect 97280 76132 97336 76188
rect 97336 76132 97340 76188
rect 97276 76128 97340 76132
rect 4216 75644 4280 75648
rect 4216 75588 4220 75644
rect 4220 75588 4276 75644
rect 4276 75588 4280 75644
rect 4216 75584 4280 75588
rect 4296 75644 4360 75648
rect 4296 75588 4300 75644
rect 4300 75588 4356 75644
rect 4356 75588 4360 75644
rect 4296 75584 4360 75588
rect 4376 75644 4440 75648
rect 4376 75588 4380 75644
rect 4380 75588 4436 75644
rect 4436 75588 4440 75644
rect 4376 75584 4440 75588
rect 4456 75644 4520 75648
rect 4456 75588 4460 75644
rect 4460 75588 4516 75644
rect 4516 75588 4520 75644
rect 4456 75584 4520 75588
rect 34936 75644 35000 75648
rect 34936 75588 34940 75644
rect 34940 75588 34996 75644
rect 34996 75588 35000 75644
rect 34936 75584 35000 75588
rect 35016 75644 35080 75648
rect 35016 75588 35020 75644
rect 35020 75588 35076 75644
rect 35076 75588 35080 75644
rect 35016 75584 35080 75588
rect 35096 75644 35160 75648
rect 35096 75588 35100 75644
rect 35100 75588 35156 75644
rect 35156 75588 35160 75644
rect 35096 75584 35160 75588
rect 35176 75644 35240 75648
rect 35176 75588 35180 75644
rect 35180 75588 35236 75644
rect 35236 75588 35240 75644
rect 35176 75584 35240 75588
rect 65656 75644 65720 75648
rect 65656 75588 65660 75644
rect 65660 75588 65716 75644
rect 65716 75588 65720 75644
rect 65656 75584 65720 75588
rect 65736 75644 65800 75648
rect 65736 75588 65740 75644
rect 65740 75588 65796 75644
rect 65796 75588 65800 75644
rect 65736 75584 65800 75588
rect 65816 75644 65880 75648
rect 65816 75588 65820 75644
rect 65820 75588 65876 75644
rect 65876 75588 65880 75644
rect 65816 75584 65880 75588
rect 65896 75644 65960 75648
rect 65896 75588 65900 75644
rect 65900 75588 65956 75644
rect 65956 75588 65960 75644
rect 65896 75584 65960 75588
rect 96376 75644 96440 75648
rect 96376 75588 96380 75644
rect 96380 75588 96436 75644
rect 96436 75588 96440 75644
rect 96376 75584 96440 75588
rect 96456 75644 96520 75648
rect 96456 75588 96460 75644
rect 96460 75588 96516 75644
rect 96516 75588 96520 75644
rect 96456 75584 96520 75588
rect 96536 75644 96600 75648
rect 96536 75588 96540 75644
rect 96540 75588 96596 75644
rect 96596 75588 96600 75644
rect 96536 75584 96600 75588
rect 96616 75644 96680 75648
rect 96616 75588 96620 75644
rect 96620 75588 96676 75644
rect 96676 75588 96680 75644
rect 96616 75584 96680 75588
rect 4876 75100 4940 75104
rect 4876 75044 4880 75100
rect 4880 75044 4936 75100
rect 4936 75044 4940 75100
rect 4876 75040 4940 75044
rect 4956 75100 5020 75104
rect 4956 75044 4960 75100
rect 4960 75044 5016 75100
rect 5016 75044 5020 75100
rect 4956 75040 5020 75044
rect 5036 75100 5100 75104
rect 5036 75044 5040 75100
rect 5040 75044 5096 75100
rect 5096 75044 5100 75100
rect 5036 75040 5100 75044
rect 5116 75100 5180 75104
rect 5116 75044 5120 75100
rect 5120 75044 5176 75100
rect 5176 75044 5180 75100
rect 5116 75040 5180 75044
rect 35596 75100 35660 75104
rect 35596 75044 35600 75100
rect 35600 75044 35656 75100
rect 35656 75044 35660 75100
rect 35596 75040 35660 75044
rect 35676 75100 35740 75104
rect 35676 75044 35680 75100
rect 35680 75044 35736 75100
rect 35736 75044 35740 75100
rect 35676 75040 35740 75044
rect 35756 75100 35820 75104
rect 35756 75044 35760 75100
rect 35760 75044 35816 75100
rect 35816 75044 35820 75100
rect 35756 75040 35820 75044
rect 35836 75100 35900 75104
rect 35836 75044 35840 75100
rect 35840 75044 35896 75100
rect 35896 75044 35900 75100
rect 35836 75040 35900 75044
rect 66316 75100 66380 75104
rect 66316 75044 66320 75100
rect 66320 75044 66376 75100
rect 66376 75044 66380 75100
rect 66316 75040 66380 75044
rect 66396 75100 66460 75104
rect 66396 75044 66400 75100
rect 66400 75044 66456 75100
rect 66456 75044 66460 75100
rect 66396 75040 66460 75044
rect 66476 75100 66540 75104
rect 66476 75044 66480 75100
rect 66480 75044 66536 75100
rect 66536 75044 66540 75100
rect 66476 75040 66540 75044
rect 66556 75100 66620 75104
rect 66556 75044 66560 75100
rect 66560 75044 66616 75100
rect 66616 75044 66620 75100
rect 66556 75040 66620 75044
rect 97036 75100 97100 75104
rect 97036 75044 97040 75100
rect 97040 75044 97096 75100
rect 97096 75044 97100 75100
rect 97036 75040 97100 75044
rect 97116 75100 97180 75104
rect 97116 75044 97120 75100
rect 97120 75044 97176 75100
rect 97176 75044 97180 75100
rect 97116 75040 97180 75044
rect 97196 75100 97260 75104
rect 97196 75044 97200 75100
rect 97200 75044 97256 75100
rect 97256 75044 97260 75100
rect 97196 75040 97260 75044
rect 97276 75100 97340 75104
rect 97276 75044 97280 75100
rect 97280 75044 97336 75100
rect 97336 75044 97340 75100
rect 97276 75040 97340 75044
rect 4216 74556 4280 74560
rect 4216 74500 4220 74556
rect 4220 74500 4276 74556
rect 4276 74500 4280 74556
rect 4216 74496 4280 74500
rect 4296 74556 4360 74560
rect 4296 74500 4300 74556
rect 4300 74500 4356 74556
rect 4356 74500 4360 74556
rect 4296 74496 4360 74500
rect 4376 74556 4440 74560
rect 4376 74500 4380 74556
rect 4380 74500 4436 74556
rect 4436 74500 4440 74556
rect 4376 74496 4440 74500
rect 4456 74556 4520 74560
rect 4456 74500 4460 74556
rect 4460 74500 4516 74556
rect 4516 74500 4520 74556
rect 4456 74496 4520 74500
rect 34936 74556 35000 74560
rect 34936 74500 34940 74556
rect 34940 74500 34996 74556
rect 34996 74500 35000 74556
rect 34936 74496 35000 74500
rect 35016 74556 35080 74560
rect 35016 74500 35020 74556
rect 35020 74500 35076 74556
rect 35076 74500 35080 74556
rect 35016 74496 35080 74500
rect 35096 74556 35160 74560
rect 35096 74500 35100 74556
rect 35100 74500 35156 74556
rect 35156 74500 35160 74556
rect 35096 74496 35160 74500
rect 35176 74556 35240 74560
rect 35176 74500 35180 74556
rect 35180 74500 35236 74556
rect 35236 74500 35240 74556
rect 35176 74496 35240 74500
rect 65656 74556 65720 74560
rect 65656 74500 65660 74556
rect 65660 74500 65716 74556
rect 65716 74500 65720 74556
rect 65656 74496 65720 74500
rect 65736 74556 65800 74560
rect 65736 74500 65740 74556
rect 65740 74500 65796 74556
rect 65796 74500 65800 74556
rect 65736 74496 65800 74500
rect 65816 74556 65880 74560
rect 65816 74500 65820 74556
rect 65820 74500 65876 74556
rect 65876 74500 65880 74556
rect 65816 74496 65880 74500
rect 65896 74556 65960 74560
rect 65896 74500 65900 74556
rect 65900 74500 65956 74556
rect 65956 74500 65960 74556
rect 65896 74496 65960 74500
rect 96376 74556 96440 74560
rect 96376 74500 96380 74556
rect 96380 74500 96436 74556
rect 96436 74500 96440 74556
rect 96376 74496 96440 74500
rect 96456 74556 96520 74560
rect 96456 74500 96460 74556
rect 96460 74500 96516 74556
rect 96516 74500 96520 74556
rect 96456 74496 96520 74500
rect 96536 74556 96600 74560
rect 96536 74500 96540 74556
rect 96540 74500 96596 74556
rect 96596 74500 96600 74556
rect 96536 74496 96600 74500
rect 96616 74556 96680 74560
rect 96616 74500 96620 74556
rect 96620 74500 96676 74556
rect 96676 74500 96680 74556
rect 96616 74496 96680 74500
rect 4876 74012 4940 74016
rect 4876 73956 4880 74012
rect 4880 73956 4936 74012
rect 4936 73956 4940 74012
rect 4876 73952 4940 73956
rect 4956 74012 5020 74016
rect 4956 73956 4960 74012
rect 4960 73956 5016 74012
rect 5016 73956 5020 74012
rect 4956 73952 5020 73956
rect 5036 74012 5100 74016
rect 5036 73956 5040 74012
rect 5040 73956 5096 74012
rect 5096 73956 5100 74012
rect 5036 73952 5100 73956
rect 5116 74012 5180 74016
rect 5116 73956 5120 74012
rect 5120 73956 5176 74012
rect 5176 73956 5180 74012
rect 5116 73952 5180 73956
rect 35596 74012 35660 74016
rect 35596 73956 35600 74012
rect 35600 73956 35656 74012
rect 35656 73956 35660 74012
rect 35596 73952 35660 73956
rect 35676 74012 35740 74016
rect 35676 73956 35680 74012
rect 35680 73956 35736 74012
rect 35736 73956 35740 74012
rect 35676 73952 35740 73956
rect 35756 74012 35820 74016
rect 35756 73956 35760 74012
rect 35760 73956 35816 74012
rect 35816 73956 35820 74012
rect 35756 73952 35820 73956
rect 35836 74012 35900 74016
rect 35836 73956 35840 74012
rect 35840 73956 35896 74012
rect 35896 73956 35900 74012
rect 35836 73952 35900 73956
rect 66316 74012 66380 74016
rect 66316 73956 66320 74012
rect 66320 73956 66376 74012
rect 66376 73956 66380 74012
rect 66316 73952 66380 73956
rect 66396 74012 66460 74016
rect 66396 73956 66400 74012
rect 66400 73956 66456 74012
rect 66456 73956 66460 74012
rect 66396 73952 66460 73956
rect 66476 74012 66540 74016
rect 66476 73956 66480 74012
rect 66480 73956 66536 74012
rect 66536 73956 66540 74012
rect 66476 73952 66540 73956
rect 66556 74012 66620 74016
rect 66556 73956 66560 74012
rect 66560 73956 66616 74012
rect 66616 73956 66620 74012
rect 66556 73952 66620 73956
rect 97036 74012 97100 74016
rect 97036 73956 97040 74012
rect 97040 73956 97096 74012
rect 97096 73956 97100 74012
rect 97036 73952 97100 73956
rect 97116 74012 97180 74016
rect 97116 73956 97120 74012
rect 97120 73956 97176 74012
rect 97176 73956 97180 74012
rect 97116 73952 97180 73956
rect 97196 74012 97260 74016
rect 97196 73956 97200 74012
rect 97200 73956 97256 74012
rect 97256 73956 97260 74012
rect 97196 73952 97260 73956
rect 97276 74012 97340 74016
rect 97276 73956 97280 74012
rect 97280 73956 97336 74012
rect 97336 73956 97340 74012
rect 97276 73952 97340 73956
rect 4216 73468 4280 73472
rect 4216 73412 4220 73468
rect 4220 73412 4276 73468
rect 4276 73412 4280 73468
rect 4216 73408 4280 73412
rect 4296 73468 4360 73472
rect 4296 73412 4300 73468
rect 4300 73412 4356 73468
rect 4356 73412 4360 73468
rect 4296 73408 4360 73412
rect 4376 73468 4440 73472
rect 4376 73412 4380 73468
rect 4380 73412 4436 73468
rect 4436 73412 4440 73468
rect 4376 73408 4440 73412
rect 4456 73468 4520 73472
rect 4456 73412 4460 73468
rect 4460 73412 4516 73468
rect 4516 73412 4520 73468
rect 4456 73408 4520 73412
rect 34936 73468 35000 73472
rect 34936 73412 34940 73468
rect 34940 73412 34996 73468
rect 34996 73412 35000 73468
rect 34936 73408 35000 73412
rect 35016 73468 35080 73472
rect 35016 73412 35020 73468
rect 35020 73412 35076 73468
rect 35076 73412 35080 73468
rect 35016 73408 35080 73412
rect 35096 73468 35160 73472
rect 35096 73412 35100 73468
rect 35100 73412 35156 73468
rect 35156 73412 35160 73468
rect 35096 73408 35160 73412
rect 35176 73468 35240 73472
rect 35176 73412 35180 73468
rect 35180 73412 35236 73468
rect 35236 73412 35240 73468
rect 35176 73408 35240 73412
rect 65656 73468 65720 73472
rect 65656 73412 65660 73468
rect 65660 73412 65716 73468
rect 65716 73412 65720 73468
rect 65656 73408 65720 73412
rect 65736 73468 65800 73472
rect 65736 73412 65740 73468
rect 65740 73412 65796 73468
rect 65796 73412 65800 73468
rect 65736 73408 65800 73412
rect 65816 73468 65880 73472
rect 65816 73412 65820 73468
rect 65820 73412 65876 73468
rect 65876 73412 65880 73468
rect 65816 73408 65880 73412
rect 65896 73468 65960 73472
rect 65896 73412 65900 73468
rect 65900 73412 65956 73468
rect 65956 73412 65960 73468
rect 65896 73408 65960 73412
rect 96376 73468 96440 73472
rect 96376 73412 96380 73468
rect 96380 73412 96436 73468
rect 96436 73412 96440 73468
rect 96376 73408 96440 73412
rect 96456 73468 96520 73472
rect 96456 73412 96460 73468
rect 96460 73412 96516 73468
rect 96516 73412 96520 73468
rect 96456 73408 96520 73412
rect 96536 73468 96600 73472
rect 96536 73412 96540 73468
rect 96540 73412 96596 73468
rect 96596 73412 96600 73468
rect 96536 73408 96600 73412
rect 96616 73468 96680 73472
rect 96616 73412 96620 73468
rect 96620 73412 96676 73468
rect 96676 73412 96680 73468
rect 96616 73408 96680 73412
rect 4876 72924 4940 72928
rect 4876 72868 4880 72924
rect 4880 72868 4936 72924
rect 4936 72868 4940 72924
rect 4876 72864 4940 72868
rect 4956 72924 5020 72928
rect 4956 72868 4960 72924
rect 4960 72868 5016 72924
rect 5016 72868 5020 72924
rect 4956 72864 5020 72868
rect 5036 72924 5100 72928
rect 5036 72868 5040 72924
rect 5040 72868 5096 72924
rect 5096 72868 5100 72924
rect 5036 72864 5100 72868
rect 5116 72924 5180 72928
rect 5116 72868 5120 72924
rect 5120 72868 5176 72924
rect 5176 72868 5180 72924
rect 5116 72864 5180 72868
rect 35596 72924 35660 72928
rect 35596 72868 35600 72924
rect 35600 72868 35656 72924
rect 35656 72868 35660 72924
rect 35596 72864 35660 72868
rect 35676 72924 35740 72928
rect 35676 72868 35680 72924
rect 35680 72868 35736 72924
rect 35736 72868 35740 72924
rect 35676 72864 35740 72868
rect 35756 72924 35820 72928
rect 35756 72868 35760 72924
rect 35760 72868 35816 72924
rect 35816 72868 35820 72924
rect 35756 72864 35820 72868
rect 35836 72924 35900 72928
rect 35836 72868 35840 72924
rect 35840 72868 35896 72924
rect 35896 72868 35900 72924
rect 35836 72864 35900 72868
rect 66316 72924 66380 72928
rect 66316 72868 66320 72924
rect 66320 72868 66376 72924
rect 66376 72868 66380 72924
rect 66316 72864 66380 72868
rect 66396 72924 66460 72928
rect 66396 72868 66400 72924
rect 66400 72868 66456 72924
rect 66456 72868 66460 72924
rect 66396 72864 66460 72868
rect 66476 72924 66540 72928
rect 66476 72868 66480 72924
rect 66480 72868 66536 72924
rect 66536 72868 66540 72924
rect 66476 72864 66540 72868
rect 66556 72924 66620 72928
rect 66556 72868 66560 72924
rect 66560 72868 66616 72924
rect 66616 72868 66620 72924
rect 66556 72864 66620 72868
rect 97036 72924 97100 72928
rect 97036 72868 97040 72924
rect 97040 72868 97096 72924
rect 97096 72868 97100 72924
rect 97036 72864 97100 72868
rect 97116 72924 97180 72928
rect 97116 72868 97120 72924
rect 97120 72868 97176 72924
rect 97176 72868 97180 72924
rect 97116 72864 97180 72868
rect 97196 72924 97260 72928
rect 97196 72868 97200 72924
rect 97200 72868 97256 72924
rect 97256 72868 97260 72924
rect 97196 72864 97260 72868
rect 97276 72924 97340 72928
rect 97276 72868 97280 72924
rect 97280 72868 97336 72924
rect 97336 72868 97340 72924
rect 97276 72864 97340 72868
rect 4216 72380 4280 72384
rect 4216 72324 4220 72380
rect 4220 72324 4276 72380
rect 4276 72324 4280 72380
rect 4216 72320 4280 72324
rect 4296 72380 4360 72384
rect 4296 72324 4300 72380
rect 4300 72324 4356 72380
rect 4356 72324 4360 72380
rect 4296 72320 4360 72324
rect 4376 72380 4440 72384
rect 4376 72324 4380 72380
rect 4380 72324 4436 72380
rect 4436 72324 4440 72380
rect 4376 72320 4440 72324
rect 4456 72380 4520 72384
rect 4456 72324 4460 72380
rect 4460 72324 4516 72380
rect 4516 72324 4520 72380
rect 4456 72320 4520 72324
rect 34936 72380 35000 72384
rect 34936 72324 34940 72380
rect 34940 72324 34996 72380
rect 34996 72324 35000 72380
rect 34936 72320 35000 72324
rect 35016 72380 35080 72384
rect 35016 72324 35020 72380
rect 35020 72324 35076 72380
rect 35076 72324 35080 72380
rect 35016 72320 35080 72324
rect 35096 72380 35160 72384
rect 35096 72324 35100 72380
rect 35100 72324 35156 72380
rect 35156 72324 35160 72380
rect 35096 72320 35160 72324
rect 35176 72380 35240 72384
rect 35176 72324 35180 72380
rect 35180 72324 35236 72380
rect 35236 72324 35240 72380
rect 35176 72320 35240 72324
rect 65656 72380 65720 72384
rect 65656 72324 65660 72380
rect 65660 72324 65716 72380
rect 65716 72324 65720 72380
rect 65656 72320 65720 72324
rect 65736 72380 65800 72384
rect 65736 72324 65740 72380
rect 65740 72324 65796 72380
rect 65796 72324 65800 72380
rect 65736 72320 65800 72324
rect 65816 72380 65880 72384
rect 65816 72324 65820 72380
rect 65820 72324 65876 72380
rect 65876 72324 65880 72380
rect 65816 72320 65880 72324
rect 65896 72380 65960 72384
rect 65896 72324 65900 72380
rect 65900 72324 65956 72380
rect 65956 72324 65960 72380
rect 65896 72320 65960 72324
rect 96376 72380 96440 72384
rect 96376 72324 96380 72380
rect 96380 72324 96436 72380
rect 96436 72324 96440 72380
rect 96376 72320 96440 72324
rect 96456 72380 96520 72384
rect 96456 72324 96460 72380
rect 96460 72324 96516 72380
rect 96516 72324 96520 72380
rect 96456 72320 96520 72324
rect 96536 72380 96600 72384
rect 96536 72324 96540 72380
rect 96540 72324 96596 72380
rect 96596 72324 96600 72380
rect 96536 72320 96600 72324
rect 96616 72380 96680 72384
rect 96616 72324 96620 72380
rect 96620 72324 96676 72380
rect 96676 72324 96680 72380
rect 96616 72320 96680 72324
rect 4876 71836 4940 71840
rect 4876 71780 4880 71836
rect 4880 71780 4936 71836
rect 4936 71780 4940 71836
rect 4876 71776 4940 71780
rect 4956 71836 5020 71840
rect 4956 71780 4960 71836
rect 4960 71780 5016 71836
rect 5016 71780 5020 71836
rect 4956 71776 5020 71780
rect 5036 71836 5100 71840
rect 5036 71780 5040 71836
rect 5040 71780 5096 71836
rect 5096 71780 5100 71836
rect 5036 71776 5100 71780
rect 5116 71836 5180 71840
rect 5116 71780 5120 71836
rect 5120 71780 5176 71836
rect 5176 71780 5180 71836
rect 5116 71776 5180 71780
rect 35596 71836 35660 71840
rect 35596 71780 35600 71836
rect 35600 71780 35656 71836
rect 35656 71780 35660 71836
rect 35596 71776 35660 71780
rect 35676 71836 35740 71840
rect 35676 71780 35680 71836
rect 35680 71780 35736 71836
rect 35736 71780 35740 71836
rect 35676 71776 35740 71780
rect 35756 71836 35820 71840
rect 35756 71780 35760 71836
rect 35760 71780 35816 71836
rect 35816 71780 35820 71836
rect 35756 71776 35820 71780
rect 35836 71836 35900 71840
rect 35836 71780 35840 71836
rect 35840 71780 35896 71836
rect 35896 71780 35900 71836
rect 35836 71776 35900 71780
rect 66316 71836 66380 71840
rect 66316 71780 66320 71836
rect 66320 71780 66376 71836
rect 66376 71780 66380 71836
rect 66316 71776 66380 71780
rect 66396 71836 66460 71840
rect 66396 71780 66400 71836
rect 66400 71780 66456 71836
rect 66456 71780 66460 71836
rect 66396 71776 66460 71780
rect 66476 71836 66540 71840
rect 66476 71780 66480 71836
rect 66480 71780 66536 71836
rect 66536 71780 66540 71836
rect 66476 71776 66540 71780
rect 66556 71836 66620 71840
rect 66556 71780 66560 71836
rect 66560 71780 66616 71836
rect 66616 71780 66620 71836
rect 66556 71776 66620 71780
rect 97036 71836 97100 71840
rect 97036 71780 97040 71836
rect 97040 71780 97096 71836
rect 97096 71780 97100 71836
rect 97036 71776 97100 71780
rect 97116 71836 97180 71840
rect 97116 71780 97120 71836
rect 97120 71780 97176 71836
rect 97176 71780 97180 71836
rect 97116 71776 97180 71780
rect 97196 71836 97260 71840
rect 97196 71780 97200 71836
rect 97200 71780 97256 71836
rect 97256 71780 97260 71836
rect 97196 71776 97260 71780
rect 97276 71836 97340 71840
rect 97276 71780 97280 71836
rect 97280 71780 97336 71836
rect 97336 71780 97340 71836
rect 97276 71776 97340 71780
rect 4216 71292 4280 71296
rect 4216 71236 4220 71292
rect 4220 71236 4276 71292
rect 4276 71236 4280 71292
rect 4216 71232 4280 71236
rect 4296 71292 4360 71296
rect 4296 71236 4300 71292
rect 4300 71236 4356 71292
rect 4356 71236 4360 71292
rect 4296 71232 4360 71236
rect 4376 71292 4440 71296
rect 4376 71236 4380 71292
rect 4380 71236 4436 71292
rect 4436 71236 4440 71292
rect 4376 71232 4440 71236
rect 4456 71292 4520 71296
rect 4456 71236 4460 71292
rect 4460 71236 4516 71292
rect 4516 71236 4520 71292
rect 4456 71232 4520 71236
rect 34936 71292 35000 71296
rect 34936 71236 34940 71292
rect 34940 71236 34996 71292
rect 34996 71236 35000 71292
rect 34936 71232 35000 71236
rect 35016 71292 35080 71296
rect 35016 71236 35020 71292
rect 35020 71236 35076 71292
rect 35076 71236 35080 71292
rect 35016 71232 35080 71236
rect 35096 71292 35160 71296
rect 35096 71236 35100 71292
rect 35100 71236 35156 71292
rect 35156 71236 35160 71292
rect 35096 71232 35160 71236
rect 35176 71292 35240 71296
rect 35176 71236 35180 71292
rect 35180 71236 35236 71292
rect 35236 71236 35240 71292
rect 35176 71232 35240 71236
rect 65656 71292 65720 71296
rect 65656 71236 65660 71292
rect 65660 71236 65716 71292
rect 65716 71236 65720 71292
rect 65656 71232 65720 71236
rect 65736 71292 65800 71296
rect 65736 71236 65740 71292
rect 65740 71236 65796 71292
rect 65796 71236 65800 71292
rect 65736 71232 65800 71236
rect 65816 71292 65880 71296
rect 65816 71236 65820 71292
rect 65820 71236 65876 71292
rect 65876 71236 65880 71292
rect 65816 71232 65880 71236
rect 65896 71292 65960 71296
rect 65896 71236 65900 71292
rect 65900 71236 65956 71292
rect 65956 71236 65960 71292
rect 65896 71232 65960 71236
rect 96376 71292 96440 71296
rect 96376 71236 96380 71292
rect 96380 71236 96436 71292
rect 96436 71236 96440 71292
rect 96376 71232 96440 71236
rect 96456 71292 96520 71296
rect 96456 71236 96460 71292
rect 96460 71236 96516 71292
rect 96516 71236 96520 71292
rect 96456 71232 96520 71236
rect 96536 71292 96600 71296
rect 96536 71236 96540 71292
rect 96540 71236 96596 71292
rect 96596 71236 96600 71292
rect 96536 71232 96600 71236
rect 96616 71292 96680 71296
rect 96616 71236 96620 71292
rect 96620 71236 96676 71292
rect 96676 71236 96680 71292
rect 96616 71232 96680 71236
rect 4876 70748 4940 70752
rect 4876 70692 4880 70748
rect 4880 70692 4936 70748
rect 4936 70692 4940 70748
rect 4876 70688 4940 70692
rect 4956 70748 5020 70752
rect 4956 70692 4960 70748
rect 4960 70692 5016 70748
rect 5016 70692 5020 70748
rect 4956 70688 5020 70692
rect 5036 70748 5100 70752
rect 5036 70692 5040 70748
rect 5040 70692 5096 70748
rect 5096 70692 5100 70748
rect 5036 70688 5100 70692
rect 5116 70748 5180 70752
rect 5116 70692 5120 70748
rect 5120 70692 5176 70748
rect 5176 70692 5180 70748
rect 5116 70688 5180 70692
rect 35596 70748 35660 70752
rect 35596 70692 35600 70748
rect 35600 70692 35656 70748
rect 35656 70692 35660 70748
rect 35596 70688 35660 70692
rect 35676 70748 35740 70752
rect 35676 70692 35680 70748
rect 35680 70692 35736 70748
rect 35736 70692 35740 70748
rect 35676 70688 35740 70692
rect 35756 70748 35820 70752
rect 35756 70692 35760 70748
rect 35760 70692 35816 70748
rect 35816 70692 35820 70748
rect 35756 70688 35820 70692
rect 35836 70748 35900 70752
rect 35836 70692 35840 70748
rect 35840 70692 35896 70748
rect 35896 70692 35900 70748
rect 35836 70688 35900 70692
rect 66316 70748 66380 70752
rect 66316 70692 66320 70748
rect 66320 70692 66376 70748
rect 66376 70692 66380 70748
rect 66316 70688 66380 70692
rect 66396 70748 66460 70752
rect 66396 70692 66400 70748
rect 66400 70692 66456 70748
rect 66456 70692 66460 70748
rect 66396 70688 66460 70692
rect 66476 70748 66540 70752
rect 66476 70692 66480 70748
rect 66480 70692 66536 70748
rect 66536 70692 66540 70748
rect 66476 70688 66540 70692
rect 66556 70748 66620 70752
rect 66556 70692 66560 70748
rect 66560 70692 66616 70748
rect 66616 70692 66620 70748
rect 66556 70688 66620 70692
rect 97036 70748 97100 70752
rect 97036 70692 97040 70748
rect 97040 70692 97096 70748
rect 97096 70692 97100 70748
rect 97036 70688 97100 70692
rect 97116 70748 97180 70752
rect 97116 70692 97120 70748
rect 97120 70692 97176 70748
rect 97176 70692 97180 70748
rect 97116 70688 97180 70692
rect 97196 70748 97260 70752
rect 97196 70692 97200 70748
rect 97200 70692 97256 70748
rect 97256 70692 97260 70748
rect 97196 70688 97260 70692
rect 97276 70748 97340 70752
rect 97276 70692 97280 70748
rect 97280 70692 97336 70748
rect 97336 70692 97340 70748
rect 97276 70688 97340 70692
rect 4216 70204 4280 70208
rect 4216 70148 4220 70204
rect 4220 70148 4276 70204
rect 4276 70148 4280 70204
rect 4216 70144 4280 70148
rect 4296 70204 4360 70208
rect 4296 70148 4300 70204
rect 4300 70148 4356 70204
rect 4356 70148 4360 70204
rect 4296 70144 4360 70148
rect 4376 70204 4440 70208
rect 4376 70148 4380 70204
rect 4380 70148 4436 70204
rect 4436 70148 4440 70204
rect 4376 70144 4440 70148
rect 4456 70204 4520 70208
rect 4456 70148 4460 70204
rect 4460 70148 4516 70204
rect 4516 70148 4520 70204
rect 4456 70144 4520 70148
rect 34936 70204 35000 70208
rect 34936 70148 34940 70204
rect 34940 70148 34996 70204
rect 34996 70148 35000 70204
rect 34936 70144 35000 70148
rect 35016 70204 35080 70208
rect 35016 70148 35020 70204
rect 35020 70148 35076 70204
rect 35076 70148 35080 70204
rect 35016 70144 35080 70148
rect 35096 70204 35160 70208
rect 35096 70148 35100 70204
rect 35100 70148 35156 70204
rect 35156 70148 35160 70204
rect 35096 70144 35160 70148
rect 35176 70204 35240 70208
rect 35176 70148 35180 70204
rect 35180 70148 35236 70204
rect 35236 70148 35240 70204
rect 35176 70144 35240 70148
rect 65656 70204 65720 70208
rect 65656 70148 65660 70204
rect 65660 70148 65716 70204
rect 65716 70148 65720 70204
rect 65656 70144 65720 70148
rect 65736 70204 65800 70208
rect 65736 70148 65740 70204
rect 65740 70148 65796 70204
rect 65796 70148 65800 70204
rect 65736 70144 65800 70148
rect 65816 70204 65880 70208
rect 65816 70148 65820 70204
rect 65820 70148 65876 70204
rect 65876 70148 65880 70204
rect 65816 70144 65880 70148
rect 65896 70204 65960 70208
rect 65896 70148 65900 70204
rect 65900 70148 65956 70204
rect 65956 70148 65960 70204
rect 65896 70144 65960 70148
rect 96376 70204 96440 70208
rect 96376 70148 96380 70204
rect 96380 70148 96436 70204
rect 96436 70148 96440 70204
rect 96376 70144 96440 70148
rect 96456 70204 96520 70208
rect 96456 70148 96460 70204
rect 96460 70148 96516 70204
rect 96516 70148 96520 70204
rect 96456 70144 96520 70148
rect 96536 70204 96600 70208
rect 96536 70148 96540 70204
rect 96540 70148 96596 70204
rect 96596 70148 96600 70204
rect 96536 70144 96600 70148
rect 96616 70204 96680 70208
rect 96616 70148 96620 70204
rect 96620 70148 96676 70204
rect 96676 70148 96680 70204
rect 96616 70144 96680 70148
rect 4876 69660 4940 69664
rect 4876 69604 4880 69660
rect 4880 69604 4936 69660
rect 4936 69604 4940 69660
rect 4876 69600 4940 69604
rect 4956 69660 5020 69664
rect 4956 69604 4960 69660
rect 4960 69604 5016 69660
rect 5016 69604 5020 69660
rect 4956 69600 5020 69604
rect 5036 69660 5100 69664
rect 5036 69604 5040 69660
rect 5040 69604 5096 69660
rect 5096 69604 5100 69660
rect 5036 69600 5100 69604
rect 5116 69660 5180 69664
rect 5116 69604 5120 69660
rect 5120 69604 5176 69660
rect 5176 69604 5180 69660
rect 5116 69600 5180 69604
rect 35596 69660 35660 69664
rect 35596 69604 35600 69660
rect 35600 69604 35656 69660
rect 35656 69604 35660 69660
rect 35596 69600 35660 69604
rect 35676 69660 35740 69664
rect 35676 69604 35680 69660
rect 35680 69604 35736 69660
rect 35736 69604 35740 69660
rect 35676 69600 35740 69604
rect 35756 69660 35820 69664
rect 35756 69604 35760 69660
rect 35760 69604 35816 69660
rect 35816 69604 35820 69660
rect 35756 69600 35820 69604
rect 35836 69660 35900 69664
rect 35836 69604 35840 69660
rect 35840 69604 35896 69660
rect 35896 69604 35900 69660
rect 35836 69600 35900 69604
rect 66316 69660 66380 69664
rect 66316 69604 66320 69660
rect 66320 69604 66376 69660
rect 66376 69604 66380 69660
rect 66316 69600 66380 69604
rect 66396 69660 66460 69664
rect 66396 69604 66400 69660
rect 66400 69604 66456 69660
rect 66456 69604 66460 69660
rect 66396 69600 66460 69604
rect 66476 69660 66540 69664
rect 66476 69604 66480 69660
rect 66480 69604 66536 69660
rect 66536 69604 66540 69660
rect 66476 69600 66540 69604
rect 66556 69660 66620 69664
rect 66556 69604 66560 69660
rect 66560 69604 66616 69660
rect 66616 69604 66620 69660
rect 66556 69600 66620 69604
rect 97036 69660 97100 69664
rect 97036 69604 97040 69660
rect 97040 69604 97096 69660
rect 97096 69604 97100 69660
rect 97036 69600 97100 69604
rect 97116 69660 97180 69664
rect 97116 69604 97120 69660
rect 97120 69604 97176 69660
rect 97176 69604 97180 69660
rect 97116 69600 97180 69604
rect 97196 69660 97260 69664
rect 97196 69604 97200 69660
rect 97200 69604 97256 69660
rect 97256 69604 97260 69660
rect 97196 69600 97260 69604
rect 97276 69660 97340 69664
rect 97276 69604 97280 69660
rect 97280 69604 97336 69660
rect 97336 69604 97340 69660
rect 97276 69600 97340 69604
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 34936 69116 35000 69120
rect 34936 69060 34940 69116
rect 34940 69060 34996 69116
rect 34996 69060 35000 69116
rect 34936 69056 35000 69060
rect 35016 69116 35080 69120
rect 35016 69060 35020 69116
rect 35020 69060 35076 69116
rect 35076 69060 35080 69116
rect 35016 69056 35080 69060
rect 35096 69116 35160 69120
rect 35096 69060 35100 69116
rect 35100 69060 35156 69116
rect 35156 69060 35160 69116
rect 35096 69056 35160 69060
rect 35176 69116 35240 69120
rect 35176 69060 35180 69116
rect 35180 69060 35236 69116
rect 35236 69060 35240 69116
rect 35176 69056 35240 69060
rect 65656 69116 65720 69120
rect 65656 69060 65660 69116
rect 65660 69060 65716 69116
rect 65716 69060 65720 69116
rect 65656 69056 65720 69060
rect 65736 69116 65800 69120
rect 65736 69060 65740 69116
rect 65740 69060 65796 69116
rect 65796 69060 65800 69116
rect 65736 69056 65800 69060
rect 65816 69116 65880 69120
rect 65816 69060 65820 69116
rect 65820 69060 65876 69116
rect 65876 69060 65880 69116
rect 65816 69056 65880 69060
rect 65896 69116 65960 69120
rect 65896 69060 65900 69116
rect 65900 69060 65956 69116
rect 65956 69060 65960 69116
rect 65896 69056 65960 69060
rect 96376 69116 96440 69120
rect 96376 69060 96380 69116
rect 96380 69060 96436 69116
rect 96436 69060 96440 69116
rect 96376 69056 96440 69060
rect 96456 69116 96520 69120
rect 96456 69060 96460 69116
rect 96460 69060 96516 69116
rect 96516 69060 96520 69116
rect 96456 69056 96520 69060
rect 96536 69116 96600 69120
rect 96536 69060 96540 69116
rect 96540 69060 96596 69116
rect 96596 69060 96600 69116
rect 96536 69056 96600 69060
rect 96616 69116 96680 69120
rect 96616 69060 96620 69116
rect 96620 69060 96676 69116
rect 96676 69060 96680 69116
rect 96616 69056 96680 69060
rect 87276 68988 87340 69052
rect 4876 68572 4940 68576
rect 4876 68516 4880 68572
rect 4880 68516 4936 68572
rect 4936 68516 4940 68572
rect 4876 68512 4940 68516
rect 4956 68572 5020 68576
rect 4956 68516 4960 68572
rect 4960 68516 5016 68572
rect 5016 68516 5020 68572
rect 4956 68512 5020 68516
rect 5036 68572 5100 68576
rect 5036 68516 5040 68572
rect 5040 68516 5096 68572
rect 5096 68516 5100 68572
rect 5036 68512 5100 68516
rect 5116 68572 5180 68576
rect 5116 68516 5120 68572
rect 5120 68516 5176 68572
rect 5176 68516 5180 68572
rect 5116 68512 5180 68516
rect 35596 68572 35660 68576
rect 35596 68516 35600 68572
rect 35600 68516 35656 68572
rect 35656 68516 35660 68572
rect 35596 68512 35660 68516
rect 35676 68572 35740 68576
rect 35676 68516 35680 68572
rect 35680 68516 35736 68572
rect 35736 68516 35740 68572
rect 35676 68512 35740 68516
rect 35756 68572 35820 68576
rect 35756 68516 35760 68572
rect 35760 68516 35816 68572
rect 35816 68516 35820 68572
rect 35756 68512 35820 68516
rect 35836 68572 35900 68576
rect 35836 68516 35840 68572
rect 35840 68516 35896 68572
rect 35896 68516 35900 68572
rect 35836 68512 35900 68516
rect 66316 68572 66380 68576
rect 66316 68516 66320 68572
rect 66320 68516 66376 68572
rect 66376 68516 66380 68572
rect 66316 68512 66380 68516
rect 66396 68572 66460 68576
rect 66396 68516 66400 68572
rect 66400 68516 66456 68572
rect 66456 68516 66460 68572
rect 66396 68512 66460 68516
rect 66476 68572 66540 68576
rect 66476 68516 66480 68572
rect 66480 68516 66536 68572
rect 66536 68516 66540 68572
rect 66476 68512 66540 68516
rect 66556 68572 66620 68576
rect 66556 68516 66560 68572
rect 66560 68516 66616 68572
rect 66616 68516 66620 68572
rect 66556 68512 66620 68516
rect 97036 68572 97100 68576
rect 97036 68516 97040 68572
rect 97040 68516 97096 68572
rect 97096 68516 97100 68572
rect 97036 68512 97100 68516
rect 97116 68572 97180 68576
rect 97116 68516 97120 68572
rect 97120 68516 97176 68572
rect 97176 68516 97180 68572
rect 97116 68512 97180 68516
rect 97196 68572 97260 68576
rect 97196 68516 97200 68572
rect 97200 68516 97256 68572
rect 97256 68516 97260 68572
rect 97196 68512 97260 68516
rect 97276 68572 97340 68576
rect 97276 68516 97280 68572
rect 97280 68516 97336 68572
rect 97336 68516 97340 68572
rect 97276 68512 97340 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 34936 68028 35000 68032
rect 34936 67972 34940 68028
rect 34940 67972 34996 68028
rect 34996 67972 35000 68028
rect 34936 67968 35000 67972
rect 35016 68028 35080 68032
rect 35016 67972 35020 68028
rect 35020 67972 35076 68028
rect 35076 67972 35080 68028
rect 35016 67968 35080 67972
rect 35096 68028 35160 68032
rect 35096 67972 35100 68028
rect 35100 67972 35156 68028
rect 35156 67972 35160 68028
rect 35096 67968 35160 67972
rect 35176 68028 35240 68032
rect 35176 67972 35180 68028
rect 35180 67972 35236 68028
rect 35236 67972 35240 68028
rect 35176 67968 35240 67972
rect 65656 68028 65720 68032
rect 65656 67972 65660 68028
rect 65660 67972 65716 68028
rect 65716 67972 65720 68028
rect 65656 67968 65720 67972
rect 65736 68028 65800 68032
rect 65736 67972 65740 68028
rect 65740 67972 65796 68028
rect 65796 67972 65800 68028
rect 65736 67968 65800 67972
rect 65816 68028 65880 68032
rect 65816 67972 65820 68028
rect 65820 67972 65876 68028
rect 65876 67972 65880 68028
rect 65816 67968 65880 67972
rect 65896 68028 65960 68032
rect 65896 67972 65900 68028
rect 65900 67972 65956 68028
rect 65956 67972 65960 68028
rect 65896 67968 65960 67972
rect 96376 68028 96440 68032
rect 96376 67972 96380 68028
rect 96380 67972 96436 68028
rect 96436 67972 96440 68028
rect 96376 67968 96440 67972
rect 96456 68028 96520 68032
rect 96456 67972 96460 68028
rect 96460 67972 96516 68028
rect 96516 67972 96520 68028
rect 96456 67968 96520 67972
rect 96536 68028 96600 68032
rect 96536 67972 96540 68028
rect 96540 67972 96596 68028
rect 96596 67972 96600 68028
rect 96536 67968 96600 67972
rect 96616 68028 96680 68032
rect 96616 67972 96620 68028
rect 96620 67972 96676 68028
rect 96676 67972 96680 68028
rect 96616 67968 96680 67972
rect 4876 67484 4940 67488
rect 4876 67428 4880 67484
rect 4880 67428 4936 67484
rect 4936 67428 4940 67484
rect 4876 67424 4940 67428
rect 4956 67484 5020 67488
rect 4956 67428 4960 67484
rect 4960 67428 5016 67484
rect 5016 67428 5020 67484
rect 4956 67424 5020 67428
rect 5036 67484 5100 67488
rect 5036 67428 5040 67484
rect 5040 67428 5096 67484
rect 5096 67428 5100 67484
rect 5036 67424 5100 67428
rect 5116 67484 5180 67488
rect 5116 67428 5120 67484
rect 5120 67428 5176 67484
rect 5176 67428 5180 67484
rect 5116 67424 5180 67428
rect 35596 67484 35660 67488
rect 35596 67428 35600 67484
rect 35600 67428 35656 67484
rect 35656 67428 35660 67484
rect 35596 67424 35660 67428
rect 35676 67484 35740 67488
rect 35676 67428 35680 67484
rect 35680 67428 35736 67484
rect 35736 67428 35740 67484
rect 35676 67424 35740 67428
rect 35756 67484 35820 67488
rect 35756 67428 35760 67484
rect 35760 67428 35816 67484
rect 35816 67428 35820 67484
rect 35756 67424 35820 67428
rect 35836 67484 35900 67488
rect 35836 67428 35840 67484
rect 35840 67428 35896 67484
rect 35896 67428 35900 67484
rect 35836 67424 35900 67428
rect 66316 67484 66380 67488
rect 66316 67428 66320 67484
rect 66320 67428 66376 67484
rect 66376 67428 66380 67484
rect 66316 67424 66380 67428
rect 66396 67484 66460 67488
rect 66396 67428 66400 67484
rect 66400 67428 66456 67484
rect 66456 67428 66460 67484
rect 66396 67424 66460 67428
rect 66476 67484 66540 67488
rect 66476 67428 66480 67484
rect 66480 67428 66536 67484
rect 66536 67428 66540 67484
rect 66476 67424 66540 67428
rect 66556 67484 66620 67488
rect 66556 67428 66560 67484
rect 66560 67428 66616 67484
rect 66616 67428 66620 67484
rect 66556 67424 66620 67428
rect 97036 67484 97100 67488
rect 97036 67428 97040 67484
rect 97040 67428 97096 67484
rect 97096 67428 97100 67484
rect 97036 67424 97100 67428
rect 97116 67484 97180 67488
rect 97116 67428 97120 67484
rect 97120 67428 97176 67484
rect 97176 67428 97180 67484
rect 97116 67424 97180 67428
rect 97196 67484 97260 67488
rect 97196 67428 97200 67484
rect 97200 67428 97256 67484
rect 97256 67428 97260 67484
rect 97196 67424 97260 67428
rect 97276 67484 97340 67488
rect 97276 67428 97280 67484
rect 97280 67428 97336 67484
rect 97336 67428 97340 67484
rect 97276 67424 97340 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 96376 66940 96440 66944
rect 96376 66884 96380 66940
rect 96380 66884 96436 66940
rect 96436 66884 96440 66940
rect 96376 66880 96440 66884
rect 96456 66940 96520 66944
rect 96456 66884 96460 66940
rect 96460 66884 96516 66940
rect 96516 66884 96520 66940
rect 96456 66880 96520 66884
rect 96536 66940 96600 66944
rect 96536 66884 96540 66940
rect 96540 66884 96596 66940
rect 96596 66884 96600 66940
rect 96536 66880 96600 66884
rect 96616 66940 96680 66944
rect 96616 66884 96620 66940
rect 96620 66884 96676 66940
rect 96676 66884 96680 66940
rect 96616 66880 96680 66884
rect 4876 66396 4940 66400
rect 4876 66340 4880 66396
rect 4880 66340 4936 66396
rect 4936 66340 4940 66396
rect 4876 66336 4940 66340
rect 4956 66396 5020 66400
rect 4956 66340 4960 66396
rect 4960 66340 5016 66396
rect 5016 66340 5020 66396
rect 4956 66336 5020 66340
rect 5036 66396 5100 66400
rect 5036 66340 5040 66396
rect 5040 66340 5096 66396
rect 5096 66340 5100 66396
rect 5036 66336 5100 66340
rect 5116 66396 5180 66400
rect 5116 66340 5120 66396
rect 5120 66340 5176 66396
rect 5176 66340 5180 66396
rect 5116 66336 5180 66340
rect 35596 66396 35660 66400
rect 35596 66340 35600 66396
rect 35600 66340 35656 66396
rect 35656 66340 35660 66396
rect 35596 66336 35660 66340
rect 35676 66396 35740 66400
rect 35676 66340 35680 66396
rect 35680 66340 35736 66396
rect 35736 66340 35740 66396
rect 35676 66336 35740 66340
rect 35756 66396 35820 66400
rect 35756 66340 35760 66396
rect 35760 66340 35816 66396
rect 35816 66340 35820 66396
rect 35756 66336 35820 66340
rect 35836 66396 35900 66400
rect 35836 66340 35840 66396
rect 35840 66340 35896 66396
rect 35896 66340 35900 66396
rect 35836 66336 35900 66340
rect 66316 66396 66380 66400
rect 66316 66340 66320 66396
rect 66320 66340 66376 66396
rect 66376 66340 66380 66396
rect 66316 66336 66380 66340
rect 66396 66396 66460 66400
rect 66396 66340 66400 66396
rect 66400 66340 66456 66396
rect 66456 66340 66460 66396
rect 66396 66336 66460 66340
rect 66476 66396 66540 66400
rect 66476 66340 66480 66396
rect 66480 66340 66536 66396
rect 66536 66340 66540 66396
rect 66476 66336 66540 66340
rect 66556 66396 66620 66400
rect 66556 66340 66560 66396
rect 66560 66340 66616 66396
rect 66616 66340 66620 66396
rect 66556 66336 66620 66340
rect 97036 66396 97100 66400
rect 97036 66340 97040 66396
rect 97040 66340 97096 66396
rect 97096 66340 97100 66396
rect 97036 66336 97100 66340
rect 97116 66396 97180 66400
rect 97116 66340 97120 66396
rect 97120 66340 97176 66396
rect 97176 66340 97180 66396
rect 97116 66336 97180 66340
rect 97196 66396 97260 66400
rect 97196 66340 97200 66396
rect 97200 66340 97256 66396
rect 97256 66340 97260 66396
rect 97196 66336 97260 66340
rect 97276 66396 97340 66400
rect 97276 66340 97280 66396
rect 97280 66340 97336 66396
rect 97336 66340 97340 66396
rect 97276 66336 97340 66340
rect 106660 66396 106724 66400
rect 106660 66340 106664 66396
rect 106664 66340 106720 66396
rect 106720 66340 106724 66396
rect 106660 66336 106724 66340
rect 106740 66396 106804 66400
rect 106740 66340 106744 66396
rect 106744 66340 106800 66396
rect 106800 66340 106804 66396
rect 106740 66336 106804 66340
rect 106820 66396 106884 66400
rect 106820 66340 106824 66396
rect 106824 66340 106880 66396
rect 106880 66340 106884 66396
rect 106820 66336 106884 66340
rect 106900 66396 106964 66400
rect 106900 66340 106904 66396
rect 106904 66340 106960 66396
rect 106960 66340 106964 66396
rect 106900 66336 106964 66340
rect 36124 66192 36188 66196
rect 36124 66136 36138 66192
rect 36138 66136 36188 66192
rect 36124 66132 36188 66136
rect 38516 66192 38580 66196
rect 38516 66136 38530 66192
rect 38530 66136 38580 66192
rect 38516 66132 38580 66136
rect 41092 66192 41156 66196
rect 41092 66136 41142 66192
rect 41142 66136 41156 66192
rect 41092 66132 41156 66136
rect 43668 66192 43732 66196
rect 43668 66136 43682 66192
rect 43682 66136 43732 66192
rect 43668 66132 43732 66136
rect 46060 66192 46124 66196
rect 46060 66136 46110 66192
rect 46110 66136 46124 66192
rect 46060 66132 46124 66136
rect 48636 66192 48700 66196
rect 48636 66136 48650 66192
rect 48650 66136 48700 66192
rect 48636 66132 48700 66136
rect 51028 66192 51092 66196
rect 51028 66136 51078 66192
rect 51078 66136 51092 66192
rect 51028 66132 51092 66136
rect 53604 66192 53668 66196
rect 53604 66136 53618 66192
rect 53618 66136 53668 66192
rect 53604 66132 53668 66136
rect 55996 66132 56060 66196
rect 58572 66192 58636 66196
rect 58572 66136 58622 66192
rect 58622 66136 58636 66192
rect 58572 66132 58636 66136
rect 61148 66192 61212 66196
rect 61148 66136 61162 66192
rect 61162 66136 61212 66192
rect 61148 66132 61212 66136
rect 63540 66192 63604 66196
rect 63540 66136 63590 66192
rect 63590 66136 63604 66192
rect 63540 66132 63604 66136
rect 66116 66192 66180 66196
rect 66116 66136 66130 66192
rect 66130 66136 66180 66192
rect 66116 66132 66180 66136
rect 68508 66192 68572 66196
rect 68508 66136 68558 66192
rect 68558 66136 68572 66192
rect 68508 66132 68572 66136
rect 71084 66192 71148 66196
rect 71084 66136 71098 66192
rect 71098 66136 71148 66192
rect 71084 66132 71148 66136
rect 73476 66192 73540 66196
rect 73476 66136 73526 66192
rect 73526 66136 73540 66192
rect 73476 66132 73540 66136
rect 86172 66132 86236 66196
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 96376 65852 96440 65856
rect 96376 65796 96380 65852
rect 96380 65796 96436 65852
rect 96436 65796 96440 65852
rect 96376 65792 96440 65796
rect 96456 65852 96520 65856
rect 96456 65796 96460 65852
rect 96460 65796 96516 65852
rect 96516 65796 96520 65852
rect 96456 65792 96520 65796
rect 96536 65852 96600 65856
rect 96536 65796 96540 65852
rect 96540 65796 96596 65852
rect 96596 65796 96600 65852
rect 96536 65792 96600 65796
rect 96616 65852 96680 65856
rect 96616 65796 96620 65852
rect 96620 65796 96676 65852
rect 96676 65796 96680 65852
rect 96616 65792 96680 65796
rect 105924 65852 105988 65856
rect 105924 65796 105928 65852
rect 105928 65796 105984 65852
rect 105984 65796 105988 65852
rect 105924 65792 105988 65796
rect 106004 65852 106068 65856
rect 106004 65796 106008 65852
rect 106008 65796 106064 65852
rect 106064 65796 106068 65852
rect 106004 65792 106068 65796
rect 106084 65852 106148 65856
rect 106084 65796 106088 65852
rect 106088 65796 106144 65852
rect 106144 65796 106148 65852
rect 106084 65792 106148 65796
rect 106164 65852 106228 65856
rect 106164 65796 106168 65852
rect 106168 65796 106224 65852
rect 106224 65796 106228 65852
rect 106164 65792 106228 65796
rect 4876 65308 4940 65312
rect 4876 65252 4880 65308
rect 4880 65252 4936 65308
rect 4936 65252 4940 65308
rect 4876 65248 4940 65252
rect 4956 65308 5020 65312
rect 4956 65252 4960 65308
rect 4960 65252 5016 65308
rect 5016 65252 5020 65308
rect 4956 65248 5020 65252
rect 5036 65308 5100 65312
rect 5036 65252 5040 65308
rect 5040 65252 5096 65308
rect 5096 65252 5100 65308
rect 5036 65248 5100 65252
rect 5116 65308 5180 65312
rect 5116 65252 5120 65308
rect 5120 65252 5176 65308
rect 5176 65252 5180 65308
rect 5116 65248 5180 65252
rect 106660 65308 106724 65312
rect 106660 65252 106664 65308
rect 106664 65252 106720 65308
rect 106720 65252 106724 65308
rect 106660 65248 106724 65252
rect 106740 65308 106804 65312
rect 106740 65252 106744 65308
rect 106744 65252 106800 65308
rect 106800 65252 106804 65308
rect 106740 65248 106804 65252
rect 106820 65308 106884 65312
rect 106820 65252 106824 65308
rect 106824 65252 106880 65308
rect 106880 65252 106884 65308
rect 106820 65248 106884 65252
rect 106900 65308 106964 65312
rect 106900 65252 106904 65308
rect 106904 65252 106960 65308
rect 106960 65252 106964 65308
rect 106900 65248 106964 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 105924 64764 105988 64768
rect 105924 64708 105928 64764
rect 105928 64708 105984 64764
rect 105984 64708 105988 64764
rect 105924 64704 105988 64708
rect 106004 64764 106068 64768
rect 106004 64708 106008 64764
rect 106008 64708 106064 64764
rect 106064 64708 106068 64764
rect 106004 64704 106068 64708
rect 106084 64764 106148 64768
rect 106084 64708 106088 64764
rect 106088 64708 106144 64764
rect 106144 64708 106148 64764
rect 106084 64704 106148 64708
rect 106164 64764 106228 64768
rect 106164 64708 106168 64764
rect 106168 64708 106224 64764
rect 106224 64708 106228 64764
rect 106164 64704 106228 64708
rect 4876 64220 4940 64224
rect 4876 64164 4880 64220
rect 4880 64164 4936 64220
rect 4936 64164 4940 64220
rect 4876 64160 4940 64164
rect 4956 64220 5020 64224
rect 4956 64164 4960 64220
rect 4960 64164 5016 64220
rect 5016 64164 5020 64220
rect 4956 64160 5020 64164
rect 5036 64220 5100 64224
rect 5036 64164 5040 64220
rect 5040 64164 5096 64220
rect 5096 64164 5100 64220
rect 5036 64160 5100 64164
rect 5116 64220 5180 64224
rect 5116 64164 5120 64220
rect 5120 64164 5176 64220
rect 5176 64164 5180 64220
rect 5116 64160 5180 64164
rect 106660 64220 106724 64224
rect 106660 64164 106664 64220
rect 106664 64164 106720 64220
rect 106720 64164 106724 64220
rect 106660 64160 106724 64164
rect 106740 64220 106804 64224
rect 106740 64164 106744 64220
rect 106744 64164 106800 64220
rect 106800 64164 106804 64220
rect 106740 64160 106804 64164
rect 106820 64220 106884 64224
rect 106820 64164 106824 64220
rect 106824 64164 106880 64220
rect 106880 64164 106884 64220
rect 106820 64160 106884 64164
rect 106900 64220 106964 64224
rect 106900 64164 106904 64220
rect 106904 64164 106960 64220
rect 106960 64164 106964 64220
rect 106900 64160 106964 64164
rect 95858 64152 95922 64156
rect 95858 64096 95882 64152
rect 95882 64096 95922 64152
rect 95858 64092 95922 64096
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 105924 63676 105988 63680
rect 105924 63620 105928 63676
rect 105928 63620 105984 63676
rect 105984 63620 105988 63676
rect 105924 63616 105988 63620
rect 106004 63676 106068 63680
rect 106004 63620 106008 63676
rect 106008 63620 106064 63676
rect 106064 63620 106068 63676
rect 106004 63616 106068 63620
rect 106084 63676 106148 63680
rect 106084 63620 106088 63676
rect 106088 63620 106144 63676
rect 106144 63620 106148 63676
rect 106084 63616 106148 63620
rect 106164 63676 106228 63680
rect 106164 63620 106168 63676
rect 106168 63620 106224 63676
rect 106224 63620 106228 63676
rect 106164 63616 106228 63620
rect 4876 63132 4940 63136
rect 4876 63076 4880 63132
rect 4880 63076 4936 63132
rect 4936 63076 4940 63132
rect 4876 63072 4940 63076
rect 4956 63132 5020 63136
rect 4956 63076 4960 63132
rect 4960 63076 5016 63132
rect 5016 63076 5020 63132
rect 4956 63072 5020 63076
rect 5036 63132 5100 63136
rect 5036 63076 5040 63132
rect 5040 63076 5096 63132
rect 5096 63076 5100 63132
rect 5036 63072 5100 63076
rect 5116 63132 5180 63136
rect 5116 63076 5120 63132
rect 5120 63076 5176 63132
rect 5176 63076 5180 63132
rect 5116 63072 5180 63076
rect 106660 63132 106724 63136
rect 106660 63076 106664 63132
rect 106664 63076 106720 63132
rect 106720 63076 106724 63132
rect 106660 63072 106724 63076
rect 106740 63132 106804 63136
rect 106740 63076 106744 63132
rect 106744 63076 106800 63132
rect 106800 63076 106804 63132
rect 106740 63072 106804 63076
rect 106820 63132 106884 63136
rect 106820 63076 106824 63132
rect 106824 63076 106880 63132
rect 106880 63076 106884 63132
rect 106820 63072 106884 63076
rect 106900 63132 106964 63136
rect 106900 63076 106904 63132
rect 106904 63076 106960 63132
rect 106960 63076 106964 63132
rect 106900 63072 106964 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 105924 62588 105988 62592
rect 105924 62532 105928 62588
rect 105928 62532 105984 62588
rect 105984 62532 105988 62588
rect 105924 62528 105988 62532
rect 106004 62588 106068 62592
rect 106004 62532 106008 62588
rect 106008 62532 106064 62588
rect 106064 62532 106068 62588
rect 106004 62528 106068 62532
rect 106084 62588 106148 62592
rect 106084 62532 106088 62588
rect 106088 62532 106144 62588
rect 106144 62532 106148 62588
rect 106084 62528 106148 62532
rect 106164 62588 106228 62592
rect 106164 62532 106168 62588
rect 106168 62532 106224 62588
rect 106224 62532 106228 62588
rect 106164 62528 106228 62532
rect 4876 62044 4940 62048
rect 4876 61988 4880 62044
rect 4880 61988 4936 62044
rect 4936 61988 4940 62044
rect 4876 61984 4940 61988
rect 4956 62044 5020 62048
rect 4956 61988 4960 62044
rect 4960 61988 5016 62044
rect 5016 61988 5020 62044
rect 4956 61984 5020 61988
rect 5036 62044 5100 62048
rect 5036 61988 5040 62044
rect 5040 61988 5096 62044
rect 5096 61988 5100 62044
rect 5036 61984 5100 61988
rect 5116 62044 5180 62048
rect 5116 61988 5120 62044
rect 5120 61988 5176 62044
rect 5176 61988 5180 62044
rect 5116 61984 5180 61988
rect 106660 62044 106724 62048
rect 106660 61988 106664 62044
rect 106664 61988 106720 62044
rect 106720 61988 106724 62044
rect 106660 61984 106724 61988
rect 106740 62044 106804 62048
rect 106740 61988 106744 62044
rect 106744 61988 106800 62044
rect 106800 61988 106804 62044
rect 106740 61984 106804 61988
rect 106820 62044 106884 62048
rect 106820 61988 106824 62044
rect 106824 61988 106880 62044
rect 106880 61988 106884 62044
rect 106820 61984 106884 61988
rect 106900 62044 106964 62048
rect 106900 61988 106904 62044
rect 106904 61988 106960 62044
rect 106960 61988 106964 62044
rect 106900 61984 106964 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 105924 61500 105988 61504
rect 105924 61444 105928 61500
rect 105928 61444 105984 61500
rect 105984 61444 105988 61500
rect 105924 61440 105988 61444
rect 106004 61500 106068 61504
rect 106004 61444 106008 61500
rect 106008 61444 106064 61500
rect 106064 61444 106068 61500
rect 106004 61440 106068 61444
rect 106084 61500 106148 61504
rect 106084 61444 106088 61500
rect 106088 61444 106144 61500
rect 106144 61444 106148 61500
rect 106084 61440 106148 61444
rect 106164 61500 106228 61504
rect 106164 61444 106168 61500
rect 106168 61444 106224 61500
rect 106224 61444 106228 61500
rect 106164 61440 106228 61444
rect 4876 60956 4940 60960
rect 4876 60900 4880 60956
rect 4880 60900 4936 60956
rect 4936 60900 4940 60956
rect 4876 60896 4940 60900
rect 4956 60956 5020 60960
rect 4956 60900 4960 60956
rect 4960 60900 5016 60956
rect 5016 60900 5020 60956
rect 4956 60896 5020 60900
rect 5036 60956 5100 60960
rect 5036 60900 5040 60956
rect 5040 60900 5096 60956
rect 5096 60900 5100 60956
rect 5036 60896 5100 60900
rect 5116 60956 5180 60960
rect 5116 60900 5120 60956
rect 5120 60900 5176 60956
rect 5176 60900 5180 60956
rect 5116 60896 5180 60900
rect 106660 60956 106724 60960
rect 106660 60900 106664 60956
rect 106664 60900 106720 60956
rect 106720 60900 106724 60956
rect 106660 60896 106724 60900
rect 106740 60956 106804 60960
rect 106740 60900 106744 60956
rect 106744 60900 106800 60956
rect 106800 60900 106804 60956
rect 106740 60896 106804 60900
rect 106820 60956 106884 60960
rect 106820 60900 106824 60956
rect 106824 60900 106880 60956
rect 106880 60900 106884 60956
rect 106820 60896 106884 60900
rect 106900 60956 106964 60960
rect 106900 60900 106904 60956
rect 106904 60900 106960 60956
rect 106960 60900 106964 60956
rect 106900 60896 106964 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 105924 60412 105988 60416
rect 105924 60356 105928 60412
rect 105928 60356 105984 60412
rect 105984 60356 105988 60412
rect 105924 60352 105988 60356
rect 106004 60412 106068 60416
rect 106004 60356 106008 60412
rect 106008 60356 106064 60412
rect 106064 60356 106068 60412
rect 106004 60352 106068 60356
rect 106084 60412 106148 60416
rect 106084 60356 106088 60412
rect 106088 60356 106144 60412
rect 106144 60356 106148 60412
rect 106084 60352 106148 60356
rect 106164 60412 106228 60416
rect 106164 60356 106168 60412
rect 106168 60356 106224 60412
rect 106224 60356 106228 60412
rect 106164 60352 106228 60356
rect 4876 59868 4940 59872
rect 4876 59812 4880 59868
rect 4880 59812 4936 59868
rect 4936 59812 4940 59868
rect 4876 59808 4940 59812
rect 4956 59868 5020 59872
rect 4956 59812 4960 59868
rect 4960 59812 5016 59868
rect 5016 59812 5020 59868
rect 4956 59808 5020 59812
rect 5036 59868 5100 59872
rect 5036 59812 5040 59868
rect 5040 59812 5096 59868
rect 5096 59812 5100 59868
rect 5036 59808 5100 59812
rect 5116 59868 5180 59872
rect 5116 59812 5120 59868
rect 5120 59812 5176 59868
rect 5176 59812 5180 59868
rect 5116 59808 5180 59812
rect 106660 59868 106724 59872
rect 106660 59812 106664 59868
rect 106664 59812 106720 59868
rect 106720 59812 106724 59868
rect 106660 59808 106724 59812
rect 106740 59868 106804 59872
rect 106740 59812 106744 59868
rect 106744 59812 106800 59868
rect 106800 59812 106804 59868
rect 106740 59808 106804 59812
rect 106820 59868 106884 59872
rect 106820 59812 106824 59868
rect 106824 59812 106880 59868
rect 106880 59812 106884 59868
rect 106820 59808 106884 59812
rect 106900 59868 106964 59872
rect 106900 59812 106904 59868
rect 106904 59812 106960 59868
rect 106960 59812 106964 59868
rect 106900 59808 106964 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 105924 59324 105988 59328
rect 105924 59268 105928 59324
rect 105928 59268 105984 59324
rect 105984 59268 105988 59324
rect 105924 59264 105988 59268
rect 106004 59324 106068 59328
rect 106004 59268 106008 59324
rect 106008 59268 106064 59324
rect 106064 59268 106068 59324
rect 106004 59264 106068 59268
rect 106084 59324 106148 59328
rect 106084 59268 106088 59324
rect 106088 59268 106144 59324
rect 106144 59268 106148 59324
rect 106084 59264 106148 59268
rect 106164 59324 106228 59328
rect 106164 59268 106168 59324
rect 106168 59268 106224 59324
rect 106224 59268 106228 59324
rect 106164 59264 106228 59268
rect 4876 58780 4940 58784
rect 4876 58724 4880 58780
rect 4880 58724 4936 58780
rect 4936 58724 4940 58780
rect 4876 58720 4940 58724
rect 4956 58780 5020 58784
rect 4956 58724 4960 58780
rect 4960 58724 5016 58780
rect 5016 58724 5020 58780
rect 4956 58720 5020 58724
rect 5036 58780 5100 58784
rect 5036 58724 5040 58780
rect 5040 58724 5096 58780
rect 5096 58724 5100 58780
rect 5036 58720 5100 58724
rect 5116 58780 5180 58784
rect 5116 58724 5120 58780
rect 5120 58724 5176 58780
rect 5176 58724 5180 58780
rect 5116 58720 5180 58724
rect 106660 58780 106724 58784
rect 106660 58724 106664 58780
rect 106664 58724 106720 58780
rect 106720 58724 106724 58780
rect 106660 58720 106724 58724
rect 106740 58780 106804 58784
rect 106740 58724 106744 58780
rect 106744 58724 106800 58780
rect 106800 58724 106804 58780
rect 106740 58720 106804 58724
rect 106820 58780 106884 58784
rect 106820 58724 106824 58780
rect 106824 58724 106880 58780
rect 106880 58724 106884 58780
rect 106820 58720 106884 58724
rect 106900 58780 106964 58784
rect 106900 58724 106904 58780
rect 106904 58724 106960 58780
rect 106960 58724 106964 58780
rect 106900 58720 106964 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 105924 58236 105988 58240
rect 105924 58180 105928 58236
rect 105928 58180 105984 58236
rect 105984 58180 105988 58236
rect 105924 58176 105988 58180
rect 106004 58236 106068 58240
rect 106004 58180 106008 58236
rect 106008 58180 106064 58236
rect 106064 58180 106068 58236
rect 106004 58176 106068 58180
rect 106084 58236 106148 58240
rect 106084 58180 106088 58236
rect 106088 58180 106144 58236
rect 106144 58180 106148 58236
rect 106084 58176 106148 58180
rect 106164 58236 106228 58240
rect 106164 58180 106168 58236
rect 106168 58180 106224 58236
rect 106224 58180 106228 58236
rect 106164 58176 106228 58180
rect 4876 57692 4940 57696
rect 4876 57636 4880 57692
rect 4880 57636 4936 57692
rect 4936 57636 4940 57692
rect 4876 57632 4940 57636
rect 4956 57692 5020 57696
rect 4956 57636 4960 57692
rect 4960 57636 5016 57692
rect 5016 57636 5020 57692
rect 4956 57632 5020 57636
rect 5036 57692 5100 57696
rect 5036 57636 5040 57692
rect 5040 57636 5096 57692
rect 5096 57636 5100 57692
rect 5036 57632 5100 57636
rect 5116 57692 5180 57696
rect 5116 57636 5120 57692
rect 5120 57636 5176 57692
rect 5176 57636 5180 57692
rect 5116 57632 5180 57636
rect 106660 57692 106724 57696
rect 106660 57636 106664 57692
rect 106664 57636 106720 57692
rect 106720 57636 106724 57692
rect 106660 57632 106724 57636
rect 106740 57692 106804 57696
rect 106740 57636 106744 57692
rect 106744 57636 106800 57692
rect 106800 57636 106804 57692
rect 106740 57632 106804 57636
rect 106820 57692 106884 57696
rect 106820 57636 106824 57692
rect 106824 57636 106880 57692
rect 106880 57636 106884 57692
rect 106820 57632 106884 57636
rect 106900 57692 106964 57696
rect 106900 57636 106904 57692
rect 106904 57636 106960 57692
rect 106960 57636 106964 57692
rect 106900 57632 106964 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 105924 57148 105988 57152
rect 105924 57092 105928 57148
rect 105928 57092 105984 57148
rect 105984 57092 105988 57148
rect 105924 57088 105988 57092
rect 106004 57148 106068 57152
rect 106004 57092 106008 57148
rect 106008 57092 106064 57148
rect 106064 57092 106068 57148
rect 106004 57088 106068 57092
rect 106084 57148 106148 57152
rect 106084 57092 106088 57148
rect 106088 57092 106144 57148
rect 106144 57092 106148 57148
rect 106084 57088 106148 57092
rect 106164 57148 106228 57152
rect 106164 57092 106168 57148
rect 106168 57092 106224 57148
rect 106224 57092 106228 57148
rect 106164 57088 106228 57092
rect 4876 56604 4940 56608
rect 4876 56548 4880 56604
rect 4880 56548 4936 56604
rect 4936 56548 4940 56604
rect 4876 56544 4940 56548
rect 4956 56604 5020 56608
rect 4956 56548 4960 56604
rect 4960 56548 5016 56604
rect 5016 56548 5020 56604
rect 4956 56544 5020 56548
rect 5036 56604 5100 56608
rect 5036 56548 5040 56604
rect 5040 56548 5096 56604
rect 5096 56548 5100 56604
rect 5036 56544 5100 56548
rect 5116 56604 5180 56608
rect 5116 56548 5120 56604
rect 5120 56548 5176 56604
rect 5176 56548 5180 56604
rect 5116 56544 5180 56548
rect 106660 56604 106724 56608
rect 106660 56548 106664 56604
rect 106664 56548 106720 56604
rect 106720 56548 106724 56604
rect 106660 56544 106724 56548
rect 106740 56604 106804 56608
rect 106740 56548 106744 56604
rect 106744 56548 106800 56604
rect 106800 56548 106804 56604
rect 106740 56544 106804 56548
rect 106820 56604 106884 56608
rect 106820 56548 106824 56604
rect 106824 56548 106880 56604
rect 106880 56548 106884 56604
rect 106820 56544 106884 56548
rect 106900 56604 106964 56608
rect 106900 56548 106904 56604
rect 106904 56548 106960 56604
rect 106960 56548 106964 56604
rect 106900 56544 106964 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 105924 56060 105988 56064
rect 105924 56004 105928 56060
rect 105928 56004 105984 56060
rect 105984 56004 105988 56060
rect 105924 56000 105988 56004
rect 106004 56060 106068 56064
rect 106004 56004 106008 56060
rect 106008 56004 106064 56060
rect 106064 56004 106068 56060
rect 106004 56000 106068 56004
rect 106084 56060 106148 56064
rect 106084 56004 106088 56060
rect 106088 56004 106144 56060
rect 106144 56004 106148 56060
rect 106084 56000 106148 56004
rect 106164 56060 106228 56064
rect 106164 56004 106168 56060
rect 106168 56004 106224 56060
rect 106224 56004 106228 56060
rect 106164 56000 106228 56004
rect 4876 55516 4940 55520
rect 4876 55460 4880 55516
rect 4880 55460 4936 55516
rect 4936 55460 4940 55516
rect 4876 55456 4940 55460
rect 4956 55516 5020 55520
rect 4956 55460 4960 55516
rect 4960 55460 5016 55516
rect 5016 55460 5020 55516
rect 4956 55456 5020 55460
rect 5036 55516 5100 55520
rect 5036 55460 5040 55516
rect 5040 55460 5096 55516
rect 5096 55460 5100 55516
rect 5036 55456 5100 55460
rect 5116 55516 5180 55520
rect 5116 55460 5120 55516
rect 5120 55460 5176 55516
rect 5176 55460 5180 55516
rect 5116 55456 5180 55460
rect 106660 55516 106724 55520
rect 106660 55460 106664 55516
rect 106664 55460 106720 55516
rect 106720 55460 106724 55516
rect 106660 55456 106724 55460
rect 106740 55516 106804 55520
rect 106740 55460 106744 55516
rect 106744 55460 106800 55516
rect 106800 55460 106804 55516
rect 106740 55456 106804 55460
rect 106820 55516 106884 55520
rect 106820 55460 106824 55516
rect 106824 55460 106880 55516
rect 106880 55460 106884 55516
rect 106820 55456 106884 55460
rect 106900 55516 106964 55520
rect 106900 55460 106904 55516
rect 106904 55460 106960 55516
rect 106960 55460 106964 55516
rect 106900 55456 106964 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 105924 54972 105988 54976
rect 105924 54916 105928 54972
rect 105928 54916 105984 54972
rect 105984 54916 105988 54972
rect 105924 54912 105988 54916
rect 106004 54972 106068 54976
rect 106004 54916 106008 54972
rect 106008 54916 106064 54972
rect 106064 54916 106068 54972
rect 106004 54912 106068 54916
rect 106084 54972 106148 54976
rect 106084 54916 106088 54972
rect 106088 54916 106144 54972
rect 106144 54916 106148 54972
rect 106084 54912 106148 54916
rect 106164 54972 106228 54976
rect 106164 54916 106168 54972
rect 106168 54916 106224 54972
rect 106224 54916 106228 54972
rect 106164 54912 106228 54916
rect 4876 54428 4940 54432
rect 4876 54372 4880 54428
rect 4880 54372 4936 54428
rect 4936 54372 4940 54428
rect 4876 54368 4940 54372
rect 4956 54428 5020 54432
rect 4956 54372 4960 54428
rect 4960 54372 5016 54428
rect 5016 54372 5020 54428
rect 4956 54368 5020 54372
rect 5036 54428 5100 54432
rect 5036 54372 5040 54428
rect 5040 54372 5096 54428
rect 5096 54372 5100 54428
rect 5036 54368 5100 54372
rect 5116 54428 5180 54432
rect 5116 54372 5120 54428
rect 5120 54372 5176 54428
rect 5176 54372 5180 54428
rect 5116 54368 5180 54372
rect 106660 54428 106724 54432
rect 106660 54372 106664 54428
rect 106664 54372 106720 54428
rect 106720 54372 106724 54428
rect 106660 54368 106724 54372
rect 106740 54428 106804 54432
rect 106740 54372 106744 54428
rect 106744 54372 106800 54428
rect 106800 54372 106804 54428
rect 106740 54368 106804 54372
rect 106820 54428 106884 54432
rect 106820 54372 106824 54428
rect 106824 54372 106880 54428
rect 106880 54372 106884 54428
rect 106820 54368 106884 54372
rect 106900 54428 106964 54432
rect 106900 54372 106904 54428
rect 106904 54372 106960 54428
rect 106960 54372 106964 54428
rect 106900 54368 106964 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 105924 53884 105988 53888
rect 105924 53828 105928 53884
rect 105928 53828 105984 53884
rect 105984 53828 105988 53884
rect 105924 53824 105988 53828
rect 106004 53884 106068 53888
rect 106004 53828 106008 53884
rect 106008 53828 106064 53884
rect 106064 53828 106068 53884
rect 106004 53824 106068 53828
rect 106084 53884 106148 53888
rect 106084 53828 106088 53884
rect 106088 53828 106144 53884
rect 106144 53828 106148 53884
rect 106084 53824 106148 53828
rect 106164 53884 106228 53888
rect 106164 53828 106168 53884
rect 106168 53828 106224 53884
rect 106224 53828 106228 53884
rect 106164 53824 106228 53828
rect 4876 53340 4940 53344
rect 4876 53284 4880 53340
rect 4880 53284 4936 53340
rect 4936 53284 4940 53340
rect 4876 53280 4940 53284
rect 4956 53340 5020 53344
rect 4956 53284 4960 53340
rect 4960 53284 5016 53340
rect 5016 53284 5020 53340
rect 4956 53280 5020 53284
rect 5036 53340 5100 53344
rect 5036 53284 5040 53340
rect 5040 53284 5096 53340
rect 5096 53284 5100 53340
rect 5036 53280 5100 53284
rect 5116 53340 5180 53344
rect 5116 53284 5120 53340
rect 5120 53284 5176 53340
rect 5176 53284 5180 53340
rect 5116 53280 5180 53284
rect 106660 53340 106724 53344
rect 106660 53284 106664 53340
rect 106664 53284 106720 53340
rect 106720 53284 106724 53340
rect 106660 53280 106724 53284
rect 106740 53340 106804 53344
rect 106740 53284 106744 53340
rect 106744 53284 106800 53340
rect 106800 53284 106804 53340
rect 106740 53280 106804 53284
rect 106820 53340 106884 53344
rect 106820 53284 106824 53340
rect 106824 53284 106880 53340
rect 106880 53284 106884 53340
rect 106820 53280 106884 53284
rect 106900 53340 106964 53344
rect 106900 53284 106904 53340
rect 106904 53284 106960 53340
rect 106960 53284 106964 53340
rect 106900 53280 106964 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 105924 52796 105988 52800
rect 105924 52740 105928 52796
rect 105928 52740 105984 52796
rect 105984 52740 105988 52796
rect 105924 52736 105988 52740
rect 106004 52796 106068 52800
rect 106004 52740 106008 52796
rect 106008 52740 106064 52796
rect 106064 52740 106068 52796
rect 106004 52736 106068 52740
rect 106084 52796 106148 52800
rect 106084 52740 106088 52796
rect 106088 52740 106144 52796
rect 106144 52740 106148 52796
rect 106084 52736 106148 52740
rect 106164 52796 106228 52800
rect 106164 52740 106168 52796
rect 106168 52740 106224 52796
rect 106224 52740 106228 52796
rect 106164 52736 106228 52740
rect 4876 52252 4940 52256
rect 4876 52196 4880 52252
rect 4880 52196 4936 52252
rect 4936 52196 4940 52252
rect 4876 52192 4940 52196
rect 4956 52252 5020 52256
rect 4956 52196 4960 52252
rect 4960 52196 5016 52252
rect 5016 52196 5020 52252
rect 4956 52192 5020 52196
rect 5036 52252 5100 52256
rect 5036 52196 5040 52252
rect 5040 52196 5096 52252
rect 5096 52196 5100 52252
rect 5036 52192 5100 52196
rect 5116 52252 5180 52256
rect 5116 52196 5120 52252
rect 5120 52196 5176 52252
rect 5176 52196 5180 52252
rect 5116 52192 5180 52196
rect 106660 52252 106724 52256
rect 106660 52196 106664 52252
rect 106664 52196 106720 52252
rect 106720 52196 106724 52252
rect 106660 52192 106724 52196
rect 106740 52252 106804 52256
rect 106740 52196 106744 52252
rect 106744 52196 106800 52252
rect 106800 52196 106804 52252
rect 106740 52192 106804 52196
rect 106820 52252 106884 52256
rect 106820 52196 106824 52252
rect 106824 52196 106880 52252
rect 106880 52196 106884 52252
rect 106820 52192 106884 52196
rect 106900 52252 106964 52256
rect 106900 52196 106904 52252
rect 106904 52196 106960 52252
rect 106960 52196 106964 52252
rect 106900 52192 106964 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 105924 51708 105988 51712
rect 105924 51652 105928 51708
rect 105928 51652 105984 51708
rect 105984 51652 105988 51708
rect 105924 51648 105988 51652
rect 106004 51708 106068 51712
rect 106004 51652 106008 51708
rect 106008 51652 106064 51708
rect 106064 51652 106068 51708
rect 106004 51648 106068 51652
rect 106084 51708 106148 51712
rect 106084 51652 106088 51708
rect 106088 51652 106144 51708
rect 106144 51652 106148 51708
rect 106084 51648 106148 51652
rect 106164 51708 106228 51712
rect 106164 51652 106168 51708
rect 106168 51652 106224 51708
rect 106224 51652 106228 51708
rect 106164 51648 106228 51652
rect 4876 51164 4940 51168
rect 4876 51108 4880 51164
rect 4880 51108 4936 51164
rect 4936 51108 4940 51164
rect 4876 51104 4940 51108
rect 4956 51164 5020 51168
rect 4956 51108 4960 51164
rect 4960 51108 5016 51164
rect 5016 51108 5020 51164
rect 4956 51104 5020 51108
rect 5036 51164 5100 51168
rect 5036 51108 5040 51164
rect 5040 51108 5096 51164
rect 5096 51108 5100 51164
rect 5036 51104 5100 51108
rect 5116 51164 5180 51168
rect 5116 51108 5120 51164
rect 5120 51108 5176 51164
rect 5176 51108 5180 51164
rect 5116 51104 5180 51108
rect 106660 51164 106724 51168
rect 106660 51108 106664 51164
rect 106664 51108 106720 51164
rect 106720 51108 106724 51164
rect 106660 51104 106724 51108
rect 106740 51164 106804 51168
rect 106740 51108 106744 51164
rect 106744 51108 106800 51164
rect 106800 51108 106804 51164
rect 106740 51104 106804 51108
rect 106820 51164 106884 51168
rect 106820 51108 106824 51164
rect 106824 51108 106880 51164
rect 106880 51108 106884 51164
rect 106820 51104 106884 51108
rect 106900 51164 106964 51168
rect 106900 51108 106904 51164
rect 106904 51108 106960 51164
rect 106960 51108 106964 51164
rect 106900 51104 106964 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 105924 50620 105988 50624
rect 105924 50564 105928 50620
rect 105928 50564 105984 50620
rect 105984 50564 105988 50620
rect 105924 50560 105988 50564
rect 106004 50620 106068 50624
rect 106004 50564 106008 50620
rect 106008 50564 106064 50620
rect 106064 50564 106068 50620
rect 106004 50560 106068 50564
rect 106084 50620 106148 50624
rect 106084 50564 106088 50620
rect 106088 50564 106144 50620
rect 106144 50564 106148 50620
rect 106084 50560 106148 50564
rect 106164 50620 106228 50624
rect 106164 50564 106168 50620
rect 106168 50564 106224 50620
rect 106224 50564 106228 50620
rect 106164 50560 106228 50564
rect 4876 50076 4940 50080
rect 4876 50020 4880 50076
rect 4880 50020 4936 50076
rect 4936 50020 4940 50076
rect 4876 50016 4940 50020
rect 4956 50076 5020 50080
rect 4956 50020 4960 50076
rect 4960 50020 5016 50076
rect 5016 50020 5020 50076
rect 4956 50016 5020 50020
rect 5036 50076 5100 50080
rect 5036 50020 5040 50076
rect 5040 50020 5096 50076
rect 5096 50020 5100 50076
rect 5036 50016 5100 50020
rect 5116 50076 5180 50080
rect 5116 50020 5120 50076
rect 5120 50020 5176 50076
rect 5176 50020 5180 50076
rect 5116 50016 5180 50020
rect 106660 50076 106724 50080
rect 106660 50020 106664 50076
rect 106664 50020 106720 50076
rect 106720 50020 106724 50076
rect 106660 50016 106724 50020
rect 106740 50076 106804 50080
rect 106740 50020 106744 50076
rect 106744 50020 106800 50076
rect 106800 50020 106804 50076
rect 106740 50016 106804 50020
rect 106820 50076 106884 50080
rect 106820 50020 106824 50076
rect 106824 50020 106880 50076
rect 106880 50020 106884 50076
rect 106820 50016 106884 50020
rect 106900 50076 106964 50080
rect 106900 50020 106904 50076
rect 106904 50020 106960 50076
rect 106960 50020 106964 50076
rect 106900 50016 106964 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 105924 49532 105988 49536
rect 105924 49476 105928 49532
rect 105928 49476 105984 49532
rect 105984 49476 105988 49532
rect 105924 49472 105988 49476
rect 106004 49532 106068 49536
rect 106004 49476 106008 49532
rect 106008 49476 106064 49532
rect 106064 49476 106068 49532
rect 106004 49472 106068 49476
rect 106084 49532 106148 49536
rect 106084 49476 106088 49532
rect 106088 49476 106144 49532
rect 106144 49476 106148 49532
rect 106084 49472 106148 49476
rect 106164 49532 106228 49536
rect 106164 49476 106168 49532
rect 106168 49476 106224 49532
rect 106224 49476 106228 49532
rect 106164 49472 106228 49476
rect 4876 48988 4940 48992
rect 4876 48932 4880 48988
rect 4880 48932 4936 48988
rect 4936 48932 4940 48988
rect 4876 48928 4940 48932
rect 4956 48988 5020 48992
rect 4956 48932 4960 48988
rect 4960 48932 5016 48988
rect 5016 48932 5020 48988
rect 4956 48928 5020 48932
rect 5036 48988 5100 48992
rect 5036 48932 5040 48988
rect 5040 48932 5096 48988
rect 5096 48932 5100 48988
rect 5036 48928 5100 48932
rect 5116 48988 5180 48992
rect 5116 48932 5120 48988
rect 5120 48932 5176 48988
rect 5176 48932 5180 48988
rect 5116 48928 5180 48932
rect 106660 48988 106724 48992
rect 106660 48932 106664 48988
rect 106664 48932 106720 48988
rect 106720 48932 106724 48988
rect 106660 48928 106724 48932
rect 106740 48988 106804 48992
rect 106740 48932 106744 48988
rect 106744 48932 106800 48988
rect 106800 48932 106804 48988
rect 106740 48928 106804 48932
rect 106820 48988 106884 48992
rect 106820 48932 106824 48988
rect 106824 48932 106880 48988
rect 106880 48932 106884 48988
rect 106820 48928 106884 48932
rect 106900 48988 106964 48992
rect 106900 48932 106904 48988
rect 106904 48932 106960 48988
rect 106960 48932 106964 48988
rect 106900 48928 106964 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 105924 48444 105988 48448
rect 105924 48388 105928 48444
rect 105928 48388 105984 48444
rect 105984 48388 105988 48444
rect 105924 48384 105988 48388
rect 106004 48444 106068 48448
rect 106004 48388 106008 48444
rect 106008 48388 106064 48444
rect 106064 48388 106068 48444
rect 106004 48384 106068 48388
rect 106084 48444 106148 48448
rect 106084 48388 106088 48444
rect 106088 48388 106144 48444
rect 106144 48388 106148 48444
rect 106084 48384 106148 48388
rect 106164 48444 106228 48448
rect 106164 48388 106168 48444
rect 106168 48388 106224 48444
rect 106224 48388 106228 48444
rect 106164 48384 106228 48388
rect 4876 47900 4940 47904
rect 4876 47844 4880 47900
rect 4880 47844 4936 47900
rect 4936 47844 4940 47900
rect 4876 47840 4940 47844
rect 4956 47900 5020 47904
rect 4956 47844 4960 47900
rect 4960 47844 5016 47900
rect 5016 47844 5020 47900
rect 4956 47840 5020 47844
rect 5036 47900 5100 47904
rect 5036 47844 5040 47900
rect 5040 47844 5096 47900
rect 5096 47844 5100 47900
rect 5036 47840 5100 47844
rect 5116 47900 5180 47904
rect 5116 47844 5120 47900
rect 5120 47844 5176 47900
rect 5176 47844 5180 47900
rect 5116 47840 5180 47844
rect 106660 47900 106724 47904
rect 106660 47844 106664 47900
rect 106664 47844 106720 47900
rect 106720 47844 106724 47900
rect 106660 47840 106724 47844
rect 106740 47900 106804 47904
rect 106740 47844 106744 47900
rect 106744 47844 106800 47900
rect 106800 47844 106804 47900
rect 106740 47840 106804 47844
rect 106820 47900 106884 47904
rect 106820 47844 106824 47900
rect 106824 47844 106880 47900
rect 106880 47844 106884 47900
rect 106820 47840 106884 47844
rect 106900 47900 106964 47904
rect 106900 47844 106904 47900
rect 106904 47844 106960 47900
rect 106960 47844 106964 47900
rect 106900 47840 106964 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 105924 47356 105988 47360
rect 105924 47300 105928 47356
rect 105928 47300 105984 47356
rect 105984 47300 105988 47356
rect 105924 47296 105988 47300
rect 106004 47356 106068 47360
rect 106004 47300 106008 47356
rect 106008 47300 106064 47356
rect 106064 47300 106068 47356
rect 106004 47296 106068 47300
rect 106084 47356 106148 47360
rect 106084 47300 106088 47356
rect 106088 47300 106144 47356
rect 106144 47300 106148 47356
rect 106084 47296 106148 47300
rect 106164 47356 106228 47360
rect 106164 47300 106168 47356
rect 106168 47300 106224 47356
rect 106224 47300 106228 47356
rect 106164 47296 106228 47300
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 106660 46812 106724 46816
rect 106660 46756 106664 46812
rect 106664 46756 106720 46812
rect 106720 46756 106724 46812
rect 106660 46752 106724 46756
rect 106740 46812 106804 46816
rect 106740 46756 106744 46812
rect 106744 46756 106800 46812
rect 106800 46756 106804 46812
rect 106740 46752 106804 46756
rect 106820 46812 106884 46816
rect 106820 46756 106824 46812
rect 106824 46756 106880 46812
rect 106880 46756 106884 46812
rect 106820 46752 106884 46756
rect 106900 46812 106964 46816
rect 106900 46756 106904 46812
rect 106904 46756 106960 46812
rect 106960 46756 106964 46812
rect 106900 46752 106964 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 105924 46268 105988 46272
rect 105924 46212 105928 46268
rect 105928 46212 105984 46268
rect 105984 46212 105988 46268
rect 105924 46208 105988 46212
rect 106004 46268 106068 46272
rect 106004 46212 106008 46268
rect 106008 46212 106064 46268
rect 106064 46212 106068 46268
rect 106004 46208 106068 46212
rect 106084 46268 106148 46272
rect 106084 46212 106088 46268
rect 106088 46212 106144 46268
rect 106144 46212 106148 46268
rect 106084 46208 106148 46212
rect 106164 46268 106228 46272
rect 106164 46212 106168 46268
rect 106168 46212 106224 46268
rect 106224 46212 106228 46268
rect 106164 46208 106228 46212
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 106660 45724 106724 45728
rect 106660 45668 106664 45724
rect 106664 45668 106720 45724
rect 106720 45668 106724 45724
rect 106660 45664 106724 45668
rect 106740 45724 106804 45728
rect 106740 45668 106744 45724
rect 106744 45668 106800 45724
rect 106800 45668 106804 45724
rect 106740 45664 106804 45668
rect 106820 45724 106884 45728
rect 106820 45668 106824 45724
rect 106824 45668 106880 45724
rect 106880 45668 106884 45724
rect 106820 45664 106884 45668
rect 106900 45724 106964 45728
rect 106900 45668 106904 45724
rect 106904 45668 106960 45724
rect 106960 45668 106964 45724
rect 106900 45664 106964 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 105924 45180 105988 45184
rect 105924 45124 105928 45180
rect 105928 45124 105984 45180
rect 105984 45124 105988 45180
rect 105924 45120 105988 45124
rect 106004 45180 106068 45184
rect 106004 45124 106008 45180
rect 106008 45124 106064 45180
rect 106064 45124 106068 45180
rect 106004 45120 106068 45124
rect 106084 45180 106148 45184
rect 106084 45124 106088 45180
rect 106088 45124 106144 45180
rect 106144 45124 106148 45180
rect 106084 45120 106148 45124
rect 106164 45180 106228 45184
rect 106164 45124 106168 45180
rect 106168 45124 106224 45180
rect 106224 45124 106228 45180
rect 106164 45120 106228 45124
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 106660 44636 106724 44640
rect 106660 44580 106664 44636
rect 106664 44580 106720 44636
rect 106720 44580 106724 44636
rect 106660 44576 106724 44580
rect 106740 44636 106804 44640
rect 106740 44580 106744 44636
rect 106744 44580 106800 44636
rect 106800 44580 106804 44636
rect 106740 44576 106804 44580
rect 106820 44636 106884 44640
rect 106820 44580 106824 44636
rect 106824 44580 106880 44636
rect 106880 44580 106884 44636
rect 106820 44576 106884 44580
rect 106900 44636 106964 44640
rect 106900 44580 106904 44636
rect 106904 44580 106960 44636
rect 106960 44580 106964 44636
rect 106900 44576 106964 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 105924 44092 105988 44096
rect 105924 44036 105928 44092
rect 105928 44036 105984 44092
rect 105984 44036 105988 44092
rect 105924 44032 105988 44036
rect 106004 44092 106068 44096
rect 106004 44036 106008 44092
rect 106008 44036 106064 44092
rect 106064 44036 106068 44092
rect 106004 44032 106068 44036
rect 106084 44092 106148 44096
rect 106084 44036 106088 44092
rect 106088 44036 106144 44092
rect 106144 44036 106148 44092
rect 106084 44032 106148 44036
rect 106164 44092 106228 44096
rect 106164 44036 106168 44092
rect 106168 44036 106224 44092
rect 106224 44036 106228 44092
rect 106164 44032 106228 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 106660 43548 106724 43552
rect 106660 43492 106664 43548
rect 106664 43492 106720 43548
rect 106720 43492 106724 43548
rect 106660 43488 106724 43492
rect 106740 43548 106804 43552
rect 106740 43492 106744 43548
rect 106744 43492 106800 43548
rect 106800 43492 106804 43548
rect 106740 43488 106804 43492
rect 106820 43548 106884 43552
rect 106820 43492 106824 43548
rect 106824 43492 106880 43548
rect 106880 43492 106884 43548
rect 106820 43488 106884 43492
rect 106900 43548 106964 43552
rect 106900 43492 106904 43548
rect 106904 43492 106960 43548
rect 106960 43492 106964 43548
rect 106900 43488 106964 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 105924 43004 105988 43008
rect 105924 42948 105928 43004
rect 105928 42948 105984 43004
rect 105984 42948 105988 43004
rect 105924 42944 105988 42948
rect 106004 43004 106068 43008
rect 106004 42948 106008 43004
rect 106008 42948 106064 43004
rect 106064 42948 106068 43004
rect 106004 42944 106068 42948
rect 106084 43004 106148 43008
rect 106084 42948 106088 43004
rect 106088 42948 106144 43004
rect 106144 42948 106148 43004
rect 106084 42944 106148 42948
rect 106164 43004 106228 43008
rect 106164 42948 106168 43004
rect 106168 42948 106224 43004
rect 106224 42948 106228 43004
rect 106164 42944 106228 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 106660 42460 106724 42464
rect 106660 42404 106664 42460
rect 106664 42404 106720 42460
rect 106720 42404 106724 42460
rect 106660 42400 106724 42404
rect 106740 42460 106804 42464
rect 106740 42404 106744 42460
rect 106744 42404 106800 42460
rect 106800 42404 106804 42460
rect 106740 42400 106804 42404
rect 106820 42460 106884 42464
rect 106820 42404 106824 42460
rect 106824 42404 106880 42460
rect 106880 42404 106884 42460
rect 106820 42400 106884 42404
rect 106900 42460 106964 42464
rect 106900 42404 106904 42460
rect 106904 42404 106960 42460
rect 106960 42404 106964 42460
rect 106900 42400 106964 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 105924 41916 105988 41920
rect 105924 41860 105928 41916
rect 105928 41860 105984 41916
rect 105984 41860 105988 41916
rect 105924 41856 105988 41860
rect 106004 41916 106068 41920
rect 106004 41860 106008 41916
rect 106008 41860 106064 41916
rect 106064 41860 106068 41916
rect 106004 41856 106068 41860
rect 106084 41916 106148 41920
rect 106084 41860 106088 41916
rect 106088 41860 106144 41916
rect 106144 41860 106148 41916
rect 106084 41856 106148 41860
rect 106164 41916 106228 41920
rect 106164 41860 106168 41916
rect 106168 41860 106224 41916
rect 106224 41860 106228 41916
rect 106164 41856 106228 41860
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 106660 41372 106724 41376
rect 106660 41316 106664 41372
rect 106664 41316 106720 41372
rect 106720 41316 106724 41372
rect 106660 41312 106724 41316
rect 106740 41372 106804 41376
rect 106740 41316 106744 41372
rect 106744 41316 106800 41372
rect 106800 41316 106804 41372
rect 106740 41312 106804 41316
rect 106820 41372 106884 41376
rect 106820 41316 106824 41372
rect 106824 41316 106880 41372
rect 106880 41316 106884 41372
rect 106820 41312 106884 41316
rect 106900 41372 106964 41376
rect 106900 41316 106904 41372
rect 106904 41316 106960 41372
rect 106960 41316 106964 41372
rect 106900 41312 106964 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 105924 40828 105988 40832
rect 105924 40772 105928 40828
rect 105928 40772 105984 40828
rect 105984 40772 105988 40828
rect 105924 40768 105988 40772
rect 106004 40828 106068 40832
rect 106004 40772 106008 40828
rect 106008 40772 106064 40828
rect 106064 40772 106068 40828
rect 106004 40768 106068 40772
rect 106084 40828 106148 40832
rect 106084 40772 106088 40828
rect 106088 40772 106144 40828
rect 106144 40772 106148 40828
rect 106084 40768 106148 40772
rect 106164 40828 106228 40832
rect 106164 40772 106168 40828
rect 106168 40772 106224 40828
rect 106224 40772 106228 40828
rect 106164 40768 106228 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 106660 40284 106724 40288
rect 106660 40228 106664 40284
rect 106664 40228 106720 40284
rect 106720 40228 106724 40284
rect 106660 40224 106724 40228
rect 106740 40284 106804 40288
rect 106740 40228 106744 40284
rect 106744 40228 106800 40284
rect 106800 40228 106804 40284
rect 106740 40224 106804 40228
rect 106820 40284 106884 40288
rect 106820 40228 106824 40284
rect 106824 40228 106880 40284
rect 106880 40228 106884 40284
rect 106820 40224 106884 40228
rect 106900 40284 106964 40288
rect 106900 40228 106904 40284
rect 106904 40228 106960 40284
rect 106960 40228 106964 40284
rect 106900 40224 106964 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 105924 39740 105988 39744
rect 105924 39684 105928 39740
rect 105928 39684 105984 39740
rect 105984 39684 105988 39740
rect 105924 39680 105988 39684
rect 106004 39740 106068 39744
rect 106004 39684 106008 39740
rect 106008 39684 106064 39740
rect 106064 39684 106068 39740
rect 106004 39680 106068 39684
rect 106084 39740 106148 39744
rect 106084 39684 106088 39740
rect 106088 39684 106144 39740
rect 106144 39684 106148 39740
rect 106084 39680 106148 39684
rect 106164 39740 106228 39744
rect 106164 39684 106168 39740
rect 106168 39684 106224 39740
rect 106224 39684 106228 39740
rect 106164 39680 106228 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 106660 39196 106724 39200
rect 106660 39140 106664 39196
rect 106664 39140 106720 39196
rect 106720 39140 106724 39196
rect 106660 39136 106724 39140
rect 106740 39196 106804 39200
rect 106740 39140 106744 39196
rect 106744 39140 106800 39196
rect 106800 39140 106804 39196
rect 106740 39136 106804 39140
rect 106820 39196 106884 39200
rect 106820 39140 106824 39196
rect 106824 39140 106880 39196
rect 106880 39140 106884 39196
rect 106820 39136 106884 39140
rect 106900 39196 106964 39200
rect 106900 39140 106904 39196
rect 106904 39140 106960 39196
rect 106960 39140 106964 39196
rect 106900 39136 106964 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 105924 38652 105988 38656
rect 105924 38596 105928 38652
rect 105928 38596 105984 38652
rect 105984 38596 105988 38652
rect 105924 38592 105988 38596
rect 106004 38652 106068 38656
rect 106004 38596 106008 38652
rect 106008 38596 106064 38652
rect 106064 38596 106068 38652
rect 106004 38592 106068 38596
rect 106084 38652 106148 38656
rect 106084 38596 106088 38652
rect 106088 38596 106144 38652
rect 106144 38596 106148 38652
rect 106084 38592 106148 38596
rect 106164 38652 106228 38656
rect 106164 38596 106168 38652
rect 106168 38596 106224 38652
rect 106224 38596 106228 38652
rect 106164 38592 106228 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 106660 38108 106724 38112
rect 106660 38052 106664 38108
rect 106664 38052 106720 38108
rect 106720 38052 106724 38108
rect 106660 38048 106724 38052
rect 106740 38108 106804 38112
rect 106740 38052 106744 38108
rect 106744 38052 106800 38108
rect 106800 38052 106804 38108
rect 106740 38048 106804 38052
rect 106820 38108 106884 38112
rect 106820 38052 106824 38108
rect 106824 38052 106880 38108
rect 106880 38052 106884 38108
rect 106820 38048 106884 38052
rect 106900 38108 106964 38112
rect 106900 38052 106904 38108
rect 106904 38052 106960 38108
rect 106960 38052 106964 38108
rect 106900 38048 106964 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 105924 37564 105988 37568
rect 105924 37508 105928 37564
rect 105928 37508 105984 37564
rect 105984 37508 105988 37564
rect 105924 37504 105988 37508
rect 106004 37564 106068 37568
rect 106004 37508 106008 37564
rect 106008 37508 106064 37564
rect 106064 37508 106068 37564
rect 106004 37504 106068 37508
rect 106084 37564 106148 37568
rect 106084 37508 106088 37564
rect 106088 37508 106144 37564
rect 106144 37508 106148 37564
rect 106084 37504 106148 37508
rect 106164 37564 106228 37568
rect 106164 37508 106168 37564
rect 106168 37508 106224 37564
rect 106224 37508 106228 37564
rect 106164 37504 106228 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 106660 37020 106724 37024
rect 106660 36964 106664 37020
rect 106664 36964 106720 37020
rect 106720 36964 106724 37020
rect 106660 36960 106724 36964
rect 106740 37020 106804 37024
rect 106740 36964 106744 37020
rect 106744 36964 106800 37020
rect 106800 36964 106804 37020
rect 106740 36960 106804 36964
rect 106820 37020 106884 37024
rect 106820 36964 106824 37020
rect 106824 36964 106880 37020
rect 106880 36964 106884 37020
rect 106820 36960 106884 36964
rect 106900 37020 106964 37024
rect 106900 36964 106904 37020
rect 106904 36964 106960 37020
rect 106960 36964 106964 37020
rect 106900 36960 106964 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 105924 36476 105988 36480
rect 105924 36420 105928 36476
rect 105928 36420 105984 36476
rect 105984 36420 105988 36476
rect 105924 36416 105988 36420
rect 106004 36476 106068 36480
rect 106004 36420 106008 36476
rect 106008 36420 106064 36476
rect 106064 36420 106068 36476
rect 106004 36416 106068 36420
rect 106084 36476 106148 36480
rect 106084 36420 106088 36476
rect 106088 36420 106144 36476
rect 106144 36420 106148 36476
rect 106084 36416 106148 36420
rect 106164 36476 106228 36480
rect 106164 36420 106168 36476
rect 106168 36420 106224 36476
rect 106224 36420 106228 36476
rect 106164 36416 106228 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 106660 35932 106724 35936
rect 106660 35876 106664 35932
rect 106664 35876 106720 35932
rect 106720 35876 106724 35932
rect 106660 35872 106724 35876
rect 106740 35932 106804 35936
rect 106740 35876 106744 35932
rect 106744 35876 106800 35932
rect 106800 35876 106804 35932
rect 106740 35872 106804 35876
rect 106820 35932 106884 35936
rect 106820 35876 106824 35932
rect 106824 35876 106880 35932
rect 106880 35876 106884 35932
rect 106820 35872 106884 35876
rect 106900 35932 106964 35936
rect 106900 35876 106904 35932
rect 106904 35876 106960 35932
rect 106960 35876 106964 35932
rect 106900 35872 106964 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 105924 35388 105988 35392
rect 105924 35332 105928 35388
rect 105928 35332 105984 35388
rect 105984 35332 105988 35388
rect 105924 35328 105988 35332
rect 106004 35388 106068 35392
rect 106004 35332 106008 35388
rect 106008 35332 106064 35388
rect 106064 35332 106068 35388
rect 106004 35328 106068 35332
rect 106084 35388 106148 35392
rect 106084 35332 106088 35388
rect 106088 35332 106144 35388
rect 106144 35332 106148 35388
rect 106084 35328 106148 35332
rect 106164 35388 106228 35392
rect 106164 35332 106168 35388
rect 106168 35332 106224 35388
rect 106224 35332 106228 35388
rect 106164 35328 106228 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 106660 34844 106724 34848
rect 106660 34788 106664 34844
rect 106664 34788 106720 34844
rect 106720 34788 106724 34844
rect 106660 34784 106724 34788
rect 106740 34844 106804 34848
rect 106740 34788 106744 34844
rect 106744 34788 106800 34844
rect 106800 34788 106804 34844
rect 106740 34784 106804 34788
rect 106820 34844 106884 34848
rect 106820 34788 106824 34844
rect 106824 34788 106880 34844
rect 106880 34788 106884 34844
rect 106820 34784 106884 34788
rect 106900 34844 106964 34848
rect 106900 34788 106904 34844
rect 106904 34788 106960 34844
rect 106960 34788 106964 34844
rect 106900 34784 106964 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 105924 34300 105988 34304
rect 105924 34244 105928 34300
rect 105928 34244 105984 34300
rect 105984 34244 105988 34300
rect 105924 34240 105988 34244
rect 106004 34300 106068 34304
rect 106004 34244 106008 34300
rect 106008 34244 106064 34300
rect 106064 34244 106068 34300
rect 106004 34240 106068 34244
rect 106084 34300 106148 34304
rect 106084 34244 106088 34300
rect 106088 34244 106144 34300
rect 106144 34244 106148 34300
rect 106084 34240 106148 34244
rect 106164 34300 106228 34304
rect 106164 34244 106168 34300
rect 106168 34244 106224 34300
rect 106224 34244 106228 34300
rect 106164 34240 106228 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 106660 33756 106724 33760
rect 106660 33700 106664 33756
rect 106664 33700 106720 33756
rect 106720 33700 106724 33756
rect 106660 33696 106724 33700
rect 106740 33756 106804 33760
rect 106740 33700 106744 33756
rect 106744 33700 106800 33756
rect 106800 33700 106804 33756
rect 106740 33696 106804 33700
rect 106820 33756 106884 33760
rect 106820 33700 106824 33756
rect 106824 33700 106880 33756
rect 106880 33700 106884 33756
rect 106820 33696 106884 33700
rect 106900 33756 106964 33760
rect 106900 33700 106904 33756
rect 106904 33700 106960 33756
rect 106960 33700 106964 33756
rect 106900 33696 106964 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 105924 33212 105988 33216
rect 105924 33156 105928 33212
rect 105928 33156 105984 33212
rect 105984 33156 105988 33212
rect 105924 33152 105988 33156
rect 106004 33212 106068 33216
rect 106004 33156 106008 33212
rect 106008 33156 106064 33212
rect 106064 33156 106068 33212
rect 106004 33152 106068 33156
rect 106084 33212 106148 33216
rect 106084 33156 106088 33212
rect 106088 33156 106144 33212
rect 106144 33156 106148 33212
rect 106084 33152 106148 33156
rect 106164 33212 106228 33216
rect 106164 33156 106168 33212
rect 106168 33156 106224 33212
rect 106224 33156 106228 33212
rect 106164 33152 106228 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 106660 32668 106724 32672
rect 106660 32612 106664 32668
rect 106664 32612 106720 32668
rect 106720 32612 106724 32668
rect 106660 32608 106724 32612
rect 106740 32668 106804 32672
rect 106740 32612 106744 32668
rect 106744 32612 106800 32668
rect 106800 32612 106804 32668
rect 106740 32608 106804 32612
rect 106820 32668 106884 32672
rect 106820 32612 106824 32668
rect 106824 32612 106880 32668
rect 106880 32612 106884 32668
rect 106820 32608 106884 32612
rect 106900 32668 106964 32672
rect 106900 32612 106904 32668
rect 106904 32612 106960 32668
rect 106960 32612 106964 32668
rect 106900 32608 106964 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 105924 32124 105988 32128
rect 105924 32068 105928 32124
rect 105928 32068 105984 32124
rect 105984 32068 105988 32124
rect 105924 32064 105988 32068
rect 106004 32124 106068 32128
rect 106004 32068 106008 32124
rect 106008 32068 106064 32124
rect 106064 32068 106068 32124
rect 106004 32064 106068 32068
rect 106084 32124 106148 32128
rect 106084 32068 106088 32124
rect 106088 32068 106144 32124
rect 106144 32068 106148 32124
rect 106084 32064 106148 32068
rect 106164 32124 106228 32128
rect 106164 32068 106168 32124
rect 106168 32068 106224 32124
rect 106224 32068 106228 32124
rect 106164 32064 106228 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 106660 31580 106724 31584
rect 106660 31524 106664 31580
rect 106664 31524 106720 31580
rect 106720 31524 106724 31580
rect 106660 31520 106724 31524
rect 106740 31580 106804 31584
rect 106740 31524 106744 31580
rect 106744 31524 106800 31580
rect 106800 31524 106804 31580
rect 106740 31520 106804 31524
rect 106820 31580 106884 31584
rect 106820 31524 106824 31580
rect 106824 31524 106880 31580
rect 106880 31524 106884 31580
rect 106820 31520 106884 31524
rect 106900 31580 106964 31584
rect 106900 31524 106904 31580
rect 106904 31524 106960 31580
rect 106960 31524 106964 31580
rect 106900 31520 106964 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 105924 31036 105988 31040
rect 105924 30980 105928 31036
rect 105928 30980 105984 31036
rect 105984 30980 105988 31036
rect 105924 30976 105988 30980
rect 106004 31036 106068 31040
rect 106004 30980 106008 31036
rect 106008 30980 106064 31036
rect 106064 30980 106068 31036
rect 106004 30976 106068 30980
rect 106084 31036 106148 31040
rect 106084 30980 106088 31036
rect 106088 30980 106144 31036
rect 106144 30980 106148 31036
rect 106084 30976 106148 30980
rect 106164 31036 106228 31040
rect 106164 30980 106168 31036
rect 106168 30980 106224 31036
rect 106224 30980 106228 31036
rect 106164 30976 106228 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 106660 30492 106724 30496
rect 106660 30436 106664 30492
rect 106664 30436 106720 30492
rect 106720 30436 106724 30492
rect 106660 30432 106724 30436
rect 106740 30492 106804 30496
rect 106740 30436 106744 30492
rect 106744 30436 106800 30492
rect 106800 30436 106804 30492
rect 106740 30432 106804 30436
rect 106820 30492 106884 30496
rect 106820 30436 106824 30492
rect 106824 30436 106880 30492
rect 106880 30436 106884 30492
rect 106820 30432 106884 30436
rect 106900 30492 106964 30496
rect 106900 30436 106904 30492
rect 106904 30436 106960 30492
rect 106960 30436 106964 30492
rect 106900 30432 106964 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 105924 29948 105988 29952
rect 105924 29892 105928 29948
rect 105928 29892 105984 29948
rect 105984 29892 105988 29948
rect 105924 29888 105988 29892
rect 106004 29948 106068 29952
rect 106004 29892 106008 29948
rect 106008 29892 106064 29948
rect 106064 29892 106068 29948
rect 106004 29888 106068 29892
rect 106084 29948 106148 29952
rect 106084 29892 106088 29948
rect 106088 29892 106144 29948
rect 106144 29892 106148 29948
rect 106084 29888 106148 29892
rect 106164 29948 106228 29952
rect 106164 29892 106168 29948
rect 106168 29892 106224 29948
rect 106224 29892 106228 29948
rect 106164 29888 106228 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 106660 29404 106724 29408
rect 106660 29348 106664 29404
rect 106664 29348 106720 29404
rect 106720 29348 106724 29404
rect 106660 29344 106724 29348
rect 106740 29404 106804 29408
rect 106740 29348 106744 29404
rect 106744 29348 106800 29404
rect 106800 29348 106804 29404
rect 106740 29344 106804 29348
rect 106820 29404 106884 29408
rect 106820 29348 106824 29404
rect 106824 29348 106880 29404
rect 106880 29348 106884 29404
rect 106820 29344 106884 29348
rect 106900 29404 106964 29408
rect 106900 29348 106904 29404
rect 106904 29348 106960 29404
rect 106960 29348 106964 29404
rect 106900 29344 106964 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 105924 28860 105988 28864
rect 105924 28804 105928 28860
rect 105928 28804 105984 28860
rect 105984 28804 105988 28860
rect 105924 28800 105988 28804
rect 106004 28860 106068 28864
rect 106004 28804 106008 28860
rect 106008 28804 106064 28860
rect 106064 28804 106068 28860
rect 106004 28800 106068 28804
rect 106084 28860 106148 28864
rect 106084 28804 106088 28860
rect 106088 28804 106144 28860
rect 106144 28804 106148 28860
rect 106084 28800 106148 28804
rect 106164 28860 106228 28864
rect 106164 28804 106168 28860
rect 106168 28804 106224 28860
rect 106224 28804 106228 28860
rect 106164 28800 106228 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 106660 28316 106724 28320
rect 106660 28260 106664 28316
rect 106664 28260 106720 28316
rect 106720 28260 106724 28316
rect 106660 28256 106724 28260
rect 106740 28316 106804 28320
rect 106740 28260 106744 28316
rect 106744 28260 106800 28316
rect 106800 28260 106804 28316
rect 106740 28256 106804 28260
rect 106820 28316 106884 28320
rect 106820 28260 106824 28316
rect 106824 28260 106880 28316
rect 106880 28260 106884 28316
rect 106820 28256 106884 28260
rect 106900 28316 106964 28320
rect 106900 28260 106904 28316
rect 106904 28260 106960 28316
rect 106960 28260 106964 28316
rect 106900 28256 106964 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 105924 27772 105988 27776
rect 105924 27716 105928 27772
rect 105928 27716 105984 27772
rect 105984 27716 105988 27772
rect 105924 27712 105988 27716
rect 106004 27772 106068 27776
rect 106004 27716 106008 27772
rect 106008 27716 106064 27772
rect 106064 27716 106068 27772
rect 106004 27712 106068 27716
rect 106084 27772 106148 27776
rect 106084 27716 106088 27772
rect 106088 27716 106144 27772
rect 106144 27716 106148 27772
rect 106084 27712 106148 27716
rect 106164 27772 106228 27776
rect 106164 27716 106168 27772
rect 106168 27716 106224 27772
rect 106224 27716 106228 27772
rect 106164 27712 106228 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 106660 27228 106724 27232
rect 106660 27172 106664 27228
rect 106664 27172 106720 27228
rect 106720 27172 106724 27228
rect 106660 27168 106724 27172
rect 106740 27228 106804 27232
rect 106740 27172 106744 27228
rect 106744 27172 106800 27228
rect 106800 27172 106804 27228
rect 106740 27168 106804 27172
rect 106820 27228 106884 27232
rect 106820 27172 106824 27228
rect 106824 27172 106880 27228
rect 106880 27172 106884 27228
rect 106820 27168 106884 27172
rect 106900 27228 106964 27232
rect 106900 27172 106904 27228
rect 106904 27172 106960 27228
rect 106960 27172 106964 27228
rect 106900 27168 106964 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 105924 26684 105988 26688
rect 105924 26628 105928 26684
rect 105928 26628 105984 26684
rect 105984 26628 105988 26684
rect 105924 26624 105988 26628
rect 106004 26684 106068 26688
rect 106004 26628 106008 26684
rect 106008 26628 106064 26684
rect 106064 26628 106068 26684
rect 106004 26624 106068 26628
rect 106084 26684 106148 26688
rect 106084 26628 106088 26684
rect 106088 26628 106144 26684
rect 106144 26628 106148 26684
rect 106084 26624 106148 26628
rect 106164 26684 106228 26688
rect 106164 26628 106168 26684
rect 106168 26628 106224 26684
rect 106224 26628 106228 26684
rect 106164 26624 106228 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 106660 26140 106724 26144
rect 106660 26084 106664 26140
rect 106664 26084 106720 26140
rect 106720 26084 106724 26140
rect 106660 26080 106724 26084
rect 106740 26140 106804 26144
rect 106740 26084 106744 26140
rect 106744 26084 106800 26140
rect 106800 26084 106804 26140
rect 106740 26080 106804 26084
rect 106820 26140 106884 26144
rect 106820 26084 106824 26140
rect 106824 26084 106880 26140
rect 106880 26084 106884 26140
rect 106820 26080 106884 26084
rect 106900 26140 106964 26144
rect 106900 26084 106904 26140
rect 106904 26084 106960 26140
rect 106960 26084 106964 26140
rect 106900 26080 106964 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 105924 25596 105988 25600
rect 105924 25540 105928 25596
rect 105928 25540 105984 25596
rect 105984 25540 105988 25596
rect 105924 25536 105988 25540
rect 106004 25596 106068 25600
rect 106004 25540 106008 25596
rect 106008 25540 106064 25596
rect 106064 25540 106068 25596
rect 106004 25536 106068 25540
rect 106084 25596 106148 25600
rect 106084 25540 106088 25596
rect 106088 25540 106144 25596
rect 106144 25540 106148 25596
rect 106084 25536 106148 25540
rect 106164 25596 106228 25600
rect 106164 25540 106168 25596
rect 106168 25540 106224 25596
rect 106224 25540 106228 25596
rect 106164 25536 106228 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 106660 25052 106724 25056
rect 106660 24996 106664 25052
rect 106664 24996 106720 25052
rect 106720 24996 106724 25052
rect 106660 24992 106724 24996
rect 106740 25052 106804 25056
rect 106740 24996 106744 25052
rect 106744 24996 106800 25052
rect 106800 24996 106804 25052
rect 106740 24992 106804 24996
rect 106820 25052 106884 25056
rect 106820 24996 106824 25052
rect 106824 24996 106880 25052
rect 106880 24996 106884 25052
rect 106820 24992 106884 24996
rect 106900 25052 106964 25056
rect 106900 24996 106904 25052
rect 106904 24996 106960 25052
rect 106960 24996 106964 25052
rect 106900 24992 106964 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 105924 24508 105988 24512
rect 105924 24452 105928 24508
rect 105928 24452 105984 24508
rect 105984 24452 105988 24508
rect 105924 24448 105988 24452
rect 106004 24508 106068 24512
rect 106004 24452 106008 24508
rect 106008 24452 106064 24508
rect 106064 24452 106068 24508
rect 106004 24448 106068 24452
rect 106084 24508 106148 24512
rect 106084 24452 106088 24508
rect 106088 24452 106144 24508
rect 106144 24452 106148 24508
rect 106084 24448 106148 24452
rect 106164 24508 106228 24512
rect 106164 24452 106168 24508
rect 106168 24452 106224 24508
rect 106224 24452 106228 24508
rect 106164 24448 106228 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 106660 23964 106724 23968
rect 106660 23908 106664 23964
rect 106664 23908 106720 23964
rect 106720 23908 106724 23964
rect 106660 23904 106724 23908
rect 106740 23964 106804 23968
rect 106740 23908 106744 23964
rect 106744 23908 106800 23964
rect 106800 23908 106804 23964
rect 106740 23904 106804 23908
rect 106820 23964 106884 23968
rect 106820 23908 106824 23964
rect 106824 23908 106880 23964
rect 106880 23908 106884 23964
rect 106820 23904 106884 23908
rect 106900 23964 106964 23968
rect 106900 23908 106904 23964
rect 106904 23908 106960 23964
rect 106960 23908 106964 23964
rect 106900 23904 106964 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 105924 23420 105988 23424
rect 105924 23364 105928 23420
rect 105928 23364 105984 23420
rect 105984 23364 105988 23420
rect 105924 23360 105988 23364
rect 106004 23420 106068 23424
rect 106004 23364 106008 23420
rect 106008 23364 106064 23420
rect 106064 23364 106068 23420
rect 106004 23360 106068 23364
rect 106084 23420 106148 23424
rect 106084 23364 106088 23420
rect 106088 23364 106144 23420
rect 106144 23364 106148 23420
rect 106084 23360 106148 23364
rect 106164 23420 106228 23424
rect 106164 23364 106168 23420
rect 106168 23364 106224 23420
rect 106224 23364 106228 23420
rect 106164 23360 106228 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 106660 22876 106724 22880
rect 106660 22820 106664 22876
rect 106664 22820 106720 22876
rect 106720 22820 106724 22876
rect 106660 22816 106724 22820
rect 106740 22876 106804 22880
rect 106740 22820 106744 22876
rect 106744 22820 106800 22876
rect 106800 22820 106804 22876
rect 106740 22816 106804 22820
rect 106820 22876 106884 22880
rect 106820 22820 106824 22876
rect 106824 22820 106880 22876
rect 106880 22820 106884 22876
rect 106820 22816 106884 22820
rect 106900 22876 106964 22880
rect 106900 22820 106904 22876
rect 106904 22820 106960 22876
rect 106960 22820 106964 22876
rect 106900 22816 106964 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 105924 22332 105988 22336
rect 105924 22276 105928 22332
rect 105928 22276 105984 22332
rect 105984 22276 105988 22332
rect 105924 22272 105988 22276
rect 106004 22332 106068 22336
rect 106004 22276 106008 22332
rect 106008 22276 106064 22332
rect 106064 22276 106068 22332
rect 106004 22272 106068 22276
rect 106084 22332 106148 22336
rect 106084 22276 106088 22332
rect 106088 22276 106144 22332
rect 106144 22276 106148 22332
rect 106084 22272 106148 22276
rect 106164 22332 106228 22336
rect 106164 22276 106168 22332
rect 106168 22276 106224 22332
rect 106224 22276 106228 22332
rect 106164 22272 106228 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 106660 21788 106724 21792
rect 106660 21732 106664 21788
rect 106664 21732 106720 21788
rect 106720 21732 106724 21788
rect 106660 21728 106724 21732
rect 106740 21788 106804 21792
rect 106740 21732 106744 21788
rect 106744 21732 106800 21788
rect 106800 21732 106804 21788
rect 106740 21728 106804 21732
rect 106820 21788 106884 21792
rect 106820 21732 106824 21788
rect 106824 21732 106880 21788
rect 106880 21732 106884 21788
rect 106820 21728 106884 21732
rect 106900 21788 106964 21792
rect 106900 21732 106904 21788
rect 106904 21732 106960 21788
rect 106960 21732 106964 21788
rect 106900 21728 106964 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 105924 21244 105988 21248
rect 105924 21188 105928 21244
rect 105928 21188 105984 21244
rect 105984 21188 105988 21244
rect 105924 21184 105988 21188
rect 106004 21244 106068 21248
rect 106004 21188 106008 21244
rect 106008 21188 106064 21244
rect 106064 21188 106068 21244
rect 106004 21184 106068 21188
rect 106084 21244 106148 21248
rect 106084 21188 106088 21244
rect 106088 21188 106144 21244
rect 106144 21188 106148 21244
rect 106084 21184 106148 21188
rect 106164 21244 106228 21248
rect 106164 21188 106168 21244
rect 106168 21188 106224 21244
rect 106224 21188 106228 21244
rect 106164 21184 106228 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 106660 20700 106724 20704
rect 106660 20644 106664 20700
rect 106664 20644 106720 20700
rect 106720 20644 106724 20700
rect 106660 20640 106724 20644
rect 106740 20700 106804 20704
rect 106740 20644 106744 20700
rect 106744 20644 106800 20700
rect 106800 20644 106804 20700
rect 106740 20640 106804 20644
rect 106820 20700 106884 20704
rect 106820 20644 106824 20700
rect 106824 20644 106880 20700
rect 106880 20644 106884 20700
rect 106820 20640 106884 20644
rect 106900 20700 106964 20704
rect 106900 20644 106904 20700
rect 106904 20644 106960 20700
rect 106960 20644 106964 20700
rect 106900 20640 106964 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 105924 20156 105988 20160
rect 105924 20100 105928 20156
rect 105928 20100 105984 20156
rect 105984 20100 105988 20156
rect 105924 20096 105988 20100
rect 106004 20156 106068 20160
rect 106004 20100 106008 20156
rect 106008 20100 106064 20156
rect 106064 20100 106068 20156
rect 106004 20096 106068 20100
rect 106084 20156 106148 20160
rect 106084 20100 106088 20156
rect 106088 20100 106144 20156
rect 106144 20100 106148 20156
rect 106084 20096 106148 20100
rect 106164 20156 106228 20160
rect 106164 20100 106168 20156
rect 106168 20100 106224 20156
rect 106224 20100 106228 20156
rect 106164 20096 106228 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 106660 19612 106724 19616
rect 106660 19556 106664 19612
rect 106664 19556 106720 19612
rect 106720 19556 106724 19612
rect 106660 19552 106724 19556
rect 106740 19612 106804 19616
rect 106740 19556 106744 19612
rect 106744 19556 106800 19612
rect 106800 19556 106804 19612
rect 106740 19552 106804 19556
rect 106820 19612 106884 19616
rect 106820 19556 106824 19612
rect 106824 19556 106880 19612
rect 106880 19556 106884 19612
rect 106820 19552 106884 19556
rect 106900 19612 106964 19616
rect 106900 19556 106904 19612
rect 106904 19556 106960 19612
rect 106960 19556 106964 19612
rect 106900 19552 106964 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 105924 19068 105988 19072
rect 105924 19012 105928 19068
rect 105928 19012 105984 19068
rect 105984 19012 105988 19068
rect 105924 19008 105988 19012
rect 106004 19068 106068 19072
rect 106004 19012 106008 19068
rect 106008 19012 106064 19068
rect 106064 19012 106068 19068
rect 106004 19008 106068 19012
rect 106084 19068 106148 19072
rect 106084 19012 106088 19068
rect 106088 19012 106144 19068
rect 106144 19012 106148 19068
rect 106084 19008 106148 19012
rect 106164 19068 106228 19072
rect 106164 19012 106168 19068
rect 106168 19012 106224 19068
rect 106224 19012 106228 19068
rect 106164 19008 106228 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 106660 18524 106724 18528
rect 106660 18468 106664 18524
rect 106664 18468 106720 18524
rect 106720 18468 106724 18524
rect 106660 18464 106724 18468
rect 106740 18524 106804 18528
rect 106740 18468 106744 18524
rect 106744 18468 106800 18524
rect 106800 18468 106804 18524
rect 106740 18464 106804 18468
rect 106820 18524 106884 18528
rect 106820 18468 106824 18524
rect 106824 18468 106880 18524
rect 106880 18468 106884 18524
rect 106820 18464 106884 18468
rect 106900 18524 106964 18528
rect 106900 18468 106904 18524
rect 106904 18468 106960 18524
rect 106960 18468 106964 18524
rect 106900 18464 106964 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 105924 17980 105988 17984
rect 105924 17924 105928 17980
rect 105928 17924 105984 17980
rect 105984 17924 105988 17980
rect 105924 17920 105988 17924
rect 106004 17980 106068 17984
rect 106004 17924 106008 17980
rect 106008 17924 106064 17980
rect 106064 17924 106068 17980
rect 106004 17920 106068 17924
rect 106084 17980 106148 17984
rect 106084 17924 106088 17980
rect 106088 17924 106144 17980
rect 106144 17924 106148 17980
rect 106084 17920 106148 17924
rect 106164 17980 106228 17984
rect 106164 17924 106168 17980
rect 106168 17924 106224 17980
rect 106224 17924 106228 17980
rect 106164 17920 106228 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 106660 17436 106724 17440
rect 106660 17380 106664 17436
rect 106664 17380 106720 17436
rect 106720 17380 106724 17436
rect 106660 17376 106724 17380
rect 106740 17436 106804 17440
rect 106740 17380 106744 17436
rect 106744 17380 106800 17436
rect 106800 17380 106804 17436
rect 106740 17376 106804 17380
rect 106820 17436 106884 17440
rect 106820 17380 106824 17436
rect 106824 17380 106880 17436
rect 106880 17380 106884 17436
rect 106820 17376 106884 17380
rect 106900 17436 106964 17440
rect 106900 17380 106904 17436
rect 106904 17380 106960 17436
rect 106960 17380 106964 17436
rect 106900 17376 106964 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 105924 16892 105988 16896
rect 105924 16836 105928 16892
rect 105928 16836 105984 16892
rect 105984 16836 105988 16892
rect 105924 16832 105988 16836
rect 106004 16892 106068 16896
rect 106004 16836 106008 16892
rect 106008 16836 106064 16892
rect 106064 16836 106068 16892
rect 106004 16832 106068 16836
rect 106084 16892 106148 16896
rect 106084 16836 106088 16892
rect 106088 16836 106144 16892
rect 106144 16836 106148 16892
rect 106084 16832 106148 16836
rect 106164 16892 106228 16896
rect 106164 16836 106168 16892
rect 106168 16836 106224 16892
rect 106224 16836 106228 16892
rect 106164 16832 106228 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 106660 16348 106724 16352
rect 106660 16292 106664 16348
rect 106664 16292 106720 16348
rect 106720 16292 106724 16348
rect 106660 16288 106724 16292
rect 106740 16348 106804 16352
rect 106740 16292 106744 16348
rect 106744 16292 106800 16348
rect 106800 16292 106804 16348
rect 106740 16288 106804 16292
rect 106820 16348 106884 16352
rect 106820 16292 106824 16348
rect 106824 16292 106880 16348
rect 106880 16292 106884 16348
rect 106820 16288 106884 16292
rect 106900 16348 106964 16352
rect 106900 16292 106904 16348
rect 106904 16292 106960 16348
rect 106960 16292 106964 16348
rect 106900 16288 106964 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 105924 15804 105988 15808
rect 105924 15748 105928 15804
rect 105928 15748 105984 15804
rect 105984 15748 105988 15804
rect 105924 15744 105988 15748
rect 106004 15804 106068 15808
rect 106004 15748 106008 15804
rect 106008 15748 106064 15804
rect 106064 15748 106068 15804
rect 106004 15744 106068 15748
rect 106084 15804 106148 15808
rect 106084 15748 106088 15804
rect 106088 15748 106144 15804
rect 106144 15748 106148 15804
rect 106084 15744 106148 15748
rect 106164 15804 106228 15808
rect 106164 15748 106168 15804
rect 106168 15748 106224 15804
rect 106224 15748 106228 15804
rect 106164 15744 106228 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 106660 15260 106724 15264
rect 106660 15204 106664 15260
rect 106664 15204 106720 15260
rect 106720 15204 106724 15260
rect 106660 15200 106724 15204
rect 106740 15260 106804 15264
rect 106740 15204 106744 15260
rect 106744 15204 106800 15260
rect 106800 15204 106804 15260
rect 106740 15200 106804 15204
rect 106820 15260 106884 15264
rect 106820 15204 106824 15260
rect 106824 15204 106880 15260
rect 106880 15204 106884 15260
rect 106820 15200 106884 15204
rect 106900 15260 106964 15264
rect 106900 15204 106904 15260
rect 106904 15204 106960 15260
rect 106960 15204 106964 15260
rect 106900 15200 106964 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 105924 14716 105988 14720
rect 105924 14660 105928 14716
rect 105928 14660 105984 14716
rect 105984 14660 105988 14716
rect 105924 14656 105988 14660
rect 106004 14716 106068 14720
rect 106004 14660 106008 14716
rect 106008 14660 106064 14716
rect 106064 14660 106068 14716
rect 106004 14656 106068 14660
rect 106084 14716 106148 14720
rect 106084 14660 106088 14716
rect 106088 14660 106144 14716
rect 106144 14660 106148 14716
rect 106084 14656 106148 14660
rect 106164 14716 106228 14720
rect 106164 14660 106168 14716
rect 106168 14660 106224 14716
rect 106224 14660 106228 14716
rect 106164 14656 106228 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 106660 14172 106724 14176
rect 106660 14116 106664 14172
rect 106664 14116 106720 14172
rect 106720 14116 106724 14172
rect 106660 14112 106724 14116
rect 106740 14172 106804 14176
rect 106740 14116 106744 14172
rect 106744 14116 106800 14172
rect 106800 14116 106804 14172
rect 106740 14112 106804 14116
rect 106820 14172 106884 14176
rect 106820 14116 106824 14172
rect 106824 14116 106880 14172
rect 106880 14116 106884 14172
rect 106820 14112 106884 14116
rect 106900 14172 106964 14176
rect 106900 14116 106904 14172
rect 106904 14116 106960 14172
rect 106960 14116 106964 14172
rect 106900 14112 106964 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 105924 13628 105988 13632
rect 105924 13572 105928 13628
rect 105928 13572 105984 13628
rect 105984 13572 105988 13628
rect 105924 13568 105988 13572
rect 106004 13628 106068 13632
rect 106004 13572 106008 13628
rect 106008 13572 106064 13628
rect 106064 13572 106068 13628
rect 106004 13568 106068 13572
rect 106084 13628 106148 13632
rect 106084 13572 106088 13628
rect 106088 13572 106144 13628
rect 106144 13572 106148 13628
rect 106084 13568 106148 13572
rect 106164 13628 106228 13632
rect 106164 13572 106168 13628
rect 106168 13572 106224 13628
rect 106224 13572 106228 13628
rect 106164 13568 106228 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 106660 13084 106724 13088
rect 106660 13028 106664 13084
rect 106664 13028 106720 13084
rect 106720 13028 106724 13084
rect 106660 13024 106724 13028
rect 106740 13084 106804 13088
rect 106740 13028 106744 13084
rect 106744 13028 106800 13084
rect 106800 13028 106804 13084
rect 106740 13024 106804 13028
rect 106820 13084 106884 13088
rect 106820 13028 106824 13084
rect 106824 13028 106880 13084
rect 106880 13028 106884 13084
rect 106820 13024 106884 13028
rect 106900 13084 106964 13088
rect 106900 13028 106904 13084
rect 106904 13028 106960 13084
rect 106960 13028 106964 13084
rect 106900 13024 106964 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 105924 12540 105988 12544
rect 105924 12484 105928 12540
rect 105928 12484 105984 12540
rect 105984 12484 105988 12540
rect 105924 12480 105988 12484
rect 106004 12540 106068 12544
rect 106004 12484 106008 12540
rect 106008 12484 106064 12540
rect 106064 12484 106068 12540
rect 106004 12480 106068 12484
rect 106084 12540 106148 12544
rect 106084 12484 106088 12540
rect 106088 12484 106144 12540
rect 106144 12484 106148 12540
rect 106084 12480 106148 12484
rect 106164 12540 106228 12544
rect 106164 12484 106168 12540
rect 106168 12484 106224 12540
rect 106224 12484 106228 12540
rect 106164 12480 106228 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 106660 11996 106724 12000
rect 106660 11940 106664 11996
rect 106664 11940 106720 11996
rect 106720 11940 106724 11996
rect 106660 11936 106724 11940
rect 106740 11996 106804 12000
rect 106740 11940 106744 11996
rect 106744 11940 106800 11996
rect 106800 11940 106804 11996
rect 106740 11936 106804 11940
rect 106820 11996 106884 12000
rect 106820 11940 106824 11996
rect 106824 11940 106880 11996
rect 106880 11940 106884 11996
rect 106820 11936 106884 11940
rect 106900 11996 106964 12000
rect 106900 11940 106904 11996
rect 106904 11940 106960 11996
rect 106960 11940 106964 11996
rect 106900 11936 106964 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 105924 11452 105988 11456
rect 105924 11396 105928 11452
rect 105928 11396 105984 11452
rect 105984 11396 105988 11452
rect 105924 11392 105988 11396
rect 106004 11452 106068 11456
rect 106004 11396 106008 11452
rect 106008 11396 106064 11452
rect 106064 11396 106068 11452
rect 106004 11392 106068 11396
rect 106084 11452 106148 11456
rect 106084 11396 106088 11452
rect 106088 11396 106144 11452
rect 106144 11396 106148 11452
rect 106084 11392 106148 11396
rect 106164 11452 106228 11456
rect 106164 11396 106168 11452
rect 106168 11396 106224 11452
rect 106224 11396 106228 11452
rect 106164 11392 106228 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 106660 10908 106724 10912
rect 106660 10852 106664 10908
rect 106664 10852 106720 10908
rect 106720 10852 106724 10908
rect 106660 10848 106724 10852
rect 106740 10908 106804 10912
rect 106740 10852 106744 10908
rect 106744 10852 106800 10908
rect 106800 10852 106804 10908
rect 106740 10848 106804 10852
rect 106820 10908 106884 10912
rect 106820 10852 106824 10908
rect 106824 10852 106880 10908
rect 106880 10852 106884 10908
rect 106820 10848 106884 10852
rect 106900 10908 106964 10912
rect 106900 10852 106904 10908
rect 106904 10852 106960 10908
rect 106960 10852 106964 10908
rect 106900 10848 106964 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 105924 10364 105988 10368
rect 105924 10308 105928 10364
rect 105928 10308 105984 10364
rect 105984 10308 105988 10364
rect 105924 10304 105988 10308
rect 106004 10364 106068 10368
rect 106004 10308 106008 10364
rect 106008 10308 106064 10364
rect 106064 10308 106068 10364
rect 106004 10304 106068 10308
rect 106084 10364 106148 10368
rect 106084 10308 106088 10364
rect 106088 10308 106144 10364
rect 106144 10308 106148 10364
rect 106084 10304 106148 10308
rect 106164 10364 106228 10368
rect 106164 10308 106168 10364
rect 106168 10308 106224 10364
rect 106224 10308 106228 10364
rect 106164 10304 106228 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 106660 9820 106724 9824
rect 106660 9764 106664 9820
rect 106664 9764 106720 9820
rect 106720 9764 106724 9820
rect 106660 9760 106724 9764
rect 106740 9820 106804 9824
rect 106740 9764 106744 9820
rect 106744 9764 106800 9820
rect 106800 9764 106804 9820
rect 106740 9760 106804 9764
rect 106820 9820 106884 9824
rect 106820 9764 106824 9820
rect 106824 9764 106880 9820
rect 106880 9764 106884 9820
rect 106820 9760 106884 9764
rect 106900 9820 106964 9824
rect 106900 9764 106904 9820
rect 106904 9764 106960 9820
rect 106960 9764 106964 9820
rect 106900 9760 106964 9764
rect 23438 9752 23502 9756
rect 23438 9696 23478 9752
rect 23478 9696 23502 9752
rect 23438 9692 23502 9696
rect 25774 9752 25838 9756
rect 25774 9696 25778 9752
rect 25778 9696 25834 9752
rect 25834 9696 25838 9752
rect 25774 9692 25838 9696
rect 28120 9752 28184 9756
rect 28120 9696 28170 9752
rect 28170 9696 28184 9752
rect 28120 9692 28184 9696
rect 29278 9692 29342 9756
rect 30446 9752 30510 9756
rect 30446 9696 30470 9752
rect 30470 9696 30510 9752
rect 30446 9692 30510 9696
rect 90527 9752 90591 9756
rect 90527 9696 90546 9752
rect 90546 9696 90591 9752
rect 90527 9692 90591 9696
rect 90956 9752 91020 9756
rect 90956 9696 90970 9752
rect 90970 9696 91020 9752
rect 90956 9692 91020 9696
rect 16058 9616 16122 9620
rect 16058 9560 16082 9616
rect 16082 9560 16122 9616
rect 16058 9556 16122 9560
rect 24624 9616 24688 9620
rect 24624 9560 24674 9616
rect 24674 9560 24688 9616
rect 24624 9556 24688 9560
rect 90680 9616 90744 9620
rect 90680 9560 90730 9616
rect 90730 9560 90744 9616
rect 90680 9556 90744 9560
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 105924 9276 105988 9280
rect 105924 9220 105928 9276
rect 105928 9220 105984 9276
rect 105984 9220 105988 9276
rect 105924 9216 105988 9220
rect 106004 9276 106068 9280
rect 106004 9220 106008 9276
rect 106008 9220 106064 9276
rect 106064 9220 106068 9276
rect 106004 9216 106068 9220
rect 106084 9276 106148 9280
rect 106084 9220 106088 9276
rect 106088 9220 106144 9276
rect 106144 9220 106148 9276
rect 106084 9216 106148 9220
rect 106164 9276 106228 9280
rect 106164 9220 106168 9276
rect 106168 9220 106224 9276
rect 106224 9220 106228 9276
rect 106164 9216 106228 9220
rect 26924 8876 26988 8940
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 106660 8732 106724 8736
rect 106660 8676 106664 8732
rect 106664 8676 106720 8732
rect 106720 8676 106724 8732
rect 106660 8672 106724 8676
rect 106740 8732 106804 8736
rect 106740 8676 106744 8732
rect 106744 8676 106800 8732
rect 106800 8676 106804 8732
rect 106740 8672 106804 8676
rect 106820 8732 106884 8736
rect 106820 8676 106824 8732
rect 106824 8676 106880 8732
rect 106880 8676 106884 8732
rect 106820 8672 106884 8676
rect 106900 8732 106964 8736
rect 106900 8676 106904 8732
rect 106904 8676 106960 8732
rect 106960 8676 106964 8732
rect 106900 8672 106964 8676
rect 31708 8256 31772 8260
rect 31708 8200 31722 8256
rect 31722 8200 31772 8256
rect 31708 8196 31772 8200
rect 32812 8196 32876 8260
rect 33916 8196 33980 8260
rect 35204 8196 35268 8260
rect 36308 8256 36372 8260
rect 36308 8200 36358 8256
rect 36358 8200 36372 8256
rect 36308 8196 36372 8200
rect 37412 8256 37476 8260
rect 37412 8200 37462 8256
rect 37462 8200 37476 8256
rect 37412 8196 37476 8200
rect 38700 8256 38764 8260
rect 38700 8200 38750 8256
rect 38750 8200 38764 8256
rect 38700 8196 38764 8200
rect 40908 8196 40972 8260
rect 42196 8256 42260 8260
rect 42196 8200 42210 8256
rect 42210 8200 42260 8256
rect 42196 8196 42260 8200
rect 43300 8196 43364 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 105924 8188 105988 8192
rect 105924 8132 105928 8188
rect 105928 8132 105984 8188
rect 105984 8132 105988 8188
rect 105924 8128 105988 8132
rect 106004 8188 106068 8192
rect 106004 8132 106008 8188
rect 106008 8132 106064 8188
rect 106064 8132 106068 8188
rect 106004 8128 106068 8132
rect 106084 8188 106148 8192
rect 106084 8132 106088 8188
rect 106088 8132 106144 8188
rect 106144 8132 106148 8188
rect 106084 8128 106148 8132
rect 106164 8188 106228 8192
rect 106164 8132 106168 8188
rect 106168 8132 106224 8188
rect 106224 8132 106228 8188
rect 106164 8128 106228 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 66316 7644 66380 7648
rect 66316 7588 66320 7644
rect 66320 7588 66376 7644
rect 66376 7588 66380 7644
rect 66316 7584 66380 7588
rect 66396 7644 66460 7648
rect 66396 7588 66400 7644
rect 66400 7588 66456 7644
rect 66456 7588 66460 7644
rect 66396 7584 66460 7588
rect 66476 7644 66540 7648
rect 66476 7588 66480 7644
rect 66480 7588 66536 7644
rect 66536 7588 66540 7644
rect 66476 7584 66540 7588
rect 66556 7644 66620 7648
rect 66556 7588 66560 7644
rect 66560 7588 66616 7644
rect 66616 7588 66620 7644
rect 66556 7584 66620 7588
rect 97036 7644 97100 7648
rect 97036 7588 97040 7644
rect 97040 7588 97096 7644
rect 97096 7588 97100 7644
rect 97036 7584 97100 7588
rect 97116 7644 97180 7648
rect 97116 7588 97120 7644
rect 97120 7588 97176 7644
rect 97176 7588 97180 7644
rect 97116 7584 97180 7588
rect 97196 7644 97260 7648
rect 97196 7588 97200 7644
rect 97200 7588 97256 7644
rect 97256 7588 97260 7644
rect 97196 7584 97260 7588
rect 97276 7644 97340 7648
rect 97276 7588 97280 7644
rect 97280 7588 97336 7644
rect 97336 7588 97340 7644
rect 97276 7584 97340 7588
rect 106660 7644 106724 7648
rect 106660 7588 106664 7644
rect 106664 7588 106720 7644
rect 106720 7588 106724 7644
rect 106660 7584 106724 7588
rect 106740 7644 106804 7648
rect 106740 7588 106744 7644
rect 106744 7588 106800 7644
rect 106800 7588 106804 7644
rect 106740 7584 106804 7588
rect 106820 7644 106884 7648
rect 106820 7588 106824 7644
rect 106824 7588 106880 7644
rect 106880 7588 106884 7644
rect 106820 7584 106884 7588
rect 106900 7644 106964 7648
rect 106900 7588 106904 7644
rect 106904 7588 106960 7644
rect 106960 7588 106964 7644
rect 106900 7584 106964 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 96376 7100 96440 7104
rect 96376 7044 96380 7100
rect 96380 7044 96436 7100
rect 96436 7044 96440 7100
rect 96376 7040 96440 7044
rect 96456 7100 96520 7104
rect 96456 7044 96460 7100
rect 96460 7044 96516 7100
rect 96516 7044 96520 7100
rect 96456 7040 96520 7044
rect 96536 7100 96600 7104
rect 96536 7044 96540 7100
rect 96540 7044 96596 7100
rect 96596 7044 96600 7100
rect 96536 7040 96600 7044
rect 96616 7100 96680 7104
rect 96616 7044 96620 7100
rect 96620 7044 96676 7100
rect 96676 7044 96680 7100
rect 96616 7040 96680 7044
rect 105924 7100 105988 7104
rect 105924 7044 105928 7100
rect 105928 7044 105984 7100
rect 105984 7044 105988 7100
rect 105924 7040 105988 7044
rect 106004 7100 106068 7104
rect 106004 7044 106008 7100
rect 106008 7044 106064 7100
rect 106064 7044 106068 7100
rect 106004 7040 106068 7044
rect 106084 7100 106148 7104
rect 106084 7044 106088 7100
rect 106088 7044 106144 7100
rect 106144 7044 106148 7100
rect 106084 7040 106148 7044
rect 106164 7100 106228 7104
rect 106164 7044 106168 7100
rect 106168 7044 106224 7100
rect 106224 7044 106228 7100
rect 106164 7040 106228 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 66316 6556 66380 6560
rect 66316 6500 66320 6556
rect 66320 6500 66376 6556
rect 66376 6500 66380 6556
rect 66316 6496 66380 6500
rect 66396 6556 66460 6560
rect 66396 6500 66400 6556
rect 66400 6500 66456 6556
rect 66456 6500 66460 6556
rect 66396 6496 66460 6500
rect 66476 6556 66540 6560
rect 66476 6500 66480 6556
rect 66480 6500 66536 6556
rect 66536 6500 66540 6556
rect 66476 6496 66540 6500
rect 66556 6556 66620 6560
rect 66556 6500 66560 6556
rect 66560 6500 66616 6556
rect 66616 6500 66620 6556
rect 66556 6496 66620 6500
rect 97036 6556 97100 6560
rect 97036 6500 97040 6556
rect 97040 6500 97096 6556
rect 97096 6500 97100 6556
rect 97036 6496 97100 6500
rect 97116 6556 97180 6560
rect 97116 6500 97120 6556
rect 97120 6500 97176 6556
rect 97176 6500 97180 6556
rect 97116 6496 97180 6500
rect 97196 6556 97260 6560
rect 97196 6500 97200 6556
rect 97200 6500 97256 6556
rect 97256 6500 97260 6556
rect 97196 6496 97260 6500
rect 97276 6556 97340 6560
rect 97276 6500 97280 6556
rect 97280 6500 97336 6556
rect 97336 6500 97340 6556
rect 97276 6496 97340 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 96376 6012 96440 6016
rect 96376 5956 96380 6012
rect 96380 5956 96436 6012
rect 96436 5956 96440 6012
rect 96376 5952 96440 5956
rect 96456 6012 96520 6016
rect 96456 5956 96460 6012
rect 96460 5956 96516 6012
rect 96516 5956 96520 6012
rect 96456 5952 96520 5956
rect 96536 6012 96600 6016
rect 96536 5956 96540 6012
rect 96540 5956 96596 6012
rect 96596 5956 96600 6012
rect 96536 5952 96600 5956
rect 96616 6012 96680 6016
rect 96616 5956 96620 6012
rect 96620 5956 96676 6012
rect 96676 5956 96680 6012
rect 96616 5952 96680 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 66316 5468 66380 5472
rect 66316 5412 66320 5468
rect 66320 5412 66376 5468
rect 66376 5412 66380 5468
rect 66316 5408 66380 5412
rect 66396 5468 66460 5472
rect 66396 5412 66400 5468
rect 66400 5412 66456 5468
rect 66456 5412 66460 5468
rect 66396 5408 66460 5412
rect 66476 5468 66540 5472
rect 66476 5412 66480 5468
rect 66480 5412 66536 5468
rect 66536 5412 66540 5468
rect 66476 5408 66540 5412
rect 66556 5468 66620 5472
rect 66556 5412 66560 5468
rect 66560 5412 66616 5468
rect 66616 5412 66620 5468
rect 66556 5408 66620 5412
rect 97036 5468 97100 5472
rect 97036 5412 97040 5468
rect 97040 5412 97096 5468
rect 97096 5412 97100 5468
rect 97036 5408 97100 5412
rect 97116 5468 97180 5472
rect 97116 5412 97120 5468
rect 97120 5412 97176 5468
rect 97176 5412 97180 5468
rect 97116 5408 97180 5412
rect 97196 5468 97260 5472
rect 97196 5412 97200 5468
rect 97200 5412 97256 5468
rect 97256 5412 97260 5468
rect 97196 5408 97260 5412
rect 97276 5468 97340 5472
rect 97276 5412 97280 5468
rect 97280 5412 97336 5468
rect 97336 5412 97340 5468
rect 97276 5408 97340 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 96376 4924 96440 4928
rect 96376 4868 96380 4924
rect 96380 4868 96436 4924
rect 96436 4868 96440 4924
rect 96376 4864 96440 4868
rect 96456 4924 96520 4928
rect 96456 4868 96460 4924
rect 96460 4868 96516 4924
rect 96516 4868 96520 4924
rect 96456 4864 96520 4868
rect 96536 4924 96600 4928
rect 96536 4868 96540 4924
rect 96540 4868 96596 4924
rect 96596 4868 96600 4924
rect 96536 4864 96600 4868
rect 96616 4924 96680 4928
rect 96616 4868 96620 4924
rect 96620 4868 96676 4924
rect 96676 4868 96680 4924
rect 96616 4864 96680 4868
rect 39804 4524 39868 4588
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 66316 4380 66380 4384
rect 66316 4324 66320 4380
rect 66320 4324 66376 4380
rect 66376 4324 66380 4380
rect 66316 4320 66380 4324
rect 66396 4380 66460 4384
rect 66396 4324 66400 4380
rect 66400 4324 66456 4380
rect 66456 4324 66460 4380
rect 66396 4320 66460 4324
rect 66476 4380 66540 4384
rect 66476 4324 66480 4380
rect 66480 4324 66536 4380
rect 66536 4324 66540 4380
rect 66476 4320 66540 4324
rect 66556 4380 66620 4384
rect 66556 4324 66560 4380
rect 66560 4324 66616 4380
rect 66616 4324 66620 4380
rect 66556 4320 66620 4324
rect 97036 4380 97100 4384
rect 97036 4324 97040 4380
rect 97040 4324 97096 4380
rect 97096 4324 97100 4380
rect 97036 4320 97100 4324
rect 97116 4380 97180 4384
rect 97116 4324 97120 4380
rect 97120 4324 97176 4380
rect 97176 4324 97180 4380
rect 97116 4320 97180 4324
rect 97196 4380 97260 4384
rect 97196 4324 97200 4380
rect 97200 4324 97256 4380
rect 97256 4324 97260 4380
rect 97196 4320 97260 4324
rect 97276 4380 97340 4384
rect 97276 4324 97280 4380
rect 97280 4324 97336 4380
rect 97336 4324 97340 4380
rect 97276 4320 97340 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 96376 3836 96440 3840
rect 96376 3780 96380 3836
rect 96380 3780 96436 3836
rect 96436 3780 96440 3836
rect 96376 3776 96440 3780
rect 96456 3836 96520 3840
rect 96456 3780 96460 3836
rect 96460 3780 96516 3836
rect 96516 3780 96520 3836
rect 96456 3776 96520 3780
rect 96536 3836 96600 3840
rect 96536 3780 96540 3836
rect 96540 3780 96596 3836
rect 96596 3780 96600 3836
rect 96536 3776 96600 3780
rect 96616 3836 96680 3840
rect 96616 3780 96620 3836
rect 96620 3780 96676 3836
rect 96676 3780 96680 3836
rect 96616 3776 96680 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 66316 3292 66380 3296
rect 66316 3236 66320 3292
rect 66320 3236 66376 3292
rect 66376 3236 66380 3292
rect 66316 3232 66380 3236
rect 66396 3292 66460 3296
rect 66396 3236 66400 3292
rect 66400 3236 66456 3292
rect 66456 3236 66460 3292
rect 66396 3232 66460 3236
rect 66476 3292 66540 3296
rect 66476 3236 66480 3292
rect 66480 3236 66536 3292
rect 66536 3236 66540 3292
rect 66476 3232 66540 3236
rect 66556 3292 66620 3296
rect 66556 3236 66560 3292
rect 66560 3236 66616 3292
rect 66616 3236 66620 3292
rect 66556 3232 66620 3236
rect 97036 3292 97100 3296
rect 97036 3236 97040 3292
rect 97040 3236 97096 3292
rect 97096 3236 97100 3292
rect 97036 3232 97100 3236
rect 97116 3292 97180 3296
rect 97116 3236 97120 3292
rect 97120 3236 97176 3292
rect 97176 3236 97180 3292
rect 97116 3232 97180 3236
rect 97196 3292 97260 3296
rect 97196 3236 97200 3292
rect 97200 3236 97256 3292
rect 97256 3236 97260 3292
rect 97196 3232 97260 3236
rect 97276 3292 97340 3296
rect 97276 3236 97280 3292
rect 97280 3236 97336 3292
rect 97336 3236 97340 3292
rect 97276 3232 97340 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 96376 2748 96440 2752
rect 96376 2692 96380 2748
rect 96380 2692 96436 2748
rect 96436 2692 96440 2748
rect 96376 2688 96440 2692
rect 96456 2748 96520 2752
rect 96456 2692 96460 2748
rect 96460 2692 96516 2748
rect 96516 2692 96520 2748
rect 96456 2688 96520 2692
rect 96536 2748 96600 2752
rect 96536 2692 96540 2748
rect 96540 2692 96596 2748
rect 96596 2692 96600 2748
rect 96536 2688 96600 2692
rect 96616 2748 96680 2752
rect 96616 2692 96620 2748
rect 96620 2692 96676 2748
rect 96676 2692 96680 2748
rect 96616 2688 96680 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
rect 66316 2204 66380 2208
rect 66316 2148 66320 2204
rect 66320 2148 66376 2204
rect 66376 2148 66380 2204
rect 66316 2144 66380 2148
rect 66396 2204 66460 2208
rect 66396 2148 66400 2204
rect 66400 2148 66456 2204
rect 66456 2148 66460 2204
rect 66396 2144 66460 2148
rect 66476 2204 66540 2208
rect 66476 2148 66480 2204
rect 66480 2148 66536 2204
rect 66536 2148 66540 2204
rect 66476 2144 66540 2148
rect 66556 2204 66620 2208
rect 66556 2148 66560 2204
rect 66560 2148 66616 2204
rect 66616 2148 66620 2204
rect 66556 2144 66620 2148
rect 97036 2204 97100 2208
rect 97036 2148 97040 2204
rect 97040 2148 97096 2204
rect 97096 2148 97100 2204
rect 97036 2144 97100 2148
rect 97116 2204 97180 2208
rect 97116 2148 97120 2204
rect 97120 2148 97176 2204
rect 97176 2148 97180 2204
rect 97116 2144 97180 2148
rect 97196 2204 97260 2208
rect 97196 2148 97200 2204
rect 97200 2148 97256 2204
rect 97256 2148 97260 2204
rect 97196 2144 97260 2148
rect 97276 2204 97340 2208
rect 97276 2148 97280 2204
rect 97280 2148 97336 2204
rect 97336 2148 97340 2204
rect 97276 2144 97340 2148
<< metal4 >>
rect 4208 147456 4528 147472
rect 4208 147392 4216 147456
rect 4280 147392 4296 147456
rect 4360 147392 4376 147456
rect 4440 147392 4456 147456
rect 4520 147392 4528 147456
rect 4208 146368 4528 147392
rect 4208 146304 4216 146368
rect 4280 146304 4296 146368
rect 4360 146304 4376 146368
rect 4440 146304 4456 146368
rect 4520 146304 4528 146368
rect 4208 145280 4528 146304
rect 4208 145216 4216 145280
rect 4280 145216 4296 145280
rect 4360 145216 4376 145280
rect 4440 145216 4456 145280
rect 4520 145216 4528 145280
rect 4208 144192 4528 145216
rect 4208 144128 4216 144192
rect 4280 144128 4296 144192
rect 4360 144128 4376 144192
rect 4440 144128 4456 144192
rect 4520 144128 4528 144192
rect 4208 143104 4528 144128
rect 4208 143040 4216 143104
rect 4280 143040 4296 143104
rect 4360 143040 4376 143104
rect 4440 143040 4456 143104
rect 4520 143040 4528 143104
rect 4208 142016 4528 143040
rect 4208 141952 4216 142016
rect 4280 141952 4296 142016
rect 4360 141952 4376 142016
rect 4440 141952 4456 142016
rect 4520 141952 4528 142016
rect 4208 141218 4528 141952
rect 4208 140982 4250 141218
rect 4486 140982 4528 141218
rect 4208 140928 4528 140982
rect 4208 140864 4216 140928
rect 4280 140864 4296 140928
rect 4360 140864 4376 140928
rect 4440 140864 4456 140928
rect 4520 140864 4528 140928
rect 4208 139840 4528 140864
rect 4208 139776 4216 139840
rect 4280 139776 4296 139840
rect 4360 139776 4376 139840
rect 4440 139776 4456 139840
rect 4520 139776 4528 139840
rect 4208 138752 4528 139776
rect 4208 138688 4216 138752
rect 4280 138688 4296 138752
rect 4360 138688 4376 138752
rect 4440 138688 4456 138752
rect 4520 138688 4528 138752
rect 4208 137664 4528 138688
rect 4208 137600 4216 137664
rect 4280 137600 4296 137664
rect 4360 137600 4376 137664
rect 4440 137600 4456 137664
rect 4520 137600 4528 137664
rect 4208 136576 4528 137600
rect 4208 136512 4216 136576
rect 4280 136512 4296 136576
rect 4360 136512 4376 136576
rect 4440 136512 4456 136576
rect 4520 136512 4528 136576
rect 4208 135488 4528 136512
rect 4208 135424 4216 135488
rect 4280 135424 4296 135488
rect 4360 135424 4376 135488
rect 4440 135424 4456 135488
rect 4520 135424 4528 135488
rect 4208 134400 4528 135424
rect 4208 134336 4216 134400
rect 4280 134336 4296 134400
rect 4360 134336 4376 134400
rect 4440 134336 4456 134400
rect 4520 134336 4528 134400
rect 4208 133312 4528 134336
rect 4208 133248 4216 133312
rect 4280 133248 4296 133312
rect 4360 133248 4376 133312
rect 4440 133248 4456 133312
rect 4520 133248 4528 133312
rect 4208 132224 4528 133248
rect 4208 132160 4216 132224
rect 4280 132160 4296 132224
rect 4360 132160 4376 132224
rect 4440 132160 4456 132224
rect 4520 132160 4528 132224
rect 4208 131136 4528 132160
rect 4208 131072 4216 131136
rect 4280 131072 4296 131136
rect 4360 131072 4376 131136
rect 4440 131072 4456 131136
rect 4520 131072 4528 131136
rect 4208 130048 4528 131072
rect 4208 129984 4216 130048
rect 4280 129984 4296 130048
rect 4360 129984 4376 130048
rect 4440 129984 4456 130048
rect 4520 129984 4528 130048
rect 4208 128960 4528 129984
rect 4208 128896 4216 128960
rect 4280 128896 4296 128960
rect 4360 128896 4376 128960
rect 4440 128896 4456 128960
rect 4520 128896 4528 128960
rect 4208 128168 4528 128896
rect 4208 127932 4250 128168
rect 4486 127932 4528 128168
rect 4208 127872 4528 127932
rect 4208 127808 4216 127872
rect 4280 127808 4296 127872
rect 4360 127808 4376 127872
rect 4440 127808 4456 127872
rect 4520 127808 4528 127872
rect 4208 126784 4528 127808
rect 4208 126720 4216 126784
rect 4280 126720 4296 126784
rect 4360 126720 4376 126784
rect 4440 126720 4456 126784
rect 4520 126720 4528 126784
rect 4208 125696 4528 126720
rect 4208 125632 4216 125696
rect 4280 125632 4296 125696
rect 4360 125632 4376 125696
rect 4440 125632 4456 125696
rect 4520 125632 4528 125696
rect 4208 124608 4528 125632
rect 4208 124544 4216 124608
rect 4280 124544 4296 124608
rect 4360 124544 4376 124608
rect 4440 124544 4456 124608
rect 4520 124544 4528 124608
rect 4208 123520 4528 124544
rect 4208 123456 4216 123520
rect 4280 123456 4296 123520
rect 4360 123456 4376 123520
rect 4440 123456 4456 123520
rect 4520 123456 4528 123520
rect 4208 122432 4528 123456
rect 4208 122368 4216 122432
rect 4280 122368 4296 122432
rect 4360 122368 4376 122432
rect 4440 122368 4456 122432
rect 4520 122368 4528 122432
rect 4208 121344 4528 122368
rect 4208 121280 4216 121344
rect 4280 121280 4296 121344
rect 4360 121280 4376 121344
rect 4440 121280 4456 121344
rect 4520 121280 4528 121344
rect 4208 120256 4528 121280
rect 4208 120192 4216 120256
rect 4280 120192 4296 120256
rect 4360 120192 4376 120256
rect 4440 120192 4456 120256
rect 4520 120192 4528 120256
rect 4208 119168 4528 120192
rect 4208 119104 4216 119168
rect 4280 119104 4296 119168
rect 4360 119104 4376 119168
rect 4440 119104 4456 119168
rect 4520 119104 4528 119168
rect 4208 118080 4528 119104
rect 4208 118016 4216 118080
rect 4280 118016 4296 118080
rect 4360 118016 4376 118080
rect 4440 118016 4456 118080
rect 4520 118016 4528 118080
rect 4208 116992 4528 118016
rect 4208 116928 4216 116992
rect 4280 116928 4296 116992
rect 4360 116928 4376 116992
rect 4440 116928 4456 116992
rect 4520 116928 4528 116992
rect 4208 115904 4528 116928
rect 4208 115840 4216 115904
rect 4280 115840 4296 115904
rect 4360 115840 4376 115904
rect 4440 115840 4456 115904
rect 4520 115840 4528 115904
rect 4208 114816 4528 115840
rect 4208 114752 4216 114816
rect 4280 114752 4296 114816
rect 4360 114752 4376 114816
rect 4440 114752 4456 114816
rect 4520 114752 4528 114816
rect 4208 113728 4528 114752
rect 4208 113664 4216 113728
rect 4280 113664 4296 113728
rect 4360 113664 4376 113728
rect 4440 113664 4456 113728
rect 4520 113664 4528 113728
rect 4208 112640 4528 113664
rect 4208 112576 4216 112640
rect 4280 112576 4296 112640
rect 4360 112576 4376 112640
rect 4440 112576 4456 112640
rect 4520 112576 4528 112640
rect 4208 111552 4528 112576
rect 4208 111488 4216 111552
rect 4280 111488 4296 111552
rect 4360 111488 4376 111552
rect 4440 111488 4456 111552
rect 4520 111488 4528 111552
rect 4208 110464 4528 111488
rect 4208 110400 4216 110464
rect 4280 110400 4296 110464
rect 4360 110400 4376 110464
rect 4440 110400 4456 110464
rect 4520 110400 4528 110464
rect 4208 109376 4528 110400
rect 4208 109312 4216 109376
rect 4280 109312 4296 109376
rect 4360 109312 4376 109376
rect 4440 109312 4456 109376
rect 4520 109312 4528 109376
rect 4208 108288 4528 109312
rect 4208 108224 4216 108288
rect 4280 108224 4296 108288
rect 4360 108224 4376 108288
rect 4440 108224 4456 108288
rect 4520 108224 4528 108288
rect 4208 107200 4528 108224
rect 4208 107136 4216 107200
rect 4280 107136 4296 107200
rect 4360 107136 4376 107200
rect 4440 107136 4456 107200
rect 4520 107136 4528 107200
rect 4208 106112 4528 107136
rect 4208 106048 4216 106112
rect 4280 106048 4296 106112
rect 4360 106048 4376 106112
rect 4440 106048 4456 106112
rect 4520 106048 4528 106112
rect 4208 105024 4528 106048
rect 4208 104960 4216 105024
rect 4280 104960 4296 105024
rect 4360 104960 4376 105024
rect 4440 104960 4456 105024
rect 4520 104960 4528 105024
rect 4208 103936 4528 104960
rect 4208 103872 4216 103936
rect 4280 103872 4296 103936
rect 4360 103872 4376 103936
rect 4440 103872 4456 103936
rect 4520 103872 4528 103936
rect 4208 102848 4528 103872
rect 4208 102784 4216 102848
rect 4280 102784 4296 102848
rect 4360 102784 4376 102848
rect 4440 102784 4456 102848
rect 4520 102784 4528 102848
rect 4208 101760 4528 102784
rect 4208 101696 4216 101760
rect 4280 101696 4296 101760
rect 4360 101696 4376 101760
rect 4440 101696 4456 101760
rect 4520 101696 4528 101760
rect 4208 100672 4528 101696
rect 4208 100608 4216 100672
rect 4280 100608 4296 100672
rect 4360 100608 4376 100672
rect 4440 100608 4456 100672
rect 4520 100608 4528 100672
rect 4208 99584 4528 100608
rect 4208 99520 4216 99584
rect 4280 99520 4296 99584
rect 4360 99520 4376 99584
rect 4440 99520 4456 99584
rect 4520 99520 4528 99584
rect 4208 98496 4528 99520
rect 4208 98432 4216 98496
rect 4280 98432 4296 98496
rect 4360 98432 4376 98496
rect 4440 98432 4456 98496
rect 4520 98432 4528 98496
rect 4208 97532 4528 98432
rect 4208 97408 4250 97532
rect 4486 97408 4528 97532
rect 4208 97344 4216 97408
rect 4520 97344 4528 97408
rect 4208 97296 4250 97344
rect 4486 97296 4528 97344
rect 4208 96320 4528 97296
rect 4208 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4528 96320
rect 4208 95232 4528 96256
rect 4208 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4528 95232
rect 4208 94144 4528 95168
rect 4208 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4528 94144
rect 4208 93056 4528 94080
rect 4208 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4528 93056
rect 4208 91968 4528 92992
rect 4208 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4528 91968
rect 4208 90880 4528 91904
rect 4208 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4528 90880
rect 4208 89792 4528 90816
rect 4208 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4528 89792
rect 4208 88704 4528 89728
rect 4208 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4528 88704
rect 4208 87616 4528 88640
rect 4208 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4528 87616
rect 4208 86528 4528 87552
rect 4208 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4528 86528
rect 4208 85440 4528 86464
rect 4208 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4528 85440
rect 4208 84352 4528 85376
rect 4208 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4528 84352
rect 4208 83264 4528 84288
rect 4208 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4528 83264
rect 4208 82176 4528 83200
rect 4208 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4528 82176
rect 4208 81088 4528 82112
rect 4208 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4528 81088
rect 4208 80000 4528 81024
rect 4208 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4528 80000
rect 4208 78912 4528 79936
rect 4208 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4528 78912
rect 4208 77824 4528 78848
rect 4208 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4528 77824
rect 4208 76736 4528 77760
rect 4208 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4528 76736
rect 4208 75648 4528 76672
rect 4208 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4528 75648
rect 4208 74560 4528 75584
rect 4208 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4528 74560
rect 4208 73472 4528 74496
rect 4208 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4528 73472
rect 4208 72384 4528 73408
rect 4208 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4528 72384
rect 4208 71296 4528 72320
rect 4208 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4528 71296
rect 4208 70208 4528 71232
rect 4208 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4528 70208
rect 4208 69120 4528 70144
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66896 4296 66944
rect 4360 66896 4376 66944
rect 4440 66896 4456 66944
rect 4520 66880 4528 66944
rect 4208 66660 4250 66880
rect 4486 66660 4528 66880
rect 4208 65856 4528 66660
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 146912 5188 147472
rect 4868 146848 4876 146912
rect 4940 146848 4956 146912
rect 5020 146848 5036 146912
rect 5100 146848 5116 146912
rect 5180 146848 5188 146912
rect 4868 145824 5188 146848
rect 4868 145760 4876 145824
rect 4940 145760 4956 145824
rect 5020 145760 5036 145824
rect 5100 145760 5116 145824
rect 5180 145760 5188 145824
rect 4868 144736 5188 145760
rect 4868 144672 4876 144736
rect 4940 144672 4956 144736
rect 5020 144672 5036 144736
rect 5100 144672 5116 144736
rect 5180 144672 5188 144736
rect 4868 143648 5188 144672
rect 4868 143584 4876 143648
rect 4940 143584 4956 143648
rect 5020 143584 5036 143648
rect 5100 143584 5116 143648
rect 5180 143584 5188 143648
rect 4868 142560 5188 143584
rect 4868 142496 4876 142560
rect 4940 142496 4956 142560
rect 5020 142496 5036 142560
rect 5100 142496 5116 142560
rect 5180 142496 5188 142560
rect 4868 141898 5188 142496
rect 4868 141662 4910 141898
rect 5146 141662 5188 141898
rect 4868 141472 5188 141662
rect 4868 141408 4876 141472
rect 4940 141408 4956 141472
rect 5020 141408 5036 141472
rect 5100 141408 5116 141472
rect 5180 141408 5188 141472
rect 4868 140384 5188 141408
rect 4868 140320 4876 140384
rect 4940 140320 4956 140384
rect 5020 140320 5036 140384
rect 5100 140320 5116 140384
rect 5180 140320 5188 140384
rect 4868 139296 5188 140320
rect 4868 139232 4876 139296
rect 4940 139232 4956 139296
rect 5020 139232 5036 139296
rect 5100 139232 5116 139296
rect 5180 139232 5188 139296
rect 4868 138208 5188 139232
rect 4868 138144 4876 138208
rect 4940 138144 4956 138208
rect 5020 138144 5036 138208
rect 5100 138144 5116 138208
rect 5180 138144 5188 138208
rect 4868 137120 5188 138144
rect 4868 137056 4876 137120
rect 4940 137056 4956 137120
rect 5020 137056 5036 137120
rect 5100 137056 5116 137120
rect 5180 137056 5188 137120
rect 4868 136032 5188 137056
rect 4868 135968 4876 136032
rect 4940 135968 4956 136032
rect 5020 135968 5036 136032
rect 5100 135968 5116 136032
rect 5180 135968 5188 136032
rect 4868 134944 5188 135968
rect 34928 147456 35248 147472
rect 34928 147392 34936 147456
rect 35000 147392 35016 147456
rect 35080 147392 35096 147456
rect 35160 147392 35176 147456
rect 35240 147392 35248 147456
rect 34928 146368 35248 147392
rect 34928 146304 34936 146368
rect 35000 146304 35016 146368
rect 35080 146304 35096 146368
rect 35160 146304 35176 146368
rect 35240 146304 35248 146368
rect 34928 145280 35248 146304
rect 34928 145216 34936 145280
rect 35000 145216 35016 145280
rect 35080 145216 35096 145280
rect 35160 145216 35176 145280
rect 35240 145216 35248 145280
rect 34928 144192 35248 145216
rect 34928 144128 34936 144192
rect 35000 144128 35016 144192
rect 35080 144128 35096 144192
rect 35160 144128 35176 144192
rect 35240 144128 35248 144192
rect 34928 143104 35248 144128
rect 34928 143040 34936 143104
rect 35000 143040 35016 143104
rect 35080 143040 35096 143104
rect 35160 143040 35176 143104
rect 35240 143040 35248 143104
rect 34928 142016 35248 143040
rect 34928 141952 34936 142016
rect 35000 141952 35016 142016
rect 35080 141952 35096 142016
rect 35160 141952 35176 142016
rect 35240 141952 35248 142016
rect 34928 141218 35248 141952
rect 34928 140982 34970 141218
rect 35206 140982 35248 141218
rect 34928 140928 35248 140982
rect 34928 140864 34936 140928
rect 35000 140864 35016 140928
rect 35080 140864 35096 140928
rect 35160 140864 35176 140928
rect 35240 140864 35248 140928
rect 34928 139840 35248 140864
rect 34928 139776 34936 139840
rect 35000 139776 35016 139840
rect 35080 139776 35096 139840
rect 35160 139776 35176 139840
rect 35240 139776 35248 139840
rect 34928 138752 35248 139776
rect 34928 138688 34936 138752
rect 35000 138688 35016 138752
rect 35080 138688 35096 138752
rect 35160 138688 35176 138752
rect 35240 138688 35248 138752
rect 34928 137664 35248 138688
rect 34928 137600 34936 137664
rect 35000 137600 35016 137664
rect 35080 137600 35096 137664
rect 35160 137600 35176 137664
rect 35240 137600 35248 137664
rect 34928 136576 35248 137600
rect 34928 136512 34936 136576
rect 35000 136512 35016 136576
rect 35080 136512 35096 136576
rect 35160 136512 35176 136576
rect 35240 136512 35248 136576
rect 34928 135650 35248 136512
rect 35588 146912 35908 147472
rect 35588 146848 35596 146912
rect 35660 146848 35676 146912
rect 35740 146848 35756 146912
rect 35820 146848 35836 146912
rect 35900 146848 35908 146912
rect 35588 145824 35908 146848
rect 35588 145760 35596 145824
rect 35660 145760 35676 145824
rect 35740 145760 35756 145824
rect 35820 145760 35836 145824
rect 35900 145760 35908 145824
rect 35588 144736 35908 145760
rect 35588 144672 35596 144736
rect 35660 144672 35676 144736
rect 35740 144672 35756 144736
rect 35820 144672 35836 144736
rect 35900 144672 35908 144736
rect 35588 143648 35908 144672
rect 35588 143584 35596 143648
rect 35660 143584 35676 143648
rect 35740 143584 35756 143648
rect 35820 143584 35836 143648
rect 35900 143584 35908 143648
rect 35588 142560 35908 143584
rect 35588 142496 35596 142560
rect 35660 142496 35676 142560
rect 35740 142496 35756 142560
rect 35820 142496 35836 142560
rect 35900 142496 35908 142560
rect 35588 141898 35908 142496
rect 35588 141662 35630 141898
rect 35866 141662 35908 141898
rect 35588 141472 35908 141662
rect 35588 141408 35596 141472
rect 35660 141408 35676 141472
rect 35740 141408 35756 141472
rect 35820 141408 35836 141472
rect 35900 141408 35908 141472
rect 35588 140384 35908 141408
rect 35588 140320 35596 140384
rect 35660 140320 35676 140384
rect 35740 140320 35756 140384
rect 35820 140320 35836 140384
rect 35900 140320 35908 140384
rect 35588 139296 35908 140320
rect 35588 139232 35596 139296
rect 35660 139232 35676 139296
rect 35740 139232 35756 139296
rect 35820 139232 35836 139296
rect 35900 139232 35908 139296
rect 35588 138208 35908 139232
rect 35588 138144 35596 138208
rect 35660 138144 35676 138208
rect 35740 138144 35756 138208
rect 35820 138144 35836 138208
rect 35900 138144 35908 138208
rect 35588 137120 35908 138144
rect 35588 137056 35596 137120
rect 35660 137056 35676 137120
rect 35740 137056 35756 137120
rect 35820 137056 35836 137120
rect 35900 137056 35908 137120
rect 35588 136032 35908 137056
rect 35588 135968 35596 136032
rect 35660 135968 35676 136032
rect 35740 135968 35756 136032
rect 35820 135968 35836 136032
rect 35900 135968 35908 136032
rect 35588 135650 35908 135968
rect 65648 147456 65968 147472
rect 65648 147392 65656 147456
rect 65720 147392 65736 147456
rect 65800 147392 65816 147456
rect 65880 147392 65896 147456
rect 65960 147392 65968 147456
rect 65648 146368 65968 147392
rect 65648 146304 65656 146368
rect 65720 146304 65736 146368
rect 65800 146304 65816 146368
rect 65880 146304 65896 146368
rect 65960 146304 65968 146368
rect 65648 145280 65968 146304
rect 65648 145216 65656 145280
rect 65720 145216 65736 145280
rect 65800 145216 65816 145280
rect 65880 145216 65896 145280
rect 65960 145216 65968 145280
rect 65648 144192 65968 145216
rect 65648 144128 65656 144192
rect 65720 144128 65736 144192
rect 65800 144128 65816 144192
rect 65880 144128 65896 144192
rect 65960 144128 65968 144192
rect 65648 143104 65968 144128
rect 65648 143040 65656 143104
rect 65720 143040 65736 143104
rect 65800 143040 65816 143104
rect 65880 143040 65896 143104
rect 65960 143040 65968 143104
rect 65648 142016 65968 143040
rect 65648 141952 65656 142016
rect 65720 141952 65736 142016
rect 65800 141952 65816 142016
rect 65880 141952 65896 142016
rect 65960 141952 65968 142016
rect 65648 141218 65968 141952
rect 65648 140982 65690 141218
rect 65926 140982 65968 141218
rect 65648 140928 65968 140982
rect 65648 140864 65656 140928
rect 65720 140864 65736 140928
rect 65800 140864 65816 140928
rect 65880 140864 65896 140928
rect 65960 140864 65968 140928
rect 65648 139840 65968 140864
rect 65648 139776 65656 139840
rect 65720 139776 65736 139840
rect 65800 139776 65816 139840
rect 65880 139776 65896 139840
rect 65960 139776 65968 139840
rect 65648 138752 65968 139776
rect 65648 138688 65656 138752
rect 65720 138688 65736 138752
rect 65800 138688 65816 138752
rect 65880 138688 65896 138752
rect 65960 138688 65968 138752
rect 65648 137664 65968 138688
rect 65648 137600 65656 137664
rect 65720 137600 65736 137664
rect 65800 137600 65816 137664
rect 65880 137600 65896 137664
rect 65960 137600 65968 137664
rect 65648 136576 65968 137600
rect 65648 136512 65656 136576
rect 65720 136512 65736 136576
rect 65800 136512 65816 136576
rect 65880 136512 65896 136576
rect 65960 136512 65968 136576
rect 65648 135834 65968 136512
rect 66308 146912 66628 147472
rect 66308 146848 66316 146912
rect 66380 146848 66396 146912
rect 66460 146848 66476 146912
rect 66540 146848 66556 146912
rect 66620 146848 66628 146912
rect 66308 145824 66628 146848
rect 66308 145760 66316 145824
rect 66380 145760 66396 145824
rect 66460 145760 66476 145824
rect 66540 145760 66556 145824
rect 66620 145760 66628 145824
rect 66308 144736 66628 145760
rect 66308 144672 66316 144736
rect 66380 144672 66396 144736
rect 66460 144672 66476 144736
rect 66540 144672 66556 144736
rect 66620 144672 66628 144736
rect 66308 143648 66628 144672
rect 66308 143584 66316 143648
rect 66380 143584 66396 143648
rect 66460 143584 66476 143648
rect 66540 143584 66556 143648
rect 66620 143584 66628 143648
rect 66308 142560 66628 143584
rect 66308 142496 66316 142560
rect 66380 142496 66396 142560
rect 66460 142496 66476 142560
rect 66540 142496 66556 142560
rect 66620 142496 66628 142560
rect 66308 141898 66628 142496
rect 66308 141662 66350 141898
rect 66586 141662 66628 141898
rect 66308 141472 66628 141662
rect 66308 141408 66316 141472
rect 66380 141408 66396 141472
rect 66460 141408 66476 141472
rect 66540 141408 66556 141472
rect 66620 141408 66628 141472
rect 66308 140384 66628 141408
rect 66308 140320 66316 140384
rect 66380 140320 66396 140384
rect 66460 140320 66476 140384
rect 66540 140320 66556 140384
rect 66620 140320 66628 140384
rect 66308 139296 66628 140320
rect 66308 139232 66316 139296
rect 66380 139232 66396 139296
rect 66460 139232 66476 139296
rect 66540 139232 66556 139296
rect 66620 139232 66628 139296
rect 66308 138208 66628 139232
rect 66308 138144 66316 138208
rect 66380 138144 66396 138208
rect 66460 138144 66476 138208
rect 66540 138144 66556 138208
rect 66620 138144 66628 138208
rect 66308 137120 66628 138144
rect 66308 137056 66316 137120
rect 66380 137056 66396 137120
rect 66460 137056 66476 137120
rect 66540 137056 66556 137120
rect 66620 137056 66628 137120
rect 66308 136032 66628 137056
rect 66308 135968 66316 136032
rect 66380 135968 66396 136032
rect 66460 135968 66476 136032
rect 66540 135968 66556 136032
rect 66620 135968 66628 136032
rect 66308 135650 66628 135968
rect 96368 147456 96688 147472
rect 96368 147392 96376 147456
rect 96440 147392 96456 147456
rect 96520 147392 96536 147456
rect 96600 147392 96616 147456
rect 96680 147392 96688 147456
rect 96368 146368 96688 147392
rect 96368 146304 96376 146368
rect 96440 146304 96456 146368
rect 96520 146304 96536 146368
rect 96600 146304 96616 146368
rect 96680 146304 96688 146368
rect 96368 145280 96688 146304
rect 96368 145216 96376 145280
rect 96440 145216 96456 145280
rect 96520 145216 96536 145280
rect 96600 145216 96616 145280
rect 96680 145216 96688 145280
rect 96368 144192 96688 145216
rect 96368 144128 96376 144192
rect 96440 144128 96456 144192
rect 96520 144128 96536 144192
rect 96600 144128 96616 144192
rect 96680 144128 96688 144192
rect 96368 143104 96688 144128
rect 96368 143040 96376 143104
rect 96440 143040 96456 143104
rect 96520 143040 96536 143104
rect 96600 143040 96616 143104
rect 96680 143040 96688 143104
rect 96368 142016 96688 143040
rect 96368 141952 96376 142016
rect 96440 141952 96456 142016
rect 96520 141952 96536 142016
rect 96600 141952 96616 142016
rect 96680 141952 96688 142016
rect 96368 141218 96688 141952
rect 96368 140982 96410 141218
rect 96646 140982 96688 141218
rect 96368 140928 96688 140982
rect 96368 140864 96376 140928
rect 96440 140864 96456 140928
rect 96520 140864 96536 140928
rect 96600 140864 96616 140928
rect 96680 140864 96688 140928
rect 96368 139840 96688 140864
rect 96368 139776 96376 139840
rect 96440 139776 96456 139840
rect 96520 139776 96536 139840
rect 96600 139776 96616 139840
rect 96680 139776 96688 139840
rect 96368 138752 96688 139776
rect 96368 138688 96376 138752
rect 96440 138688 96456 138752
rect 96520 138688 96536 138752
rect 96600 138688 96616 138752
rect 96680 138688 96688 138752
rect 96368 137664 96688 138688
rect 96368 137600 96376 137664
rect 96440 137600 96456 137664
rect 96520 137600 96536 137664
rect 96600 137600 96616 137664
rect 96680 137600 96688 137664
rect 96368 136576 96688 137600
rect 96368 136512 96376 136576
rect 96440 136512 96456 136576
rect 96520 136512 96536 136576
rect 96600 136512 96616 136576
rect 96680 136512 96688 136576
rect 96368 135650 96688 136512
rect 97028 146912 97348 147472
rect 97028 146848 97036 146912
rect 97100 146848 97116 146912
rect 97180 146848 97196 146912
rect 97260 146848 97276 146912
rect 97340 146848 97348 146912
rect 97028 145824 97348 146848
rect 97028 145760 97036 145824
rect 97100 145760 97116 145824
rect 97180 145760 97196 145824
rect 97260 145760 97276 145824
rect 97340 145760 97348 145824
rect 97028 144736 97348 145760
rect 97028 144672 97036 144736
rect 97100 144672 97116 144736
rect 97180 144672 97196 144736
rect 97260 144672 97276 144736
rect 97340 144672 97348 144736
rect 97028 143648 97348 144672
rect 97028 143584 97036 143648
rect 97100 143584 97116 143648
rect 97180 143584 97196 143648
rect 97260 143584 97276 143648
rect 97340 143584 97348 143648
rect 97028 142560 97348 143584
rect 97028 142496 97036 142560
rect 97100 142496 97116 142560
rect 97180 142496 97196 142560
rect 97260 142496 97276 142560
rect 97340 142496 97348 142560
rect 97028 141898 97348 142496
rect 97028 141662 97070 141898
rect 97306 141662 97348 141898
rect 97028 141472 97348 141662
rect 97028 141408 97036 141472
rect 97100 141408 97116 141472
rect 97180 141408 97196 141472
rect 97260 141408 97276 141472
rect 97340 141408 97348 141472
rect 97028 140384 97348 141408
rect 97028 140320 97036 140384
rect 97100 140320 97116 140384
rect 97180 140320 97196 140384
rect 97260 140320 97276 140384
rect 97340 140320 97348 140384
rect 97028 139296 97348 140320
rect 97028 139232 97036 139296
rect 97100 139232 97116 139296
rect 97180 139232 97196 139296
rect 97260 139232 97276 139296
rect 97340 139232 97348 139296
rect 97028 138208 97348 139232
rect 97028 138144 97036 138208
rect 97100 138144 97116 138208
rect 97180 138144 97196 138208
rect 97260 138144 97276 138208
rect 97340 138144 97348 138208
rect 97028 137120 97348 138144
rect 97028 137056 97036 137120
rect 97100 137056 97116 137120
rect 97180 137056 97196 137120
rect 97260 137056 97276 137120
rect 97340 137056 97348 137120
rect 97028 136032 97348 137056
rect 97028 135968 97036 136032
rect 97100 135968 97116 136032
rect 97180 135968 97196 136032
rect 97260 135968 97276 136032
rect 97340 135968 97348 136032
rect 97028 135650 97348 135968
rect 105916 136576 106236 136592
rect 105916 136512 105924 136576
rect 105988 136512 106004 136576
rect 106068 136512 106084 136576
rect 106148 136512 106164 136576
rect 106228 136512 106236 136576
rect 105916 135488 106236 136512
rect 105916 135424 105924 135488
rect 105988 135424 106004 135488
rect 106068 135424 106084 135488
rect 106148 135424 106164 135488
rect 106228 135424 106236 135488
rect 58571 135284 58637 135285
rect 58571 135220 58572 135284
rect 58636 135220 58637 135284
rect 58571 135219 58637 135220
rect 61147 135284 61213 135285
rect 61147 135220 61148 135284
rect 61212 135220 61213 135284
rect 61147 135219 61213 135220
rect 66115 135284 66181 135285
rect 66115 135220 66116 135284
rect 66180 135220 66181 135284
rect 66115 135219 66181 135220
rect 68507 135284 68573 135285
rect 68507 135220 68508 135284
rect 68572 135220 68573 135284
rect 68507 135219 68573 135220
rect 71083 135284 71149 135285
rect 71083 135220 71084 135284
rect 71148 135220 71149 135284
rect 71083 135219 71149 135220
rect 4868 134880 4876 134944
rect 4940 134880 4956 134944
rect 5020 134880 5036 134944
rect 5100 134880 5116 134944
rect 5180 134880 5188 134944
rect 4868 133856 5188 134880
rect 58574 134330 58634 135219
rect 61150 134330 61210 135219
rect 63539 135148 63605 135149
rect 63539 135084 63540 135148
rect 63604 135084 63605 135148
rect 63539 135083 63605 135084
rect 58541 134270 58634 134330
rect 61058 134270 61210 134330
rect 38570 134196 38636 134197
rect 38570 134132 38571 134196
rect 38635 134132 38636 134196
rect 38570 134131 38636 134132
rect 41066 134196 41132 134197
rect 41066 134132 41067 134196
rect 41131 134132 41132 134196
rect 41066 134131 41132 134132
rect 51050 134196 51116 134197
rect 51050 134132 51051 134196
rect 51115 134132 51116 134196
rect 51050 134131 51116 134132
rect 56042 134196 56108 134197
rect 56042 134132 56043 134196
rect 56107 134132 56108 134196
rect 56042 134131 56108 134132
rect 36074 133924 36140 133925
rect 36074 133860 36075 133924
rect 36139 133860 36140 133924
rect 36074 133859 36140 133860
rect 4868 133792 4876 133856
rect 4940 133792 4956 133856
rect 5020 133792 5036 133856
rect 5100 133792 5116 133856
rect 5180 133792 5188 133856
rect 4868 132768 5188 133792
rect 36077 133676 36137 133859
rect 38573 133676 38633 134131
rect 41069 133676 41129 134131
rect 43562 133924 43628 133925
rect 43562 133860 43563 133924
rect 43627 133860 43628 133924
rect 43562 133859 43628 133860
rect 46058 133924 46124 133925
rect 46058 133860 46059 133924
rect 46123 133860 46124 133924
rect 46058 133859 46124 133860
rect 48543 133924 48609 133925
rect 48543 133860 48544 133924
rect 48608 133860 48609 133924
rect 48543 133859 48609 133860
rect 43565 133676 43625 133859
rect 46061 133676 46121 133859
rect 48546 133676 48606 133859
rect 51053 133676 51113 134131
rect 53546 134060 53612 134061
rect 53546 133996 53547 134060
rect 53611 133996 53612 134060
rect 53546 133995 53612 133996
rect 53549 133676 53609 133995
rect 56045 133676 56105 134131
rect 58541 133676 58601 134270
rect 61058 133676 61118 134270
rect 63542 133676 63602 135083
rect 66118 134330 66178 135219
rect 66029 134270 66178 134330
rect 66029 133676 66089 134270
rect 68510 133676 68570 135219
rect 71086 134330 71146 135219
rect 95923 134468 95989 134469
rect 95923 134404 95924 134468
rect 95988 134404 95989 134468
rect 95923 134403 95989 134404
rect 95926 134330 95986 134403
rect 71021 134270 71146 134330
rect 95860 134270 95986 134330
rect 105916 134400 106236 135424
rect 105916 134336 105924 134400
rect 105988 134336 106004 134400
rect 106068 134336 106084 134400
rect 106148 134336 106164 134400
rect 106228 134336 106236 134400
rect 71021 133676 71081 134270
rect 73514 134196 73580 134197
rect 73514 134132 73515 134196
rect 73579 134132 73580 134196
rect 73514 134131 73580 134132
rect 73517 133676 73577 134131
rect 86141 133924 86207 133925
rect 86141 133860 86142 133924
rect 86206 133860 86207 133924
rect 86141 133859 86207 133860
rect 87309 133924 87375 133925
rect 87309 133860 87310 133924
rect 87374 133860 87375 133924
rect 87309 133859 87375 133860
rect 86144 133676 86204 133859
rect 87312 133676 87372 133859
rect 95860 133676 95920 134270
rect 4868 132704 4876 132768
rect 4940 132704 4956 132768
rect 5020 132704 5036 132768
rect 5100 132704 5116 132768
rect 5180 132704 5188 132768
rect 4868 131680 5188 132704
rect 4868 131616 4876 131680
rect 4940 131616 4956 131680
rect 5020 131616 5036 131680
rect 5100 131616 5116 131680
rect 5180 131616 5188 131680
rect 4868 130592 5188 131616
rect 4868 130528 4876 130592
rect 4940 130528 4956 130592
rect 5020 130528 5036 130592
rect 5100 130528 5116 130592
rect 5180 130528 5188 130592
rect 4868 129504 5188 130528
rect 4868 129440 4876 129504
rect 4940 129440 4956 129504
rect 5020 129440 5036 129504
rect 5100 129440 5116 129504
rect 5180 129440 5188 129504
rect 4868 128828 5188 129440
rect 105916 133312 106236 134336
rect 105916 133248 105924 133312
rect 105988 133248 106004 133312
rect 106068 133248 106084 133312
rect 106148 133248 106164 133312
rect 106228 133248 106236 133312
rect 105916 132224 106236 133248
rect 105916 132160 105924 132224
rect 105988 132160 106004 132224
rect 106068 132160 106084 132224
rect 106148 132160 106164 132224
rect 106228 132160 106236 132224
rect 105916 131136 106236 132160
rect 105916 131072 105924 131136
rect 105988 131072 106004 131136
rect 106068 131072 106084 131136
rect 106148 131072 106164 131136
rect 106228 131072 106236 131136
rect 105916 130048 106236 131072
rect 105916 129984 105924 130048
rect 105988 129984 106004 130048
rect 106068 129984 106084 130048
rect 106148 129984 106164 130048
rect 106228 129984 106236 130048
rect 105916 128960 106236 129984
rect 105916 128896 105924 128960
rect 105988 128896 106004 128960
rect 106068 128896 106084 128960
rect 106148 128896 106164 128960
rect 106228 128896 106236 128960
rect 4868 128592 4910 128828
rect 5146 128592 5188 128828
rect 4868 128416 5188 128592
rect 10696 128828 11044 128870
rect 10696 128592 10752 128828
rect 10988 128592 11044 128828
rect 10696 128550 11044 128592
rect 100936 128828 101284 128870
rect 100936 128592 100992 128828
rect 101228 128592 101284 128828
rect 100936 128550 101284 128592
rect 4868 128352 4876 128416
rect 4940 128352 4956 128416
rect 5020 128352 5036 128416
rect 5100 128352 5116 128416
rect 5180 128352 5188 128416
rect 4868 127328 5188 128352
rect 10000 128168 10348 128210
rect 10000 127932 10056 128168
rect 10292 127932 10348 128168
rect 10000 127890 10348 127932
rect 101632 128168 101980 128210
rect 101632 127932 101688 128168
rect 101924 127932 101980 128168
rect 101632 127890 101980 127932
rect 105916 128168 106236 128896
rect 105916 127932 105958 128168
rect 106194 127932 106236 128168
rect 4868 127264 4876 127328
rect 4940 127264 4956 127328
rect 5020 127264 5036 127328
rect 5100 127264 5116 127328
rect 5180 127264 5188 127328
rect 4868 126240 5188 127264
rect 4868 126176 4876 126240
rect 4940 126176 4956 126240
rect 5020 126176 5036 126240
rect 5100 126176 5116 126240
rect 5180 126176 5188 126240
rect 4868 125152 5188 126176
rect 4868 125088 4876 125152
rect 4940 125088 4956 125152
rect 5020 125088 5036 125152
rect 5100 125088 5116 125152
rect 5180 125088 5188 125152
rect 4868 124064 5188 125088
rect 4868 124000 4876 124064
rect 4940 124000 4956 124064
rect 5020 124000 5036 124064
rect 5100 124000 5116 124064
rect 5180 124000 5188 124064
rect 4868 122976 5188 124000
rect 4868 122912 4876 122976
rect 4940 122912 4956 122976
rect 5020 122912 5036 122976
rect 5100 122912 5116 122976
rect 5180 122912 5188 122976
rect 4868 121888 5188 122912
rect 4868 121824 4876 121888
rect 4940 121824 4956 121888
rect 5020 121824 5036 121888
rect 5100 121824 5116 121888
rect 5180 121824 5188 121888
rect 4868 120800 5188 121824
rect 4868 120736 4876 120800
rect 4940 120736 4956 120800
rect 5020 120736 5036 120800
rect 5100 120736 5116 120800
rect 5180 120736 5188 120800
rect 4868 119712 5188 120736
rect 4868 119648 4876 119712
rect 4940 119648 4956 119712
rect 5020 119648 5036 119712
rect 5100 119648 5116 119712
rect 5180 119648 5188 119712
rect 4868 118624 5188 119648
rect 4868 118560 4876 118624
rect 4940 118560 4956 118624
rect 5020 118560 5036 118624
rect 5100 118560 5116 118624
rect 5180 118560 5188 118624
rect 4868 117536 5188 118560
rect 4868 117472 4876 117536
rect 4940 117472 4956 117536
rect 5020 117472 5036 117536
rect 5100 117472 5116 117536
rect 5180 117472 5188 117536
rect 4868 116448 5188 117472
rect 4868 116384 4876 116448
rect 4940 116384 4956 116448
rect 5020 116384 5036 116448
rect 5100 116384 5116 116448
rect 5180 116384 5188 116448
rect 4868 115360 5188 116384
rect 4868 115296 4876 115360
rect 4940 115296 4956 115360
rect 5020 115296 5036 115360
rect 5100 115296 5116 115360
rect 5180 115296 5188 115360
rect 4868 114272 5188 115296
rect 4868 114208 4876 114272
rect 4940 114208 4956 114272
rect 5020 114208 5036 114272
rect 5100 114208 5116 114272
rect 5180 114208 5188 114272
rect 4868 113184 5188 114208
rect 4868 113120 4876 113184
rect 4940 113120 4956 113184
rect 5020 113120 5036 113184
rect 5100 113120 5116 113184
rect 5180 113120 5188 113184
rect 4868 112096 5188 113120
rect 4868 112032 4876 112096
rect 4940 112032 4956 112096
rect 5020 112032 5036 112096
rect 5100 112032 5116 112096
rect 5180 112032 5188 112096
rect 4868 111008 5188 112032
rect 4868 110944 4876 111008
rect 4940 110944 4956 111008
rect 5020 110944 5036 111008
rect 5100 110944 5116 111008
rect 5180 110944 5188 111008
rect 4868 109920 5188 110944
rect 4868 109856 4876 109920
rect 4940 109856 4956 109920
rect 5020 109856 5036 109920
rect 5100 109856 5116 109920
rect 5180 109856 5188 109920
rect 4868 108832 5188 109856
rect 4868 108768 4876 108832
rect 4940 108768 4956 108832
rect 5020 108768 5036 108832
rect 5100 108768 5116 108832
rect 5180 108768 5188 108832
rect 4868 107744 5188 108768
rect 4868 107680 4876 107744
rect 4940 107680 4956 107744
rect 5020 107680 5036 107744
rect 5100 107680 5116 107744
rect 5180 107680 5188 107744
rect 4868 106656 5188 107680
rect 4868 106592 4876 106656
rect 4940 106592 4956 106656
rect 5020 106592 5036 106656
rect 5100 106592 5116 106656
rect 5180 106592 5188 106656
rect 4868 105568 5188 106592
rect 4868 105504 4876 105568
rect 4940 105504 4956 105568
rect 5020 105504 5036 105568
rect 5100 105504 5116 105568
rect 5180 105504 5188 105568
rect 4868 104480 5188 105504
rect 4868 104416 4876 104480
rect 4940 104416 4956 104480
rect 5020 104416 5036 104480
rect 5100 104416 5116 104480
rect 5180 104416 5188 104480
rect 4868 103392 5188 104416
rect 4868 103328 4876 103392
rect 4940 103328 4956 103392
rect 5020 103328 5036 103392
rect 5100 103328 5116 103392
rect 5180 103328 5188 103392
rect 4868 102304 5188 103328
rect 4868 102240 4876 102304
rect 4940 102240 4956 102304
rect 5020 102240 5036 102304
rect 5100 102240 5116 102304
rect 5180 102240 5188 102304
rect 4868 101216 5188 102240
rect 4868 101152 4876 101216
rect 4940 101152 4956 101216
rect 5020 101152 5036 101216
rect 5100 101152 5116 101216
rect 5180 101152 5188 101216
rect 4868 100128 5188 101152
rect 4868 100064 4876 100128
rect 4940 100064 4956 100128
rect 5020 100064 5036 100128
rect 5100 100064 5116 100128
rect 5180 100064 5188 100128
rect 4868 99040 5188 100064
rect 4868 98976 4876 99040
rect 4940 98976 4956 99040
rect 5020 98976 5036 99040
rect 5100 98976 5116 99040
rect 5180 98976 5188 99040
rect 4868 98192 5188 98976
rect 105916 127872 106236 127932
rect 105916 127808 105924 127872
rect 105988 127808 106004 127872
rect 106068 127808 106084 127872
rect 106148 127808 106164 127872
rect 106228 127808 106236 127872
rect 105916 126784 106236 127808
rect 105916 126720 105924 126784
rect 105988 126720 106004 126784
rect 106068 126720 106084 126784
rect 106148 126720 106164 126784
rect 106228 126720 106236 126784
rect 105916 125696 106236 126720
rect 105916 125632 105924 125696
rect 105988 125632 106004 125696
rect 106068 125632 106084 125696
rect 106148 125632 106164 125696
rect 106228 125632 106236 125696
rect 105916 124608 106236 125632
rect 105916 124544 105924 124608
rect 105988 124544 106004 124608
rect 106068 124544 106084 124608
rect 106148 124544 106164 124608
rect 106228 124544 106236 124608
rect 105916 123520 106236 124544
rect 105916 123456 105924 123520
rect 105988 123456 106004 123520
rect 106068 123456 106084 123520
rect 106148 123456 106164 123520
rect 106228 123456 106236 123520
rect 105916 122432 106236 123456
rect 105916 122368 105924 122432
rect 105988 122368 106004 122432
rect 106068 122368 106084 122432
rect 106148 122368 106164 122432
rect 106228 122368 106236 122432
rect 105916 121344 106236 122368
rect 105916 121280 105924 121344
rect 105988 121280 106004 121344
rect 106068 121280 106084 121344
rect 106148 121280 106164 121344
rect 106228 121280 106236 121344
rect 105916 120256 106236 121280
rect 105916 120192 105924 120256
rect 105988 120192 106004 120256
rect 106068 120192 106084 120256
rect 106148 120192 106164 120256
rect 106228 120192 106236 120256
rect 105916 119168 106236 120192
rect 105916 119104 105924 119168
rect 105988 119104 106004 119168
rect 106068 119104 106084 119168
rect 106148 119104 106164 119168
rect 106228 119104 106236 119168
rect 105916 118080 106236 119104
rect 105916 118016 105924 118080
rect 105988 118016 106004 118080
rect 106068 118016 106084 118080
rect 106148 118016 106164 118080
rect 106228 118016 106236 118080
rect 105916 116992 106236 118016
rect 105916 116928 105924 116992
rect 105988 116928 106004 116992
rect 106068 116928 106084 116992
rect 106148 116928 106164 116992
rect 106228 116928 106236 116992
rect 105916 115904 106236 116928
rect 105916 115840 105924 115904
rect 105988 115840 106004 115904
rect 106068 115840 106084 115904
rect 106148 115840 106164 115904
rect 106228 115840 106236 115904
rect 105916 114816 106236 115840
rect 105916 114752 105924 114816
rect 105988 114752 106004 114816
rect 106068 114752 106084 114816
rect 106148 114752 106164 114816
rect 106228 114752 106236 114816
rect 105916 113728 106236 114752
rect 105916 113664 105924 113728
rect 105988 113664 106004 113728
rect 106068 113664 106084 113728
rect 106148 113664 106164 113728
rect 106228 113664 106236 113728
rect 105916 112640 106236 113664
rect 105916 112576 105924 112640
rect 105988 112576 106004 112640
rect 106068 112576 106084 112640
rect 106148 112576 106164 112640
rect 106228 112576 106236 112640
rect 105916 111552 106236 112576
rect 105916 111488 105924 111552
rect 105988 111488 106004 111552
rect 106068 111488 106084 111552
rect 106148 111488 106164 111552
rect 106228 111488 106236 111552
rect 105916 110464 106236 111488
rect 105916 110400 105924 110464
rect 105988 110400 106004 110464
rect 106068 110400 106084 110464
rect 106148 110400 106164 110464
rect 106228 110400 106236 110464
rect 105916 109376 106236 110400
rect 105916 109312 105924 109376
rect 105988 109312 106004 109376
rect 106068 109312 106084 109376
rect 106148 109312 106164 109376
rect 106228 109312 106236 109376
rect 105916 108288 106236 109312
rect 105916 108224 105924 108288
rect 105988 108224 106004 108288
rect 106068 108224 106084 108288
rect 106148 108224 106164 108288
rect 106228 108224 106236 108288
rect 105916 107200 106236 108224
rect 105916 107136 105924 107200
rect 105988 107136 106004 107200
rect 106068 107136 106084 107200
rect 106148 107136 106164 107200
rect 106228 107136 106236 107200
rect 105916 106112 106236 107136
rect 105916 106048 105924 106112
rect 105988 106048 106004 106112
rect 106068 106048 106084 106112
rect 106148 106048 106164 106112
rect 106228 106048 106236 106112
rect 105916 105024 106236 106048
rect 105916 104960 105924 105024
rect 105988 104960 106004 105024
rect 106068 104960 106084 105024
rect 106148 104960 106164 105024
rect 106228 104960 106236 105024
rect 105916 103936 106236 104960
rect 105916 103872 105924 103936
rect 105988 103872 106004 103936
rect 106068 103872 106084 103936
rect 106148 103872 106164 103936
rect 106228 103872 106236 103936
rect 105916 102848 106236 103872
rect 105916 102784 105924 102848
rect 105988 102784 106004 102848
rect 106068 102784 106084 102848
rect 106148 102784 106164 102848
rect 106228 102784 106236 102848
rect 105916 101760 106236 102784
rect 105916 101696 105924 101760
rect 105988 101696 106004 101760
rect 106068 101696 106084 101760
rect 106148 101696 106164 101760
rect 106228 101696 106236 101760
rect 105916 100672 106236 101696
rect 105916 100608 105924 100672
rect 105988 100608 106004 100672
rect 106068 100608 106084 100672
rect 106148 100608 106164 100672
rect 106228 100608 106236 100672
rect 105916 99584 106236 100608
rect 105916 99520 105924 99584
rect 105988 99520 106004 99584
rect 106068 99520 106084 99584
rect 106148 99520 106164 99584
rect 106228 99520 106236 99584
rect 105916 98496 106236 99520
rect 105916 98432 105924 98496
rect 105988 98432 106004 98496
rect 106068 98432 106084 98496
rect 106148 98432 106164 98496
rect 106228 98432 106236 98496
rect 4868 97956 4910 98192
rect 5146 97956 5188 98192
rect 4868 97952 5188 97956
rect 4868 97888 4876 97952
rect 4940 97888 4956 97952
rect 5020 97888 5036 97952
rect 5100 97888 5116 97952
rect 5180 97888 5188 97952
rect 10696 98192 11044 98234
rect 10696 97956 10752 98192
rect 10988 97956 11044 98192
rect 10696 97914 11044 97956
rect 100936 98192 101284 98234
rect 100936 97956 100992 98192
rect 101228 97956 101284 98192
rect 100936 97914 101284 97956
rect 4868 96864 5188 97888
rect 10000 97532 10348 97574
rect 10000 97296 10056 97532
rect 10292 97296 10348 97532
rect 10000 97254 10348 97296
rect 101632 97532 101980 97574
rect 101632 97296 101688 97532
rect 101924 97296 101980 97532
rect 101632 97254 101980 97296
rect 105916 97532 106236 98432
rect 105916 97408 105958 97532
rect 106194 97408 106236 97532
rect 105916 97344 105924 97408
rect 106228 97344 106236 97408
rect 105916 97296 105958 97344
rect 106194 97296 106236 97344
rect 4868 96800 4876 96864
rect 4940 96800 4956 96864
rect 5020 96800 5036 96864
rect 5100 96800 5116 96864
rect 5180 96800 5188 96864
rect 4868 95776 5188 96800
rect 4868 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5188 95776
rect 4868 94688 5188 95712
rect 4868 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5188 94688
rect 4868 93600 5188 94624
rect 4868 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5188 93600
rect 4868 92512 5188 93536
rect 4868 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5188 92512
rect 4868 91424 5188 92448
rect 4868 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5188 91424
rect 4868 90336 5188 91360
rect 4868 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5188 90336
rect 4868 89248 5188 90272
rect 4868 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5188 89248
rect 4868 88160 5188 89184
rect 4868 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5188 88160
rect 4868 87072 5188 88096
rect 4868 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5188 87072
rect 4868 85984 5188 87008
rect 4868 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5188 85984
rect 4868 84896 5188 85920
rect 4868 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5188 84896
rect 4868 83808 5188 84832
rect 4868 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5188 83808
rect 4868 82720 5188 83744
rect 4868 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5188 82720
rect 4868 81632 5188 82656
rect 4868 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5188 81632
rect 4868 80544 5188 81568
rect 4868 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5188 80544
rect 4868 79456 5188 80480
rect 105916 96320 106236 97296
rect 105916 96256 105924 96320
rect 105988 96256 106004 96320
rect 106068 96256 106084 96320
rect 106148 96256 106164 96320
rect 106228 96256 106236 96320
rect 105916 95232 106236 96256
rect 105916 95168 105924 95232
rect 105988 95168 106004 95232
rect 106068 95168 106084 95232
rect 106148 95168 106164 95232
rect 106228 95168 106236 95232
rect 105916 94144 106236 95168
rect 105916 94080 105924 94144
rect 105988 94080 106004 94144
rect 106068 94080 106084 94144
rect 106148 94080 106164 94144
rect 106228 94080 106236 94144
rect 105916 93056 106236 94080
rect 105916 92992 105924 93056
rect 105988 92992 106004 93056
rect 106068 92992 106084 93056
rect 106148 92992 106164 93056
rect 106228 92992 106236 93056
rect 105916 91968 106236 92992
rect 105916 91904 105924 91968
rect 105988 91904 106004 91968
rect 106068 91904 106084 91968
rect 106148 91904 106164 91968
rect 106228 91904 106236 91968
rect 105916 90880 106236 91904
rect 105916 90816 105924 90880
rect 105988 90816 106004 90880
rect 106068 90816 106084 90880
rect 106148 90816 106164 90880
rect 106228 90816 106236 90880
rect 105916 89792 106236 90816
rect 105916 89728 105924 89792
rect 105988 89728 106004 89792
rect 106068 89728 106084 89792
rect 106148 89728 106164 89792
rect 106228 89728 106236 89792
rect 105916 88704 106236 89728
rect 105916 88640 105924 88704
rect 105988 88640 106004 88704
rect 106068 88640 106084 88704
rect 106148 88640 106164 88704
rect 106228 88640 106236 88704
rect 105916 87616 106236 88640
rect 105916 87552 105924 87616
rect 105988 87552 106004 87616
rect 106068 87552 106084 87616
rect 106148 87552 106164 87616
rect 106228 87552 106236 87616
rect 105916 86528 106236 87552
rect 105916 86464 105924 86528
rect 105988 86464 106004 86528
rect 106068 86464 106084 86528
rect 106148 86464 106164 86528
rect 106228 86464 106236 86528
rect 105916 85440 106236 86464
rect 105916 85376 105924 85440
rect 105988 85376 106004 85440
rect 106068 85376 106084 85440
rect 106148 85376 106164 85440
rect 106228 85376 106236 85440
rect 105916 84352 106236 85376
rect 105916 84288 105924 84352
rect 105988 84288 106004 84352
rect 106068 84288 106084 84352
rect 106148 84288 106164 84352
rect 106228 84288 106236 84352
rect 105916 83264 106236 84288
rect 105916 83200 105924 83264
rect 105988 83200 106004 83264
rect 106068 83200 106084 83264
rect 106148 83200 106164 83264
rect 106228 83200 106236 83264
rect 105916 82176 106236 83200
rect 105916 82112 105924 82176
rect 105988 82112 106004 82176
rect 106068 82112 106084 82176
rect 106148 82112 106164 82176
rect 106228 82112 106236 82176
rect 105916 81088 106236 82112
rect 105916 81024 105924 81088
rect 105988 81024 106004 81088
rect 106068 81024 106084 81088
rect 106148 81024 106164 81088
rect 106228 81024 106236 81088
rect 4868 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5188 79456
rect 4868 78368 5188 79392
rect 4868 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5188 78368
rect 4868 77280 5188 78304
rect 16070 78029 16130 80038
rect 23430 79253 23490 80038
rect 24608 79525 24668 80038
rect 25776 79661 25836 80038
rect 25773 79660 25839 79661
rect 25773 79596 25774 79660
rect 25838 79596 25839 79660
rect 25773 79595 25839 79596
rect 24605 79524 24671 79525
rect 24605 79460 24606 79524
rect 24670 79460 24671 79524
rect 24605 79459 24671 79460
rect 26926 79389 26986 80038
rect 28122 79658 28182 80038
rect 28122 79598 28274 79658
rect 26923 79388 26989 79389
rect 26923 79324 26924 79388
rect 26988 79324 26989 79388
rect 26923 79323 26989 79324
rect 23427 79252 23493 79253
rect 23427 79188 23428 79252
rect 23492 79188 23493 79252
rect 23427 79187 23493 79188
rect 23430 78845 23490 79187
rect 23427 78844 23493 78845
rect 23427 78780 23428 78844
rect 23492 78780 23493 78844
rect 23427 78779 23493 78780
rect 16067 78028 16133 78029
rect 16067 77964 16068 78028
rect 16132 77964 16133 78028
rect 16067 77963 16133 77964
rect 28214 77757 28274 79598
rect 29280 79525 29340 80038
rect 30448 79797 30508 80038
rect 31616 79933 31676 80038
rect 31613 79932 31679 79933
rect 31613 79868 31614 79932
rect 31678 79868 31679 79932
rect 31613 79867 31679 79868
rect 30445 79796 30511 79797
rect 30445 79732 30446 79796
rect 30510 79732 30511 79796
rect 30445 79731 30511 79732
rect 30448 79525 30508 79731
rect 31616 79525 31676 79867
rect 32784 79797 32844 80038
rect 32781 79796 32847 79797
rect 32781 79732 32782 79796
rect 32846 79732 32847 79796
rect 32781 79731 32847 79732
rect 33952 79525 34012 80038
rect 35114 79525 35174 80038
rect 36288 79933 36348 80038
rect 36285 79932 36351 79933
rect 36285 79868 36286 79932
rect 36350 79868 36351 79932
rect 36285 79867 36351 79868
rect 37456 79661 37516 80038
rect 38624 79933 38684 80038
rect 39792 79933 39852 80038
rect 40960 79933 41020 80038
rect 38621 79932 38687 79933
rect 38621 79868 38622 79932
rect 38686 79868 38687 79932
rect 38621 79867 38687 79868
rect 39789 79932 39855 79933
rect 39789 79868 39790 79932
rect 39854 79868 39855 79932
rect 39789 79867 39855 79868
rect 40957 79932 41023 79933
rect 40957 79868 40958 79932
rect 41022 79868 41023 79932
rect 40957 79867 41023 79868
rect 37453 79660 37519 79661
rect 37453 79596 37454 79660
rect 37518 79596 37519 79660
rect 37453 79595 37519 79596
rect 42128 79525 42188 80038
rect 43296 79525 43356 80038
rect 90529 79930 90589 80038
rect 90406 79870 90589 79930
rect 29277 79524 29343 79525
rect 29277 79460 29278 79524
rect 29342 79460 29343 79524
rect 29277 79459 29343 79460
rect 30445 79524 30511 79525
rect 30445 79460 30446 79524
rect 30510 79460 30511 79524
rect 30445 79459 30511 79460
rect 31613 79524 31679 79525
rect 31613 79460 31614 79524
rect 31678 79460 31679 79524
rect 31613 79459 31679 79460
rect 33949 79524 34015 79525
rect 33949 79460 33950 79524
rect 34014 79460 34015 79524
rect 33949 79459 34015 79460
rect 35111 79524 35177 79525
rect 35111 79460 35112 79524
rect 35176 79460 35177 79524
rect 35111 79459 35177 79460
rect 42125 79524 42191 79525
rect 42125 79460 42126 79524
rect 42190 79460 42191 79524
rect 42125 79459 42191 79460
rect 43293 79524 43359 79525
rect 43293 79460 43294 79524
rect 43358 79460 43359 79524
rect 43293 79459 43359 79460
rect 34928 77824 35248 77880
rect 34928 77760 34936 77824
rect 35000 77760 35016 77824
rect 35080 77760 35096 77824
rect 35160 77760 35176 77824
rect 35240 77760 35248 77824
rect 28211 77756 28277 77757
rect 28211 77692 28212 77756
rect 28276 77692 28277 77756
rect 28211 77691 28277 77692
rect 4868 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5188 77280
rect 4868 76192 5188 77216
rect 4868 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5188 76192
rect 4868 75104 5188 76128
rect 4868 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5188 75104
rect 4868 74016 5188 75040
rect 4868 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5188 74016
rect 4868 72928 5188 73952
rect 4868 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5188 72928
rect 4868 71840 5188 72864
rect 4868 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5188 71840
rect 4868 70752 5188 71776
rect 4868 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5188 70752
rect 4868 69664 5188 70688
rect 4868 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5188 69664
rect 4868 68576 5188 69600
rect 4868 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5188 68576
rect 4868 67556 5188 68512
rect 4868 67488 4910 67556
rect 5146 67488 5188 67556
rect 4868 67424 4876 67488
rect 5180 67424 5188 67488
rect 4868 67320 4910 67424
rect 5146 67320 5188 67424
rect 4868 66400 5188 67320
rect 4868 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5188 66400
rect 4868 65312 5188 66336
rect 34928 76736 35248 77760
rect 34928 76672 34936 76736
rect 35000 76672 35016 76736
rect 35080 76672 35096 76736
rect 35160 76672 35176 76736
rect 35240 76672 35248 76736
rect 34928 75648 35248 76672
rect 34928 75584 34936 75648
rect 35000 75584 35016 75648
rect 35080 75584 35096 75648
rect 35160 75584 35176 75648
rect 35240 75584 35248 75648
rect 34928 74560 35248 75584
rect 34928 74496 34936 74560
rect 35000 74496 35016 74560
rect 35080 74496 35096 74560
rect 35160 74496 35176 74560
rect 35240 74496 35248 74560
rect 34928 73472 35248 74496
rect 34928 73408 34936 73472
rect 35000 73408 35016 73472
rect 35080 73408 35096 73472
rect 35160 73408 35176 73472
rect 35240 73408 35248 73472
rect 34928 72384 35248 73408
rect 34928 72320 34936 72384
rect 35000 72320 35016 72384
rect 35080 72320 35096 72384
rect 35160 72320 35176 72384
rect 35240 72320 35248 72384
rect 34928 71296 35248 72320
rect 34928 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35248 71296
rect 34928 70208 35248 71232
rect 34928 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35248 70208
rect 34928 69120 35248 70144
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 68032 35248 69056
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 66944 35248 67968
rect 34928 66880 34936 66944
rect 35000 66896 35016 66944
rect 35080 66896 35096 66944
rect 35160 66896 35176 66944
rect 35240 66880 35248 66944
rect 34928 66660 34970 66880
rect 35206 66660 35248 66880
rect 34928 65856 35248 66660
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 65650 35248 65792
rect 35588 77280 35908 78064
rect 35588 77216 35596 77280
rect 35660 77216 35676 77280
rect 35740 77216 35756 77280
rect 35820 77216 35836 77280
rect 35900 77216 35908 77280
rect 35588 76192 35908 77216
rect 35588 76128 35596 76192
rect 35660 76128 35676 76192
rect 35740 76128 35756 76192
rect 35820 76128 35836 76192
rect 35900 76128 35908 76192
rect 35588 75104 35908 76128
rect 35588 75040 35596 75104
rect 35660 75040 35676 75104
rect 35740 75040 35756 75104
rect 35820 75040 35836 75104
rect 35900 75040 35908 75104
rect 35588 74016 35908 75040
rect 35588 73952 35596 74016
rect 35660 73952 35676 74016
rect 35740 73952 35756 74016
rect 35820 73952 35836 74016
rect 35900 73952 35908 74016
rect 35588 72928 35908 73952
rect 35588 72864 35596 72928
rect 35660 72864 35676 72928
rect 35740 72864 35756 72928
rect 35820 72864 35836 72928
rect 35900 72864 35908 72928
rect 35588 71840 35908 72864
rect 35588 71776 35596 71840
rect 35660 71776 35676 71840
rect 35740 71776 35756 71840
rect 35820 71776 35836 71840
rect 35900 71776 35908 71840
rect 35588 70752 35908 71776
rect 35588 70688 35596 70752
rect 35660 70688 35676 70752
rect 35740 70688 35756 70752
rect 35820 70688 35836 70752
rect 35900 70688 35908 70752
rect 35588 69664 35908 70688
rect 35588 69600 35596 69664
rect 35660 69600 35676 69664
rect 35740 69600 35756 69664
rect 35820 69600 35836 69664
rect 35900 69600 35908 69664
rect 35588 68576 35908 69600
rect 35588 68512 35596 68576
rect 35660 68512 35676 68576
rect 35740 68512 35756 68576
rect 35820 68512 35836 68576
rect 35900 68512 35908 68576
rect 35588 67556 35908 68512
rect 35588 67488 35630 67556
rect 35866 67488 35908 67556
rect 35588 67424 35596 67488
rect 35900 67424 35908 67488
rect 35588 67320 35630 67424
rect 35866 67320 35908 67424
rect 35588 66400 35908 67320
rect 35588 66336 35596 66400
rect 35660 66336 35676 66400
rect 35740 66336 35756 66400
rect 35820 66336 35836 66400
rect 35900 66336 35908 66400
rect 35588 65650 35908 66336
rect 65648 77824 65968 78064
rect 65648 77760 65656 77824
rect 65720 77760 65736 77824
rect 65800 77760 65816 77824
rect 65880 77760 65896 77824
rect 65960 77760 65968 77824
rect 65648 76736 65968 77760
rect 65648 76672 65656 76736
rect 65720 76672 65736 76736
rect 65800 76672 65816 76736
rect 65880 76672 65896 76736
rect 65960 76672 65968 76736
rect 65648 75648 65968 76672
rect 65648 75584 65656 75648
rect 65720 75584 65736 75648
rect 65800 75584 65816 75648
rect 65880 75584 65896 75648
rect 65960 75584 65968 75648
rect 65648 74560 65968 75584
rect 65648 74496 65656 74560
rect 65720 74496 65736 74560
rect 65800 74496 65816 74560
rect 65880 74496 65896 74560
rect 65960 74496 65968 74560
rect 65648 73472 65968 74496
rect 65648 73408 65656 73472
rect 65720 73408 65736 73472
rect 65800 73408 65816 73472
rect 65880 73408 65896 73472
rect 65960 73408 65968 73472
rect 65648 72384 65968 73408
rect 65648 72320 65656 72384
rect 65720 72320 65736 72384
rect 65800 72320 65816 72384
rect 65880 72320 65896 72384
rect 65960 72320 65968 72384
rect 65648 71296 65968 72320
rect 65648 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65968 71296
rect 65648 70208 65968 71232
rect 65648 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65968 70208
rect 65648 69120 65968 70144
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 68032 65968 69056
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 66944 65968 67968
rect 65648 66880 65656 66944
rect 65720 66896 65736 66944
rect 65800 66896 65816 66944
rect 65880 66896 65896 66944
rect 65960 66880 65968 66944
rect 65648 66660 65690 66880
rect 65926 66660 65968 66880
rect 36123 66196 36189 66197
rect 36123 66132 36124 66196
rect 36188 66132 36189 66196
rect 36123 66131 36189 66132
rect 38515 66196 38581 66197
rect 38515 66132 38516 66196
rect 38580 66132 38581 66196
rect 38515 66131 38581 66132
rect 41091 66196 41157 66197
rect 41091 66132 41092 66196
rect 41156 66132 41157 66196
rect 41091 66131 41157 66132
rect 43667 66196 43733 66197
rect 43667 66132 43668 66196
rect 43732 66132 43733 66196
rect 43667 66131 43733 66132
rect 46059 66196 46125 66197
rect 46059 66132 46060 66196
rect 46124 66132 46125 66196
rect 46059 66131 46125 66132
rect 48635 66196 48701 66197
rect 48635 66132 48636 66196
rect 48700 66132 48701 66196
rect 48635 66131 48701 66132
rect 51027 66196 51093 66197
rect 51027 66132 51028 66196
rect 51092 66132 51093 66196
rect 51027 66131 51093 66132
rect 53603 66196 53669 66197
rect 53603 66132 53604 66196
rect 53668 66132 53669 66196
rect 53603 66131 53669 66132
rect 55995 66196 56061 66197
rect 55995 66132 55996 66196
rect 56060 66132 56061 66196
rect 55995 66131 56061 66132
rect 58571 66196 58637 66197
rect 58571 66132 58572 66196
rect 58636 66132 58637 66196
rect 58571 66131 58637 66132
rect 61147 66196 61213 66197
rect 61147 66132 61148 66196
rect 61212 66132 61213 66196
rect 61147 66131 61213 66132
rect 63539 66196 63605 66197
rect 63539 66132 63540 66196
rect 63604 66132 63605 66196
rect 63539 66131 63605 66132
rect 4868 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5188 65312
rect 4868 64224 5188 65248
rect 36126 64290 36186 66131
rect 4868 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5188 64224
rect 4868 63136 5188 64160
rect 36077 64230 36186 64290
rect 38518 64290 38578 66131
rect 41094 64290 41154 66131
rect 43670 64290 43730 66131
rect 38518 64230 38633 64290
rect 36077 63676 36137 64230
rect 38573 63676 38633 64230
rect 41069 64230 41154 64290
rect 43578 64230 43730 64290
rect 41069 63676 41129 64230
rect 43578 63676 43638 64230
rect 46062 63676 46122 66131
rect 48638 64290 48698 66131
rect 48557 64230 48698 64290
rect 51030 64290 51090 66131
rect 53606 64290 53666 66131
rect 51030 64230 51113 64290
rect 48557 63676 48617 64230
rect 51053 63676 51113 64230
rect 53549 64230 53666 64290
rect 55998 64290 56058 66131
rect 58574 64290 58634 66131
rect 61150 64290 61210 66131
rect 55998 64230 56105 64290
rect 53549 63676 53609 64230
rect 56045 63676 56105 64230
rect 58541 64230 58634 64290
rect 61058 64230 61210 64290
rect 58541 63676 58601 64230
rect 61058 63676 61118 64230
rect 63542 63676 63602 66131
rect 65648 65856 65968 66660
rect 66308 77280 66628 78064
rect 66308 77216 66316 77280
rect 66380 77216 66396 77280
rect 66460 77216 66476 77280
rect 66540 77216 66556 77280
rect 66620 77216 66628 77280
rect 66308 76192 66628 77216
rect 90406 77213 90466 79870
rect 90682 79525 90742 80038
rect 90816 79933 90876 80038
rect 105916 80000 106236 81024
rect 105916 79936 105924 80000
rect 105988 79936 106004 80000
rect 106068 79936 106084 80000
rect 106148 79936 106164 80000
rect 106228 79936 106236 80000
rect 90813 79932 90879 79933
rect 90813 79868 90814 79932
rect 90878 79868 90879 79932
rect 90813 79867 90879 79868
rect 90679 79524 90745 79525
rect 90679 79460 90680 79524
rect 90744 79460 90745 79524
rect 90679 79459 90745 79460
rect 105916 78912 106236 79936
rect 105916 78848 105924 78912
rect 105988 78848 106004 78912
rect 106068 78848 106084 78912
rect 106148 78848 106164 78912
rect 106228 78848 106236 78912
rect 96368 77824 96688 78064
rect 96368 77760 96376 77824
rect 96440 77760 96456 77824
rect 96520 77760 96536 77824
rect 96600 77760 96616 77824
rect 96680 77760 96688 77824
rect 90403 77212 90469 77213
rect 90403 77148 90404 77212
rect 90468 77148 90469 77212
rect 90403 77147 90469 77148
rect 66308 76128 66316 76192
rect 66380 76128 66396 76192
rect 66460 76128 66476 76192
rect 66540 76128 66556 76192
rect 66620 76128 66628 76192
rect 66308 75104 66628 76128
rect 66308 75040 66316 75104
rect 66380 75040 66396 75104
rect 66460 75040 66476 75104
rect 66540 75040 66556 75104
rect 66620 75040 66628 75104
rect 66308 74016 66628 75040
rect 66308 73952 66316 74016
rect 66380 73952 66396 74016
rect 66460 73952 66476 74016
rect 66540 73952 66556 74016
rect 66620 73952 66628 74016
rect 66308 72928 66628 73952
rect 66308 72864 66316 72928
rect 66380 72864 66396 72928
rect 66460 72864 66476 72928
rect 66540 72864 66556 72928
rect 66620 72864 66628 72928
rect 66308 71840 66628 72864
rect 66308 71776 66316 71840
rect 66380 71776 66396 71840
rect 66460 71776 66476 71840
rect 66540 71776 66556 71840
rect 66620 71776 66628 71840
rect 66308 70752 66628 71776
rect 66308 70688 66316 70752
rect 66380 70688 66396 70752
rect 66460 70688 66476 70752
rect 66540 70688 66556 70752
rect 66620 70688 66628 70752
rect 66308 69664 66628 70688
rect 66308 69600 66316 69664
rect 66380 69600 66396 69664
rect 66460 69600 66476 69664
rect 66540 69600 66556 69664
rect 66620 69600 66628 69664
rect 66308 68576 66628 69600
rect 96368 76736 96688 77760
rect 96368 76672 96376 76736
rect 96440 76672 96456 76736
rect 96520 76672 96536 76736
rect 96600 76672 96616 76736
rect 96680 76672 96688 76736
rect 96368 75648 96688 76672
rect 96368 75584 96376 75648
rect 96440 75584 96456 75648
rect 96520 75584 96536 75648
rect 96600 75584 96616 75648
rect 96680 75584 96688 75648
rect 96368 74560 96688 75584
rect 96368 74496 96376 74560
rect 96440 74496 96456 74560
rect 96520 74496 96536 74560
rect 96600 74496 96616 74560
rect 96680 74496 96688 74560
rect 96368 73472 96688 74496
rect 96368 73408 96376 73472
rect 96440 73408 96456 73472
rect 96520 73408 96536 73472
rect 96600 73408 96616 73472
rect 96680 73408 96688 73472
rect 96368 72384 96688 73408
rect 96368 72320 96376 72384
rect 96440 72320 96456 72384
rect 96520 72320 96536 72384
rect 96600 72320 96616 72384
rect 96680 72320 96688 72384
rect 96368 71296 96688 72320
rect 96368 71232 96376 71296
rect 96440 71232 96456 71296
rect 96520 71232 96536 71296
rect 96600 71232 96616 71296
rect 96680 71232 96688 71296
rect 96368 70208 96688 71232
rect 96368 70144 96376 70208
rect 96440 70144 96456 70208
rect 96520 70144 96536 70208
rect 96600 70144 96616 70208
rect 96680 70144 96688 70208
rect 96368 69120 96688 70144
rect 96368 69056 96376 69120
rect 96440 69056 96456 69120
rect 96520 69056 96536 69120
rect 96600 69056 96616 69120
rect 96680 69056 96688 69120
rect 87275 69052 87341 69053
rect 87275 68988 87276 69052
rect 87340 68988 87341 69052
rect 87275 68987 87341 68988
rect 66308 68512 66316 68576
rect 66380 68512 66396 68576
rect 66460 68512 66476 68576
rect 66540 68512 66556 68576
rect 66620 68512 66628 68576
rect 66308 67556 66628 68512
rect 66308 67488 66350 67556
rect 66586 67488 66628 67556
rect 66308 67424 66316 67488
rect 66620 67424 66628 67488
rect 66308 67320 66350 67424
rect 66586 67320 66628 67424
rect 66308 66400 66628 67320
rect 66308 66336 66316 66400
rect 66380 66336 66396 66400
rect 66460 66336 66476 66400
rect 66540 66336 66556 66400
rect 66620 66336 66628 66400
rect 66115 66196 66181 66197
rect 66115 66132 66116 66196
rect 66180 66132 66181 66196
rect 66115 66131 66181 66132
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 65776 65968 65792
rect 66118 64290 66178 66131
rect 66308 65650 66628 66336
rect 68507 66196 68573 66197
rect 68507 66132 68508 66196
rect 68572 66132 68573 66196
rect 68507 66131 68573 66132
rect 71083 66196 71149 66197
rect 71083 66132 71084 66196
rect 71148 66132 71149 66196
rect 71083 66131 71149 66132
rect 73475 66196 73541 66197
rect 73475 66132 73476 66196
rect 73540 66132 73541 66196
rect 73475 66131 73541 66132
rect 86171 66196 86237 66197
rect 86171 66132 86172 66196
rect 86236 66132 86237 66196
rect 86171 66131 86237 66132
rect 66029 64230 66178 64290
rect 66029 63676 66089 64230
rect 68510 63676 68570 66131
rect 71086 64290 71146 66131
rect 71021 64230 71146 64290
rect 73478 64290 73538 66131
rect 86174 64290 86234 66131
rect 73478 64230 73577 64290
rect 71021 63676 71081 64230
rect 73517 63676 73577 64230
rect 86144 64230 86234 64290
rect 87278 64290 87338 68987
rect 96368 68032 96688 69056
rect 96368 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96688 68032
rect 96368 66944 96688 67968
rect 96368 66880 96376 66944
rect 96440 66896 96456 66944
rect 96520 66896 96536 66944
rect 96600 66896 96616 66944
rect 96680 66880 96688 66944
rect 96368 66660 96410 66880
rect 96646 66660 96688 66880
rect 96368 65856 96688 66660
rect 96368 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96688 65856
rect 96368 65650 96688 65792
rect 97028 77280 97348 78064
rect 97028 77216 97036 77280
rect 97100 77216 97116 77280
rect 97180 77216 97196 77280
rect 97260 77216 97276 77280
rect 97340 77216 97348 77280
rect 97028 76192 97348 77216
rect 105916 77824 106236 78848
rect 105916 77760 105924 77824
rect 105988 77760 106004 77824
rect 106068 77760 106084 77824
rect 106148 77760 106164 77824
rect 106228 77760 106236 77824
rect 105916 77200 106236 77760
rect 106652 136032 106972 136592
rect 106652 135968 106660 136032
rect 106724 135968 106740 136032
rect 106804 135968 106820 136032
rect 106884 135968 106900 136032
rect 106964 135968 106972 136032
rect 106652 134944 106972 135968
rect 106652 134880 106660 134944
rect 106724 134880 106740 134944
rect 106804 134880 106820 134944
rect 106884 134880 106900 134944
rect 106964 134880 106972 134944
rect 106652 133856 106972 134880
rect 106652 133792 106660 133856
rect 106724 133792 106740 133856
rect 106804 133792 106820 133856
rect 106884 133792 106900 133856
rect 106964 133792 106972 133856
rect 106652 132768 106972 133792
rect 106652 132704 106660 132768
rect 106724 132704 106740 132768
rect 106804 132704 106820 132768
rect 106884 132704 106900 132768
rect 106964 132704 106972 132768
rect 106652 131680 106972 132704
rect 106652 131616 106660 131680
rect 106724 131616 106740 131680
rect 106804 131616 106820 131680
rect 106884 131616 106900 131680
rect 106964 131616 106972 131680
rect 106652 130592 106972 131616
rect 106652 130528 106660 130592
rect 106724 130528 106740 130592
rect 106804 130528 106820 130592
rect 106884 130528 106900 130592
rect 106964 130528 106972 130592
rect 106652 129504 106972 130528
rect 106652 129440 106660 129504
rect 106724 129440 106740 129504
rect 106804 129440 106820 129504
rect 106884 129440 106900 129504
rect 106964 129440 106972 129504
rect 106652 128828 106972 129440
rect 106652 128592 106694 128828
rect 106930 128592 106972 128828
rect 106652 128416 106972 128592
rect 106652 128352 106660 128416
rect 106724 128352 106740 128416
rect 106804 128352 106820 128416
rect 106884 128352 106900 128416
rect 106964 128352 106972 128416
rect 106652 127328 106972 128352
rect 106652 127264 106660 127328
rect 106724 127264 106740 127328
rect 106804 127264 106820 127328
rect 106884 127264 106900 127328
rect 106964 127264 106972 127328
rect 106652 126240 106972 127264
rect 106652 126176 106660 126240
rect 106724 126176 106740 126240
rect 106804 126176 106820 126240
rect 106884 126176 106900 126240
rect 106964 126176 106972 126240
rect 106652 125152 106972 126176
rect 106652 125088 106660 125152
rect 106724 125088 106740 125152
rect 106804 125088 106820 125152
rect 106884 125088 106900 125152
rect 106964 125088 106972 125152
rect 106652 124064 106972 125088
rect 106652 124000 106660 124064
rect 106724 124000 106740 124064
rect 106804 124000 106820 124064
rect 106884 124000 106900 124064
rect 106964 124000 106972 124064
rect 106652 122976 106972 124000
rect 106652 122912 106660 122976
rect 106724 122912 106740 122976
rect 106804 122912 106820 122976
rect 106884 122912 106900 122976
rect 106964 122912 106972 122976
rect 106652 121888 106972 122912
rect 106652 121824 106660 121888
rect 106724 121824 106740 121888
rect 106804 121824 106820 121888
rect 106884 121824 106900 121888
rect 106964 121824 106972 121888
rect 106652 120800 106972 121824
rect 106652 120736 106660 120800
rect 106724 120736 106740 120800
rect 106804 120736 106820 120800
rect 106884 120736 106900 120800
rect 106964 120736 106972 120800
rect 106652 119712 106972 120736
rect 106652 119648 106660 119712
rect 106724 119648 106740 119712
rect 106804 119648 106820 119712
rect 106884 119648 106900 119712
rect 106964 119648 106972 119712
rect 106652 118624 106972 119648
rect 106652 118560 106660 118624
rect 106724 118560 106740 118624
rect 106804 118560 106820 118624
rect 106884 118560 106900 118624
rect 106964 118560 106972 118624
rect 106652 117536 106972 118560
rect 106652 117472 106660 117536
rect 106724 117472 106740 117536
rect 106804 117472 106820 117536
rect 106884 117472 106900 117536
rect 106964 117472 106972 117536
rect 106652 116448 106972 117472
rect 106652 116384 106660 116448
rect 106724 116384 106740 116448
rect 106804 116384 106820 116448
rect 106884 116384 106900 116448
rect 106964 116384 106972 116448
rect 106652 115360 106972 116384
rect 106652 115296 106660 115360
rect 106724 115296 106740 115360
rect 106804 115296 106820 115360
rect 106884 115296 106900 115360
rect 106964 115296 106972 115360
rect 106652 114272 106972 115296
rect 106652 114208 106660 114272
rect 106724 114208 106740 114272
rect 106804 114208 106820 114272
rect 106884 114208 106900 114272
rect 106964 114208 106972 114272
rect 106652 113184 106972 114208
rect 106652 113120 106660 113184
rect 106724 113120 106740 113184
rect 106804 113120 106820 113184
rect 106884 113120 106900 113184
rect 106964 113120 106972 113184
rect 106652 112096 106972 113120
rect 106652 112032 106660 112096
rect 106724 112032 106740 112096
rect 106804 112032 106820 112096
rect 106884 112032 106900 112096
rect 106964 112032 106972 112096
rect 106652 111008 106972 112032
rect 106652 110944 106660 111008
rect 106724 110944 106740 111008
rect 106804 110944 106820 111008
rect 106884 110944 106900 111008
rect 106964 110944 106972 111008
rect 106652 109920 106972 110944
rect 106652 109856 106660 109920
rect 106724 109856 106740 109920
rect 106804 109856 106820 109920
rect 106884 109856 106900 109920
rect 106964 109856 106972 109920
rect 106652 108832 106972 109856
rect 106652 108768 106660 108832
rect 106724 108768 106740 108832
rect 106804 108768 106820 108832
rect 106884 108768 106900 108832
rect 106964 108768 106972 108832
rect 106652 107744 106972 108768
rect 106652 107680 106660 107744
rect 106724 107680 106740 107744
rect 106804 107680 106820 107744
rect 106884 107680 106900 107744
rect 106964 107680 106972 107744
rect 106652 106656 106972 107680
rect 106652 106592 106660 106656
rect 106724 106592 106740 106656
rect 106804 106592 106820 106656
rect 106884 106592 106900 106656
rect 106964 106592 106972 106656
rect 106652 105568 106972 106592
rect 106652 105504 106660 105568
rect 106724 105504 106740 105568
rect 106804 105504 106820 105568
rect 106884 105504 106900 105568
rect 106964 105504 106972 105568
rect 106652 104480 106972 105504
rect 106652 104416 106660 104480
rect 106724 104416 106740 104480
rect 106804 104416 106820 104480
rect 106884 104416 106900 104480
rect 106964 104416 106972 104480
rect 106652 103392 106972 104416
rect 106652 103328 106660 103392
rect 106724 103328 106740 103392
rect 106804 103328 106820 103392
rect 106884 103328 106900 103392
rect 106964 103328 106972 103392
rect 106652 102304 106972 103328
rect 106652 102240 106660 102304
rect 106724 102240 106740 102304
rect 106804 102240 106820 102304
rect 106884 102240 106900 102304
rect 106964 102240 106972 102304
rect 106652 101216 106972 102240
rect 106652 101152 106660 101216
rect 106724 101152 106740 101216
rect 106804 101152 106820 101216
rect 106884 101152 106900 101216
rect 106964 101152 106972 101216
rect 106652 100128 106972 101152
rect 106652 100064 106660 100128
rect 106724 100064 106740 100128
rect 106804 100064 106820 100128
rect 106884 100064 106900 100128
rect 106964 100064 106972 100128
rect 106652 99040 106972 100064
rect 106652 98976 106660 99040
rect 106724 98976 106740 99040
rect 106804 98976 106820 99040
rect 106884 98976 106900 99040
rect 106964 98976 106972 99040
rect 106652 98192 106972 98976
rect 106652 97956 106694 98192
rect 106930 97956 106972 98192
rect 106652 97952 106972 97956
rect 106652 97888 106660 97952
rect 106724 97888 106740 97952
rect 106804 97888 106820 97952
rect 106884 97888 106900 97952
rect 106964 97888 106972 97952
rect 106652 96864 106972 97888
rect 106652 96800 106660 96864
rect 106724 96800 106740 96864
rect 106804 96800 106820 96864
rect 106884 96800 106900 96864
rect 106964 96800 106972 96864
rect 106652 95776 106972 96800
rect 106652 95712 106660 95776
rect 106724 95712 106740 95776
rect 106804 95712 106820 95776
rect 106884 95712 106900 95776
rect 106964 95712 106972 95776
rect 106652 94688 106972 95712
rect 106652 94624 106660 94688
rect 106724 94624 106740 94688
rect 106804 94624 106820 94688
rect 106884 94624 106900 94688
rect 106964 94624 106972 94688
rect 106652 93600 106972 94624
rect 106652 93536 106660 93600
rect 106724 93536 106740 93600
rect 106804 93536 106820 93600
rect 106884 93536 106900 93600
rect 106964 93536 106972 93600
rect 106652 92512 106972 93536
rect 106652 92448 106660 92512
rect 106724 92448 106740 92512
rect 106804 92448 106820 92512
rect 106884 92448 106900 92512
rect 106964 92448 106972 92512
rect 106652 91424 106972 92448
rect 106652 91360 106660 91424
rect 106724 91360 106740 91424
rect 106804 91360 106820 91424
rect 106884 91360 106900 91424
rect 106964 91360 106972 91424
rect 106652 90336 106972 91360
rect 106652 90272 106660 90336
rect 106724 90272 106740 90336
rect 106804 90272 106820 90336
rect 106884 90272 106900 90336
rect 106964 90272 106972 90336
rect 106652 89248 106972 90272
rect 106652 89184 106660 89248
rect 106724 89184 106740 89248
rect 106804 89184 106820 89248
rect 106884 89184 106900 89248
rect 106964 89184 106972 89248
rect 106652 88160 106972 89184
rect 106652 88096 106660 88160
rect 106724 88096 106740 88160
rect 106804 88096 106820 88160
rect 106884 88096 106900 88160
rect 106964 88096 106972 88160
rect 106652 87072 106972 88096
rect 106652 87008 106660 87072
rect 106724 87008 106740 87072
rect 106804 87008 106820 87072
rect 106884 87008 106900 87072
rect 106964 87008 106972 87072
rect 106652 85984 106972 87008
rect 106652 85920 106660 85984
rect 106724 85920 106740 85984
rect 106804 85920 106820 85984
rect 106884 85920 106900 85984
rect 106964 85920 106972 85984
rect 106652 84896 106972 85920
rect 106652 84832 106660 84896
rect 106724 84832 106740 84896
rect 106804 84832 106820 84896
rect 106884 84832 106900 84896
rect 106964 84832 106972 84896
rect 106652 83808 106972 84832
rect 106652 83744 106660 83808
rect 106724 83744 106740 83808
rect 106804 83744 106820 83808
rect 106884 83744 106900 83808
rect 106964 83744 106972 83808
rect 106652 82720 106972 83744
rect 106652 82656 106660 82720
rect 106724 82656 106740 82720
rect 106804 82656 106820 82720
rect 106884 82656 106900 82720
rect 106964 82656 106972 82720
rect 106652 81632 106972 82656
rect 106652 81568 106660 81632
rect 106724 81568 106740 81632
rect 106804 81568 106820 81632
rect 106884 81568 106900 81632
rect 106964 81568 106972 81632
rect 106652 80544 106972 81568
rect 106652 80480 106660 80544
rect 106724 80480 106740 80544
rect 106804 80480 106820 80544
rect 106884 80480 106900 80544
rect 106964 80480 106972 80544
rect 106652 79456 106972 80480
rect 106652 79392 106660 79456
rect 106724 79392 106740 79456
rect 106804 79392 106820 79456
rect 106884 79392 106900 79456
rect 106964 79392 106972 79456
rect 106652 78368 106972 79392
rect 106652 78304 106660 78368
rect 106724 78304 106740 78368
rect 106804 78304 106820 78368
rect 106884 78304 106900 78368
rect 106964 78304 106972 78368
rect 106652 77280 106972 78304
rect 106652 77216 106660 77280
rect 106724 77216 106740 77280
rect 106804 77216 106820 77280
rect 106884 77216 106900 77280
rect 106964 77216 106972 77280
rect 106652 77200 106972 77216
rect 97028 76128 97036 76192
rect 97100 76128 97116 76192
rect 97180 76128 97196 76192
rect 97260 76128 97276 76192
rect 97340 76128 97348 76192
rect 97028 75104 97348 76128
rect 97028 75040 97036 75104
rect 97100 75040 97116 75104
rect 97180 75040 97196 75104
rect 97260 75040 97276 75104
rect 97340 75040 97348 75104
rect 97028 74016 97348 75040
rect 97028 73952 97036 74016
rect 97100 73952 97116 74016
rect 97180 73952 97196 74016
rect 97260 73952 97276 74016
rect 97340 73952 97348 74016
rect 97028 72928 97348 73952
rect 97028 72864 97036 72928
rect 97100 72864 97116 72928
rect 97180 72864 97196 72928
rect 97260 72864 97276 72928
rect 97340 72864 97348 72928
rect 97028 71840 97348 72864
rect 97028 71776 97036 71840
rect 97100 71776 97116 71840
rect 97180 71776 97196 71840
rect 97260 71776 97276 71840
rect 97340 71776 97348 71840
rect 97028 70752 97348 71776
rect 97028 70688 97036 70752
rect 97100 70688 97116 70752
rect 97180 70688 97196 70752
rect 97260 70688 97276 70752
rect 97340 70688 97348 70752
rect 97028 69664 97348 70688
rect 97028 69600 97036 69664
rect 97100 69600 97116 69664
rect 97180 69600 97196 69664
rect 97260 69600 97276 69664
rect 97340 69600 97348 69664
rect 97028 68576 97348 69600
rect 97028 68512 97036 68576
rect 97100 68512 97116 68576
rect 97180 68512 97196 68576
rect 97260 68512 97276 68576
rect 97340 68512 97348 68576
rect 97028 67556 97348 68512
rect 97028 67488 97070 67556
rect 97306 67488 97348 67556
rect 97028 67424 97036 67488
rect 97340 67424 97348 67488
rect 97028 67320 97070 67424
rect 97306 67320 97348 67424
rect 97028 66400 97348 67320
rect 97028 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97348 66400
rect 97028 65650 97348 66336
rect 105916 65856 106236 66416
rect 105916 65792 105924 65856
rect 105988 65792 106004 65856
rect 106068 65792 106084 65856
rect 106148 65792 106164 65856
rect 106228 65792 106236 65856
rect 105916 64768 106236 65792
rect 105916 64704 105924 64768
rect 105988 64704 106004 64768
rect 106068 64704 106084 64768
rect 106148 64704 106164 64768
rect 106228 64704 106236 64768
rect 87278 64230 87372 64290
rect 86144 63676 86204 64230
rect 87312 63676 87372 64230
rect 95857 64156 95923 64157
rect 95857 64092 95858 64156
rect 95922 64092 95923 64156
rect 95857 64091 95923 64092
rect 95860 63676 95920 64091
rect 105916 63680 106236 64704
rect 4868 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5188 63136
rect 4868 62048 5188 63072
rect 4868 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5188 62048
rect 4868 60960 5188 61984
rect 4868 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5188 60960
rect 4868 59872 5188 60896
rect 4868 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5188 59872
rect 4868 58784 5188 59808
rect 4868 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5188 58784
rect 4868 57696 5188 58720
rect 4868 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5188 57696
rect 4868 56608 5188 57632
rect 4868 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5188 56608
rect 4868 55520 5188 56544
rect 4868 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5188 55520
rect 4868 54432 5188 55456
rect 4868 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5188 54432
rect 4868 53344 5188 54368
rect 4868 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5188 53344
rect 4868 52256 5188 53280
rect 4868 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5188 52256
rect 4868 51168 5188 52192
rect 4868 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5188 51168
rect 4868 50080 5188 51104
rect 4868 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5188 50080
rect 4868 48992 5188 50016
rect 4868 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5188 48992
rect 4868 47904 5188 48928
rect 4868 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5188 47904
rect 4868 46816 5188 47840
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 105916 63616 105924 63680
rect 105988 63616 106004 63680
rect 106068 63616 106084 63680
rect 106148 63616 106164 63680
rect 106228 63616 106236 63680
rect 105916 62592 106236 63616
rect 105916 62528 105924 62592
rect 105988 62528 106004 62592
rect 106068 62528 106084 62592
rect 106148 62528 106164 62592
rect 106228 62528 106236 62592
rect 105916 61504 106236 62528
rect 105916 61440 105924 61504
rect 105988 61440 106004 61504
rect 106068 61440 106084 61504
rect 106148 61440 106164 61504
rect 106228 61440 106236 61504
rect 105916 60416 106236 61440
rect 105916 60352 105924 60416
rect 105988 60352 106004 60416
rect 106068 60352 106084 60416
rect 106148 60352 106164 60416
rect 106228 60352 106236 60416
rect 105916 59328 106236 60352
rect 105916 59264 105924 59328
rect 105988 59264 106004 59328
rect 106068 59264 106084 59328
rect 106148 59264 106164 59328
rect 106228 59264 106236 59328
rect 105916 58240 106236 59264
rect 105916 58176 105924 58240
rect 105988 58176 106004 58240
rect 106068 58176 106084 58240
rect 106148 58176 106164 58240
rect 106228 58176 106236 58240
rect 105916 57152 106236 58176
rect 105916 57088 105924 57152
rect 105988 57088 106004 57152
rect 106068 57088 106084 57152
rect 106148 57088 106164 57152
rect 106228 57088 106236 57152
rect 105916 56064 106236 57088
rect 105916 56000 105924 56064
rect 105988 56000 106004 56064
rect 106068 56000 106084 56064
rect 106148 56000 106164 56064
rect 106228 56000 106236 56064
rect 105916 54976 106236 56000
rect 105916 54912 105924 54976
rect 105988 54912 106004 54976
rect 106068 54912 106084 54976
rect 106148 54912 106164 54976
rect 106228 54912 106236 54976
rect 105916 53888 106236 54912
rect 105916 53824 105924 53888
rect 105988 53824 106004 53888
rect 106068 53824 106084 53888
rect 106148 53824 106164 53888
rect 106228 53824 106236 53888
rect 105916 52800 106236 53824
rect 105916 52736 105924 52800
rect 105988 52736 106004 52800
rect 106068 52736 106084 52800
rect 106148 52736 106164 52800
rect 106228 52736 106236 52800
rect 105916 51712 106236 52736
rect 105916 51648 105924 51712
rect 105988 51648 106004 51712
rect 106068 51648 106084 51712
rect 106148 51648 106164 51712
rect 106228 51648 106236 51712
rect 105916 50624 106236 51648
rect 105916 50560 105924 50624
rect 105988 50560 106004 50624
rect 106068 50560 106084 50624
rect 106148 50560 106164 50624
rect 106228 50560 106236 50624
rect 105916 49536 106236 50560
rect 105916 49472 105924 49536
rect 105988 49472 106004 49536
rect 106068 49472 106084 49536
rect 106148 49472 106164 49536
rect 106228 49472 106236 49536
rect 105916 48448 106236 49472
rect 105916 48384 105924 48448
rect 105988 48384 106004 48448
rect 106068 48384 106084 48448
rect 106148 48384 106164 48448
rect 106228 48384 106236 48448
rect 105916 47360 106236 48384
rect 105916 47296 105924 47360
rect 105988 47296 106004 47360
rect 106068 47296 106084 47360
rect 106148 47296 106164 47360
rect 106228 47296 106236 47360
rect 105916 46272 106236 47296
rect 105916 46208 105924 46272
rect 105988 46208 106004 46272
rect 106068 46208 106084 46272
rect 106148 46208 106164 46272
rect 106228 46208 106236 46272
rect 105916 45184 106236 46208
rect 105916 45120 105924 45184
rect 105988 45120 106004 45184
rect 106068 45120 106084 45184
rect 106148 45120 106164 45184
rect 106228 45120 106236 45184
rect 105916 44096 106236 45120
rect 105916 44032 105924 44096
rect 105988 44032 106004 44096
rect 106068 44032 106084 44096
rect 106148 44032 106164 44096
rect 106228 44032 106236 44096
rect 105916 43008 106236 44032
rect 105916 42944 105924 43008
rect 105988 42944 106004 43008
rect 106068 42944 106084 43008
rect 106148 42944 106164 43008
rect 106228 42944 106236 43008
rect 105916 41920 106236 42944
rect 105916 41856 105924 41920
rect 105988 41856 106004 41920
rect 106068 41856 106084 41920
rect 106148 41856 106164 41920
rect 106228 41856 106236 41920
rect 105916 40832 106236 41856
rect 105916 40768 105924 40832
rect 105988 40768 106004 40832
rect 106068 40768 106084 40832
rect 106148 40768 106164 40832
rect 106228 40768 106236 40832
rect 105916 39744 106236 40768
rect 105916 39680 105924 39744
rect 105988 39680 106004 39744
rect 106068 39680 106084 39744
rect 106148 39680 106164 39744
rect 106228 39680 106236 39744
rect 105916 38656 106236 39680
rect 105916 38592 105924 38656
rect 105988 38592 106004 38656
rect 106068 38592 106084 38656
rect 106148 38592 106164 38656
rect 106228 38592 106236 38656
rect 105916 37568 106236 38592
rect 105916 37504 105924 37568
rect 105988 37504 106004 37568
rect 106068 37504 106084 37568
rect 106148 37504 106164 37568
rect 106228 37504 106236 37568
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 10696 36920 11044 36962
rect 10696 36684 10752 36920
rect 10988 36684 11044 36920
rect 10696 36642 11044 36684
rect 100936 36920 101284 36962
rect 100936 36684 100992 36920
rect 101228 36684 101284 36920
rect 100936 36642 101284 36684
rect 105916 36480 106236 37504
rect 105916 36416 105924 36480
rect 105988 36416 106004 36480
rect 106068 36416 106084 36480
rect 106148 36416 106164 36480
rect 106228 36416 106236 36480
rect 10000 36260 10348 36302
rect 10000 36024 10056 36260
rect 10292 36024 10348 36260
rect 10000 35982 10348 36024
rect 101632 36260 101980 36302
rect 101632 36024 101688 36260
rect 101924 36024 101980 36260
rect 101632 35982 101980 36024
rect 105916 36260 106236 36416
rect 105916 36024 105958 36260
rect 106194 36024 106236 36260
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 105916 35392 106236 36024
rect 105916 35328 105924 35392
rect 105988 35328 106004 35392
rect 106068 35328 106084 35392
rect 106148 35328 106164 35392
rect 106228 35328 106236 35392
rect 105916 34304 106236 35328
rect 105916 34240 105924 34304
rect 105988 34240 106004 34304
rect 106068 34240 106084 34304
rect 106148 34240 106164 34304
rect 106228 34240 106236 34304
rect 105916 33216 106236 34240
rect 105916 33152 105924 33216
rect 105988 33152 106004 33216
rect 106068 33152 106084 33216
rect 106148 33152 106164 33216
rect 106228 33152 106236 33216
rect 105916 32128 106236 33152
rect 105916 32064 105924 32128
rect 105988 32064 106004 32128
rect 106068 32064 106084 32128
rect 106148 32064 106164 32128
rect 106228 32064 106236 32128
rect 105916 31040 106236 32064
rect 105916 30976 105924 31040
rect 105988 30976 106004 31040
rect 106068 30976 106084 31040
rect 106148 30976 106164 31040
rect 106228 30976 106236 31040
rect 105916 29952 106236 30976
rect 105916 29888 105924 29952
rect 105988 29888 106004 29952
rect 106068 29888 106084 29952
rect 106148 29888 106164 29952
rect 106228 29888 106236 29952
rect 105916 28864 106236 29888
rect 105916 28800 105924 28864
rect 105988 28800 106004 28864
rect 106068 28800 106084 28864
rect 106148 28800 106164 28864
rect 106228 28800 106236 28864
rect 105916 27776 106236 28800
rect 105916 27712 105924 27776
rect 105988 27712 106004 27776
rect 106068 27712 106084 27776
rect 106148 27712 106164 27776
rect 106228 27712 106236 27776
rect 105916 26688 106236 27712
rect 105916 26624 105924 26688
rect 105988 26624 106004 26688
rect 106068 26624 106084 26688
rect 106148 26624 106164 26688
rect 106228 26624 106236 26688
rect 105916 25600 106236 26624
rect 105916 25536 105924 25600
rect 105988 25536 106004 25600
rect 106068 25536 106084 25600
rect 106148 25536 106164 25600
rect 106228 25536 106236 25600
rect 105916 24512 106236 25536
rect 105916 24448 105924 24512
rect 105988 24448 106004 24512
rect 106068 24448 106084 24512
rect 106148 24448 106164 24512
rect 106228 24448 106236 24512
rect 105916 23424 106236 24448
rect 105916 23360 105924 23424
rect 105988 23360 106004 23424
rect 106068 23360 106084 23424
rect 106148 23360 106164 23424
rect 106228 23360 106236 23424
rect 105916 22336 106236 23360
rect 105916 22272 105924 22336
rect 105988 22272 106004 22336
rect 106068 22272 106084 22336
rect 106148 22272 106164 22336
rect 106228 22272 106236 22336
rect 105916 21248 106236 22272
rect 105916 21184 105924 21248
rect 105988 21184 106004 21248
rect 106068 21184 106084 21248
rect 106148 21184 106164 21248
rect 106228 21184 106236 21248
rect 105916 20160 106236 21184
rect 105916 20096 105924 20160
rect 105988 20096 106004 20160
rect 106068 20096 106084 20160
rect 106148 20096 106164 20160
rect 106228 20096 106236 20160
rect 105916 19072 106236 20096
rect 105916 19008 105924 19072
rect 105988 19008 106004 19072
rect 106068 19008 106084 19072
rect 106148 19008 106164 19072
rect 106228 19008 106236 19072
rect 105916 17984 106236 19008
rect 105916 17920 105924 17984
rect 105988 17920 106004 17984
rect 106068 17920 106084 17984
rect 106148 17920 106164 17984
rect 106228 17920 106236 17984
rect 105916 16896 106236 17920
rect 105916 16832 105924 16896
rect 105988 16832 106004 16896
rect 106068 16832 106084 16896
rect 106148 16832 106164 16896
rect 106228 16832 106236 16896
rect 105916 15808 106236 16832
rect 105916 15744 105924 15808
rect 105988 15744 106004 15808
rect 106068 15744 106084 15808
rect 106148 15744 106164 15808
rect 106228 15744 106236 15808
rect 105916 14720 106236 15744
rect 105916 14656 105924 14720
rect 105988 14656 106004 14720
rect 106068 14656 106084 14720
rect 106148 14656 106164 14720
rect 106228 14656 106236 14720
rect 105916 13632 106236 14656
rect 105916 13568 105924 13632
rect 105988 13568 106004 13632
rect 106068 13568 106084 13632
rect 106148 13568 106164 13632
rect 106228 13568 106236 13632
rect 105916 12544 106236 13568
rect 105916 12480 105924 12544
rect 105988 12480 106004 12544
rect 106068 12480 106084 12544
rect 106148 12480 106164 12544
rect 106228 12480 106236 12544
rect 105916 11456 106236 12480
rect 105916 11392 105924 11456
rect 105988 11392 106004 11456
rect 106068 11392 106084 11456
rect 106148 11392 106164 11456
rect 106228 11392 106236 11456
rect 105916 10368 106236 11392
rect 105916 10304 105924 10368
rect 105988 10304 106004 10368
rect 106068 10304 106084 10368
rect 106148 10304 106164 10368
rect 106228 10304 106236 10368
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 16060 9621 16120 10038
rect 23440 9757 23500 10038
rect 23437 9756 23503 9757
rect 23437 9692 23438 9756
rect 23502 9692 23503 9756
rect 23437 9691 23503 9692
rect 24626 9621 24686 10038
rect 25776 9757 25836 10038
rect 25773 9756 25839 9757
rect 25773 9692 25774 9756
rect 25838 9692 25839 9756
rect 25773 9691 25839 9692
rect 16057 9620 16123 9621
rect 16057 9556 16058 9620
rect 16122 9556 16123 9620
rect 16057 9555 16123 9556
rect 24623 9620 24689 9621
rect 24623 9556 24624 9620
rect 24688 9556 24689 9620
rect 24623 9555 24689 9556
rect 26926 8941 26986 10038
rect 28122 9757 28182 10038
rect 29280 9757 29340 10038
rect 30448 9757 30508 10038
rect 28119 9756 28185 9757
rect 28119 9692 28120 9756
rect 28184 9692 28185 9756
rect 28119 9691 28185 9692
rect 29277 9756 29343 9757
rect 29277 9692 29278 9756
rect 29342 9692 29343 9756
rect 29277 9691 29343 9692
rect 30445 9756 30511 9757
rect 30445 9692 30446 9756
rect 30510 9692 30511 9756
rect 31618 9754 31678 10038
rect 32784 9754 32844 10038
rect 33952 9754 34012 10038
rect 35120 9890 35180 10038
rect 36288 9890 36348 10038
rect 37456 9890 37516 10038
rect 35120 9830 35266 9890
rect 36288 9830 36370 9890
rect 31618 9694 31770 9754
rect 32784 9694 32874 9754
rect 30445 9691 30511 9692
rect 26923 8940 26989 8941
rect 26923 8876 26924 8940
rect 26988 8876 26989 8940
rect 26923 8875 26989 8876
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 31710 8261 31770 9694
rect 32814 8261 32874 9694
rect 33918 9694 34012 9754
rect 33918 8261 33978 9694
rect 35206 8261 35266 9830
rect 36310 8261 36370 9830
rect 37414 9830 37516 9890
rect 38624 9890 38684 10038
rect 38624 9830 38762 9890
rect 37414 8261 37474 9830
rect 38702 8261 38762 9830
rect 31707 8260 31773 8261
rect 31707 8196 31708 8260
rect 31772 8196 31773 8260
rect 31707 8195 31773 8196
rect 32811 8260 32877 8261
rect 32811 8196 32812 8260
rect 32876 8196 32877 8260
rect 32811 8195 32877 8196
rect 33915 8260 33981 8261
rect 33915 8196 33916 8260
rect 33980 8196 33981 8260
rect 33915 8195 33981 8196
rect 35203 8260 35269 8261
rect 35203 8196 35204 8260
rect 35268 8196 35269 8260
rect 35203 8195 35269 8196
rect 36307 8260 36373 8261
rect 36307 8196 36308 8260
rect 36372 8196 36373 8260
rect 36307 8195 36373 8196
rect 37411 8260 37477 8261
rect 37411 8196 37412 8260
rect 37476 8196 37477 8260
rect 37411 8195 37477 8196
rect 38699 8260 38765 8261
rect 38699 8196 38700 8260
rect 38764 8196 38765 8260
rect 38699 8195 38765 8196
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 7104 35248 7880
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 7648 35908 8064
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 39806 4589 39866 10038
rect 40960 9890 41020 10038
rect 40910 9830 41020 9890
rect 42128 9890 42188 10038
rect 42128 9830 42258 9890
rect 40910 8261 40970 9830
rect 42198 8261 42258 9830
rect 43302 8261 43362 10038
rect 90529 9757 90589 10038
rect 90526 9756 90592 9757
rect 90526 9692 90527 9756
rect 90591 9692 90592 9756
rect 90526 9691 90592 9692
rect 90682 9621 90742 10038
rect 90816 9890 90876 10038
rect 90816 9830 91018 9890
rect 90958 9757 91018 9830
rect 90955 9756 91021 9757
rect 90955 9692 90956 9756
rect 91020 9692 91021 9756
rect 90955 9691 91021 9692
rect 90679 9620 90745 9621
rect 90679 9556 90680 9620
rect 90744 9556 90745 9620
rect 90679 9555 90745 9556
rect 105916 9280 106236 10304
rect 105916 9216 105924 9280
rect 105988 9216 106004 9280
rect 106068 9216 106084 9280
rect 106148 9216 106164 9280
rect 106228 9216 106236 9280
rect 40907 8260 40973 8261
rect 40907 8196 40908 8260
rect 40972 8196 40973 8260
rect 40907 8195 40973 8196
rect 42195 8260 42261 8261
rect 42195 8196 42196 8260
rect 42260 8196 42261 8260
rect 42195 8195 42261 8196
rect 43299 8260 43365 8261
rect 43299 8196 43300 8260
rect 43364 8196 43365 8260
rect 43299 8195 43365 8196
rect 105916 8192 106236 9216
rect 105916 8128 105924 8192
rect 105988 8128 106004 8192
rect 106068 8128 106084 8192
rect 106148 8128 106164 8192
rect 106228 8128 106236 8192
rect 65648 7104 65968 8064
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 5624 65968 5952
rect 65648 5388 65690 5624
rect 65926 5388 65968 5624
rect 65648 4928 65968 5388
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 39803 4588 39869 4589
rect 39803 4524 39804 4588
rect 39868 4524 39869 4588
rect 39803 4523 39869 4524
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
rect 66308 7648 66628 8064
rect 66308 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66628 7648
rect 66308 6560 66628 7584
rect 66308 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66628 6560
rect 66308 6284 66628 6496
rect 66308 6048 66350 6284
rect 66586 6048 66628 6284
rect 66308 5472 66628 6048
rect 66308 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66628 5472
rect 66308 4384 66628 5408
rect 66308 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66628 4384
rect 66308 3296 66628 4320
rect 66308 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66628 3296
rect 66308 2208 66628 3232
rect 66308 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66628 2208
rect 66308 2128 66628 2144
rect 96368 7104 96688 8064
rect 96368 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96688 7104
rect 96368 6016 96688 7040
rect 96368 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96688 6016
rect 96368 5624 96688 5952
rect 96368 5388 96410 5624
rect 96646 5388 96688 5624
rect 96368 4928 96688 5388
rect 96368 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96688 4928
rect 96368 3840 96688 4864
rect 96368 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96688 3840
rect 96368 2752 96688 3776
rect 96368 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96688 2752
rect 96368 2128 96688 2688
rect 97028 7648 97348 8064
rect 97028 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97348 7648
rect 97028 6560 97348 7584
rect 105916 7104 106236 8128
rect 105916 7040 105924 7104
rect 105988 7040 106004 7104
rect 106068 7040 106084 7104
rect 106148 7040 106164 7104
rect 106228 7040 106236 7104
rect 105916 7024 106236 7040
rect 106652 66400 106972 66416
rect 106652 66336 106660 66400
rect 106724 66336 106740 66400
rect 106804 66336 106820 66400
rect 106884 66336 106900 66400
rect 106964 66336 106972 66400
rect 106652 65312 106972 66336
rect 106652 65248 106660 65312
rect 106724 65248 106740 65312
rect 106804 65248 106820 65312
rect 106884 65248 106900 65312
rect 106964 65248 106972 65312
rect 106652 64224 106972 65248
rect 106652 64160 106660 64224
rect 106724 64160 106740 64224
rect 106804 64160 106820 64224
rect 106884 64160 106900 64224
rect 106964 64160 106972 64224
rect 106652 63136 106972 64160
rect 106652 63072 106660 63136
rect 106724 63072 106740 63136
rect 106804 63072 106820 63136
rect 106884 63072 106900 63136
rect 106964 63072 106972 63136
rect 106652 62048 106972 63072
rect 106652 61984 106660 62048
rect 106724 61984 106740 62048
rect 106804 61984 106820 62048
rect 106884 61984 106900 62048
rect 106964 61984 106972 62048
rect 106652 60960 106972 61984
rect 106652 60896 106660 60960
rect 106724 60896 106740 60960
rect 106804 60896 106820 60960
rect 106884 60896 106900 60960
rect 106964 60896 106972 60960
rect 106652 59872 106972 60896
rect 106652 59808 106660 59872
rect 106724 59808 106740 59872
rect 106804 59808 106820 59872
rect 106884 59808 106900 59872
rect 106964 59808 106972 59872
rect 106652 58784 106972 59808
rect 106652 58720 106660 58784
rect 106724 58720 106740 58784
rect 106804 58720 106820 58784
rect 106884 58720 106900 58784
rect 106964 58720 106972 58784
rect 106652 57696 106972 58720
rect 106652 57632 106660 57696
rect 106724 57632 106740 57696
rect 106804 57632 106820 57696
rect 106884 57632 106900 57696
rect 106964 57632 106972 57696
rect 106652 56608 106972 57632
rect 106652 56544 106660 56608
rect 106724 56544 106740 56608
rect 106804 56544 106820 56608
rect 106884 56544 106900 56608
rect 106964 56544 106972 56608
rect 106652 55520 106972 56544
rect 106652 55456 106660 55520
rect 106724 55456 106740 55520
rect 106804 55456 106820 55520
rect 106884 55456 106900 55520
rect 106964 55456 106972 55520
rect 106652 54432 106972 55456
rect 106652 54368 106660 54432
rect 106724 54368 106740 54432
rect 106804 54368 106820 54432
rect 106884 54368 106900 54432
rect 106964 54368 106972 54432
rect 106652 53344 106972 54368
rect 106652 53280 106660 53344
rect 106724 53280 106740 53344
rect 106804 53280 106820 53344
rect 106884 53280 106900 53344
rect 106964 53280 106972 53344
rect 106652 52256 106972 53280
rect 106652 52192 106660 52256
rect 106724 52192 106740 52256
rect 106804 52192 106820 52256
rect 106884 52192 106900 52256
rect 106964 52192 106972 52256
rect 106652 51168 106972 52192
rect 106652 51104 106660 51168
rect 106724 51104 106740 51168
rect 106804 51104 106820 51168
rect 106884 51104 106900 51168
rect 106964 51104 106972 51168
rect 106652 50080 106972 51104
rect 106652 50016 106660 50080
rect 106724 50016 106740 50080
rect 106804 50016 106820 50080
rect 106884 50016 106900 50080
rect 106964 50016 106972 50080
rect 106652 48992 106972 50016
rect 106652 48928 106660 48992
rect 106724 48928 106740 48992
rect 106804 48928 106820 48992
rect 106884 48928 106900 48992
rect 106964 48928 106972 48992
rect 106652 47904 106972 48928
rect 106652 47840 106660 47904
rect 106724 47840 106740 47904
rect 106804 47840 106820 47904
rect 106884 47840 106900 47904
rect 106964 47840 106972 47904
rect 106652 46816 106972 47840
rect 106652 46752 106660 46816
rect 106724 46752 106740 46816
rect 106804 46752 106820 46816
rect 106884 46752 106900 46816
rect 106964 46752 106972 46816
rect 106652 45728 106972 46752
rect 106652 45664 106660 45728
rect 106724 45664 106740 45728
rect 106804 45664 106820 45728
rect 106884 45664 106900 45728
rect 106964 45664 106972 45728
rect 106652 44640 106972 45664
rect 106652 44576 106660 44640
rect 106724 44576 106740 44640
rect 106804 44576 106820 44640
rect 106884 44576 106900 44640
rect 106964 44576 106972 44640
rect 106652 43552 106972 44576
rect 106652 43488 106660 43552
rect 106724 43488 106740 43552
rect 106804 43488 106820 43552
rect 106884 43488 106900 43552
rect 106964 43488 106972 43552
rect 106652 42464 106972 43488
rect 106652 42400 106660 42464
rect 106724 42400 106740 42464
rect 106804 42400 106820 42464
rect 106884 42400 106900 42464
rect 106964 42400 106972 42464
rect 106652 41376 106972 42400
rect 106652 41312 106660 41376
rect 106724 41312 106740 41376
rect 106804 41312 106820 41376
rect 106884 41312 106900 41376
rect 106964 41312 106972 41376
rect 106652 40288 106972 41312
rect 106652 40224 106660 40288
rect 106724 40224 106740 40288
rect 106804 40224 106820 40288
rect 106884 40224 106900 40288
rect 106964 40224 106972 40288
rect 106652 39200 106972 40224
rect 106652 39136 106660 39200
rect 106724 39136 106740 39200
rect 106804 39136 106820 39200
rect 106884 39136 106900 39200
rect 106964 39136 106972 39200
rect 106652 38112 106972 39136
rect 106652 38048 106660 38112
rect 106724 38048 106740 38112
rect 106804 38048 106820 38112
rect 106884 38048 106900 38112
rect 106964 38048 106972 38112
rect 106652 37024 106972 38048
rect 106652 36960 106660 37024
rect 106724 36960 106740 37024
rect 106804 36960 106820 37024
rect 106884 36960 106900 37024
rect 106964 36960 106972 37024
rect 106652 36920 106972 36960
rect 106652 36684 106694 36920
rect 106930 36684 106972 36920
rect 106652 35936 106972 36684
rect 106652 35872 106660 35936
rect 106724 35872 106740 35936
rect 106804 35872 106820 35936
rect 106884 35872 106900 35936
rect 106964 35872 106972 35936
rect 106652 34848 106972 35872
rect 106652 34784 106660 34848
rect 106724 34784 106740 34848
rect 106804 34784 106820 34848
rect 106884 34784 106900 34848
rect 106964 34784 106972 34848
rect 106652 33760 106972 34784
rect 106652 33696 106660 33760
rect 106724 33696 106740 33760
rect 106804 33696 106820 33760
rect 106884 33696 106900 33760
rect 106964 33696 106972 33760
rect 106652 32672 106972 33696
rect 106652 32608 106660 32672
rect 106724 32608 106740 32672
rect 106804 32608 106820 32672
rect 106884 32608 106900 32672
rect 106964 32608 106972 32672
rect 106652 31584 106972 32608
rect 106652 31520 106660 31584
rect 106724 31520 106740 31584
rect 106804 31520 106820 31584
rect 106884 31520 106900 31584
rect 106964 31520 106972 31584
rect 106652 30496 106972 31520
rect 106652 30432 106660 30496
rect 106724 30432 106740 30496
rect 106804 30432 106820 30496
rect 106884 30432 106900 30496
rect 106964 30432 106972 30496
rect 106652 29408 106972 30432
rect 106652 29344 106660 29408
rect 106724 29344 106740 29408
rect 106804 29344 106820 29408
rect 106884 29344 106900 29408
rect 106964 29344 106972 29408
rect 106652 28320 106972 29344
rect 106652 28256 106660 28320
rect 106724 28256 106740 28320
rect 106804 28256 106820 28320
rect 106884 28256 106900 28320
rect 106964 28256 106972 28320
rect 106652 27232 106972 28256
rect 106652 27168 106660 27232
rect 106724 27168 106740 27232
rect 106804 27168 106820 27232
rect 106884 27168 106900 27232
rect 106964 27168 106972 27232
rect 106652 26144 106972 27168
rect 106652 26080 106660 26144
rect 106724 26080 106740 26144
rect 106804 26080 106820 26144
rect 106884 26080 106900 26144
rect 106964 26080 106972 26144
rect 106652 25056 106972 26080
rect 106652 24992 106660 25056
rect 106724 24992 106740 25056
rect 106804 24992 106820 25056
rect 106884 24992 106900 25056
rect 106964 24992 106972 25056
rect 106652 23968 106972 24992
rect 106652 23904 106660 23968
rect 106724 23904 106740 23968
rect 106804 23904 106820 23968
rect 106884 23904 106900 23968
rect 106964 23904 106972 23968
rect 106652 22880 106972 23904
rect 106652 22816 106660 22880
rect 106724 22816 106740 22880
rect 106804 22816 106820 22880
rect 106884 22816 106900 22880
rect 106964 22816 106972 22880
rect 106652 21792 106972 22816
rect 106652 21728 106660 21792
rect 106724 21728 106740 21792
rect 106804 21728 106820 21792
rect 106884 21728 106900 21792
rect 106964 21728 106972 21792
rect 106652 20704 106972 21728
rect 106652 20640 106660 20704
rect 106724 20640 106740 20704
rect 106804 20640 106820 20704
rect 106884 20640 106900 20704
rect 106964 20640 106972 20704
rect 106652 19616 106972 20640
rect 106652 19552 106660 19616
rect 106724 19552 106740 19616
rect 106804 19552 106820 19616
rect 106884 19552 106900 19616
rect 106964 19552 106972 19616
rect 106652 18528 106972 19552
rect 106652 18464 106660 18528
rect 106724 18464 106740 18528
rect 106804 18464 106820 18528
rect 106884 18464 106900 18528
rect 106964 18464 106972 18528
rect 106652 17440 106972 18464
rect 106652 17376 106660 17440
rect 106724 17376 106740 17440
rect 106804 17376 106820 17440
rect 106884 17376 106900 17440
rect 106964 17376 106972 17440
rect 106652 16352 106972 17376
rect 106652 16288 106660 16352
rect 106724 16288 106740 16352
rect 106804 16288 106820 16352
rect 106884 16288 106900 16352
rect 106964 16288 106972 16352
rect 106652 15264 106972 16288
rect 106652 15200 106660 15264
rect 106724 15200 106740 15264
rect 106804 15200 106820 15264
rect 106884 15200 106900 15264
rect 106964 15200 106972 15264
rect 106652 14176 106972 15200
rect 106652 14112 106660 14176
rect 106724 14112 106740 14176
rect 106804 14112 106820 14176
rect 106884 14112 106900 14176
rect 106964 14112 106972 14176
rect 106652 13088 106972 14112
rect 106652 13024 106660 13088
rect 106724 13024 106740 13088
rect 106804 13024 106820 13088
rect 106884 13024 106900 13088
rect 106964 13024 106972 13088
rect 106652 12000 106972 13024
rect 106652 11936 106660 12000
rect 106724 11936 106740 12000
rect 106804 11936 106820 12000
rect 106884 11936 106900 12000
rect 106964 11936 106972 12000
rect 106652 10912 106972 11936
rect 106652 10848 106660 10912
rect 106724 10848 106740 10912
rect 106804 10848 106820 10912
rect 106884 10848 106900 10912
rect 106964 10848 106972 10912
rect 106652 9824 106972 10848
rect 106652 9760 106660 9824
rect 106724 9760 106740 9824
rect 106804 9760 106820 9824
rect 106884 9760 106900 9824
rect 106964 9760 106972 9824
rect 106652 8736 106972 9760
rect 106652 8672 106660 8736
rect 106724 8672 106740 8736
rect 106804 8672 106820 8736
rect 106884 8672 106900 8736
rect 106964 8672 106972 8736
rect 106652 7648 106972 8672
rect 106652 7584 106660 7648
rect 106724 7584 106740 7648
rect 106804 7584 106820 7648
rect 106884 7584 106900 7648
rect 106964 7584 106972 7648
rect 106652 7024 106972 7584
rect 97028 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97348 6560
rect 97028 6284 97348 6496
rect 97028 6048 97070 6284
rect 97306 6048 97348 6284
rect 97028 5472 97348 6048
rect 97028 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97348 5472
rect 97028 4384 97348 5408
rect 97028 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97348 4384
rect 97028 3296 97348 4320
rect 97028 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97348 3296
rect 97028 2208 97348 3232
rect 97028 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97348 2208
rect 97028 2128 97348 2144
<< via4 >>
rect 4250 140982 4486 141218
rect 4250 127932 4486 128168
rect 4250 97408 4486 97532
rect 4250 97344 4280 97408
rect 4280 97344 4296 97408
rect 4296 97344 4360 97408
rect 4360 97344 4376 97408
rect 4376 97344 4440 97408
rect 4440 97344 4456 97408
rect 4456 97344 4486 97408
rect 4250 97296 4486 97344
rect 4250 66880 4280 66896
rect 4280 66880 4296 66896
rect 4296 66880 4360 66896
rect 4360 66880 4376 66896
rect 4376 66880 4440 66896
rect 4440 66880 4456 66896
rect 4456 66880 4486 66896
rect 4250 66660 4486 66880
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 141662 5146 141898
rect 34970 140982 35206 141218
rect 35630 141662 35866 141898
rect 65690 140982 65926 141218
rect 66350 141662 66586 141898
rect 96410 140982 96646 141218
rect 97070 141662 97306 141898
rect 4910 128592 5146 128828
rect 10752 128592 10988 128828
rect 100992 128592 101228 128828
rect 10056 127932 10292 128168
rect 101688 127932 101924 128168
rect 105958 127932 106194 128168
rect 4910 97956 5146 98192
rect 10752 97956 10988 98192
rect 100992 97956 101228 98192
rect 10056 97296 10292 97532
rect 101688 97296 101924 97532
rect 105958 97408 106194 97532
rect 105958 97344 105988 97408
rect 105988 97344 106004 97408
rect 106004 97344 106068 97408
rect 106068 97344 106084 97408
rect 106084 97344 106148 97408
rect 106148 97344 106164 97408
rect 106164 97344 106194 97408
rect 105958 97296 106194 97344
rect 4910 67488 5146 67556
rect 4910 67424 4940 67488
rect 4940 67424 4956 67488
rect 4956 67424 5020 67488
rect 5020 67424 5036 67488
rect 5036 67424 5100 67488
rect 5100 67424 5116 67488
rect 5116 67424 5146 67488
rect 4910 67320 5146 67424
rect 34970 66880 35000 66896
rect 35000 66880 35016 66896
rect 35016 66880 35080 66896
rect 35080 66880 35096 66896
rect 35096 66880 35160 66896
rect 35160 66880 35176 66896
rect 35176 66880 35206 66896
rect 34970 66660 35206 66880
rect 35630 67488 35866 67556
rect 35630 67424 35660 67488
rect 35660 67424 35676 67488
rect 35676 67424 35740 67488
rect 35740 67424 35756 67488
rect 35756 67424 35820 67488
rect 35820 67424 35836 67488
rect 35836 67424 35866 67488
rect 35630 67320 35866 67424
rect 65690 66880 65720 66896
rect 65720 66880 65736 66896
rect 65736 66880 65800 66896
rect 65800 66880 65816 66896
rect 65816 66880 65880 66896
rect 65880 66880 65896 66896
rect 65896 66880 65926 66896
rect 65690 66660 65926 66880
rect 66350 67488 66586 67556
rect 66350 67424 66380 67488
rect 66380 67424 66396 67488
rect 66396 67424 66460 67488
rect 66460 67424 66476 67488
rect 66476 67424 66540 67488
rect 66540 67424 66556 67488
rect 66556 67424 66586 67488
rect 66350 67320 66586 67424
rect 96410 66880 96440 66896
rect 96440 66880 96456 66896
rect 96456 66880 96520 66896
rect 96520 66880 96536 66896
rect 96536 66880 96600 66896
rect 96600 66880 96616 66896
rect 96616 66880 96646 66896
rect 96410 66660 96646 66880
rect 106694 128592 106930 128828
rect 106694 97956 106930 98192
rect 97070 67488 97306 67556
rect 97070 67424 97100 67488
rect 97100 67424 97116 67488
rect 97116 67424 97180 67488
rect 97180 67424 97196 67488
rect 97196 67424 97260 67488
rect 97260 67424 97276 67488
rect 97276 67424 97306 67488
rect 97070 67320 97306 67424
rect 4910 36684 5146 36920
rect 10752 36684 10988 36920
rect 100992 36684 101228 36920
rect 10056 36024 10292 36260
rect 101688 36024 101924 36260
rect 105958 36024 106194 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 6048 35866 6284
rect 65690 5388 65926 5624
rect 66350 6048 66586 6284
rect 96410 5388 96646 5624
rect 106694 36684 106930 36920
rect 97070 6048 97306 6284
<< metal5 >>
rect 4208 141898 108884 141940
rect 4208 141662 4910 141898
rect 5146 141662 35630 141898
rect 35866 141662 66350 141898
rect 66586 141662 97070 141898
rect 97306 141662 108884 141898
rect 4208 141620 108884 141662
rect 4208 141218 108884 141260
rect 4208 140982 4250 141218
rect 4486 140982 34970 141218
rect 35206 140982 65690 141218
rect 65926 140982 96410 141218
rect 96646 140982 108884 141218
rect 4208 140940 108884 140982
rect 1056 128828 108884 128870
rect 1056 128592 4910 128828
rect 5146 128592 10752 128828
rect 10988 128592 100992 128828
rect 101228 128592 106694 128828
rect 106930 128592 108884 128828
rect 1056 128550 108884 128592
rect 1056 128168 108884 128210
rect 1056 127932 4250 128168
rect 4486 127932 10056 128168
rect 10292 127932 101688 128168
rect 101924 127932 105958 128168
rect 106194 127932 108884 128168
rect 1056 127890 108884 127932
rect 1056 98192 108884 98234
rect 1056 97956 4910 98192
rect 5146 97956 10752 98192
rect 10988 97956 100992 98192
rect 101228 97956 106694 98192
rect 106930 97956 108884 98192
rect 1056 97914 108884 97956
rect 1056 97532 108884 97574
rect 1056 97296 4250 97532
rect 4486 97296 10056 97532
rect 10292 97296 101688 97532
rect 101924 97296 105958 97532
rect 106194 97296 108884 97532
rect 1056 97254 108884 97296
rect 1056 67556 108884 67598
rect 1056 67320 4910 67556
rect 5146 67320 35630 67556
rect 35866 67320 66350 67556
rect 66586 67320 97070 67556
rect 97306 67320 108884 67556
rect 1056 67278 108884 67320
rect 1056 66896 108884 66938
rect 1056 66660 4250 66896
rect 4486 66660 34970 66896
rect 35206 66660 65690 66896
rect 65926 66660 96410 66896
rect 96646 66660 108884 66896
rect 1056 66618 108884 66660
rect 1056 36920 108884 36962
rect 1056 36684 4910 36920
rect 5146 36684 10752 36920
rect 10988 36684 100992 36920
rect 101228 36684 106694 36920
rect 106930 36684 108884 36920
rect 1056 36642 108884 36684
rect 1056 36260 108884 36302
rect 1056 36024 4250 36260
rect 4486 36024 10056 36260
rect 10292 36024 101688 36260
rect 101924 36024 105958 36260
rect 106194 36024 108884 36260
rect 1056 35982 108884 36024
rect 1056 6284 108884 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 66350 6284
rect 66586 6048 97070 6284
rect 97306 6048 108884 6284
rect 1056 6006 108884 6048
rect 1056 5624 108884 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 65690 5624
rect 65926 5388 96410 5624
rect 96646 5388 108884 5624
rect 1056 5346 108884 5388
use sky130_fd_sc_hd__inv_2  _061_
timestamp 1
transform -1 0 84088 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1
transform 1 0 83628 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _063_
timestamp 1
transform 1 0 30728 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _064_
timestamp 1
transform 1 0 32660 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _065_
timestamp 1
transform 1 0 34868 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _066_
timestamp 1
transform 1 0 37260 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _067_
timestamp 1
transform 1 0 39836 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _068_
timestamp 1
transform 1 0 42412 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _069_
timestamp 1
transform -1 0 61640 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _070_
timestamp 1
transform -1 0 63848 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _071_
timestamp 1
transform -1 0 66424 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _072_
timestamp 1
transform -1 0 69000 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _073_
timestamp 1
transform -1 0 70288 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _074_
timestamp 1
transform -1 0 72036 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _075_
timestamp 1
transform -1 0 74520 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _076_
timestamp 1
transform -1 0 76728 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _077_
timestamp 1
transform -1 0 79304 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _078_
timestamp 1
transform -1 0 80960 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _079_
timestamp 1
transform -1 0 86848 0 1 77248
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _080_
timestamp 1
transform -1 0 90896 0 1 75072
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _081_
timestamp 1
transform -1 0 90344 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _082_
timestamp 1
transform 1 0 90068 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _083_
timestamp 1
transform 1 0 91540 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _084_
timestamp 1
transform 1 0 92184 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _085_
timestamp 1
transform -1 0 91172 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _086_
timestamp 1
transform -1 0 89608 0 -1 67456
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _087_
timestamp 1
transform -1 0 91816 0 -1 66368
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _088_
timestamp 1
transform -1 0 90620 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _089_
timestamp 1
transform 1 0 90988 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _090_
timestamp 1
transform -1 0 90620 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _091_
timestamp 1
transform -1 0 89976 0 -1 66368
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _092_
timestamp 1
transform -1 0 88688 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _093_
timestamp 1
transform 1 0 88780 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _094_
timestamp 1
transform -1 0 85744 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _095_
timestamp 1
transform -1 0 78016 0 -1 70720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1
transform 1 0 85468 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 1
transform 1 0 86204 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098_
timestamp 1
transform 1 0 85652 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1
transform 1 0 88044 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1
transform 1 0 88412 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1
transform 1 0 89700 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1
transform 1 0 91632 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1
transform -1 0 81696 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1
transform 1 0 82708 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105_
timestamp 1
transform 1 0 87860 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1
transform 1 0 88964 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp 1
transform 1 0 86572 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1
transform 1 0 86204 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _109_
timestamp 1
transform 1 0 84364 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp 1
transform -1 0 83996 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 1
transform 1 0 74060 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1
transform -1 0 27784 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113_
timestamp 1
transform -1 0 29164 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 1
transform -1 0 30452 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1
transform -1 0 31188 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 1
transform -1 0 31740 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 1
transform -1 0 32476 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1
transform 1 0 82156 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1
transform 1 0 82340 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _120_
timestamp 1
transform 1 0 84272 0 -1 76160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _121_
timestamp 1
transform 1 0 86204 0 1 76160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _122_
timestamp 1
transform 1 0 86664 0 -1 76160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _123_
timestamp 1
transform 1 0 86848 0 -1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _124_
timestamp 1
transform 1 0 88780 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _125_
timestamp 1
transform 1 0 89424 0 -1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _126_
timestamp 1
transform 1 0 91356 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _127_
timestamp 1
transform 1 0 93932 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _128_
timestamp 1
transform -1 0 83444 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _129_
timestamp 1
transform -1 0 86020 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _130_
timestamp 1
transform 1 0 88688 0 1 70720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _131_
timestamp 1
transform 1 0 89976 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _132_
timestamp 1
transform -1 0 89240 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _133_
timestamp 1
transform -1 0 88504 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _134_
timestamp 1
transform -1 0 88044 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _135_
timestamp 1
transform 1 0 83996 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _136_
timestamp 1
transform -1 0 75440 0 -1 72896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _137_
timestamp 1
transform -1 0 21620 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _138_
timestamp 1
transform 1 0 21712 0 1 76160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _139_
timestamp 1
transform 1 0 22448 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _140_
timestamp 1
transform -1 0 24656 0 -1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _141_
timestamp 1
transform -1 0 26496 0 -1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _142_
timestamp 1
transform -1 0 26864 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _143_
timestamp 1
transform 1 0 82432 0 1 75072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _144_
timestamp 1
transform 1 0 82984 0 1 76160
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform -1 0 22816 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1
transform 1 0 83904 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A0
timestamp 1
transform -1 0 31740 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A1
timestamp 1
transform 1 0 31740 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__S
timestamp 1
transform 1 0 32108 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A0
timestamp 1
transform -1 0 33672 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A1
timestamp 1
transform 1 0 33672 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__S
timestamp 1
transform 1 0 34132 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A0
timestamp 1
transform -1 0 35880 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A1
timestamp 1
transform 1 0 35880 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__S
timestamp 1
transform 1 0 36064 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A0
timestamp 1
transform -1 0 38272 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A1
timestamp 1
transform 1 0 38272 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__S
timestamp 1
transform 1 0 38456 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A0
timestamp 1
transform -1 0 40848 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A1
timestamp 1
transform 1 0 40848 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__S
timestamp 1
transform 1 0 41032 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A0
timestamp 1
transform -1 0 43424 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A1
timestamp 1
transform 1 0 43424 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__S
timestamp 1
transform 1 0 43608 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A0
timestamp 1
transform -1 0 60812 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A1
timestamp 1
transform 1 0 60444 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__S
timestamp 1
transform 1 0 61824 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__X
timestamp 1
transform -1 0 61824 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A0
timestamp 1
transform -1 0 62652 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A1
timestamp 1
transform 1 0 62652 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__S
timestamp 1
transform 1 0 64032 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__X
timestamp 1
transform -1 0 64032 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A0
timestamp 1
transform -1 0 65228 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A1
timestamp 1
transform 1 0 65228 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__S
timestamp 1
transform 1 0 66608 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__X
timestamp 1
transform -1 0 66608 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A0
timestamp 1
transform -1 0 67804 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A1
timestamp 1
transform 1 0 67804 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__S
timestamp 1
transform -1 0 69368 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__X
timestamp 1
transform -1 0 69184 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A0
timestamp 1
transform 1 0 69368 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A1
timestamp 1
transform 1 0 69184 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__S
timestamp 1
transform 1 0 70472 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__X
timestamp 1
transform -1 0 70472 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A0
timestamp 1
transform -1 0 71208 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A1
timestamp 1
transform 1 0 70840 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__S
timestamp 1
transform 1 0 72036 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A0
timestamp 1
transform -1 0 73692 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A1
timestamp 1
transform 1 0 73324 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__S
timestamp 1
transform 1 0 75072 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A0
timestamp 1
transform 1 0 75716 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A1
timestamp 1
transform -1 0 75716 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__S
timestamp 1
transform 1 0 75624 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A0
timestamp 1
transform -1 0 77924 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A1
timestamp 1
transform 1 0 78108 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__S
timestamp 1
transform 1 0 77924 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A0
timestamp 1
transform -1 0 80132 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A1
timestamp 1
transform 1 0 79764 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__S
timestamp 1
transform 1 0 79580 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1
transform -1 0 78200 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1
transform 1 0 89056 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1
transform 1 0 89976 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1
transform 1 0 91448 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1
transform 1 0 81696 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1
transform 1 0 82984 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1
transform 1 0 74336 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1
transform 1 0 27784 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1
transform 1 0 29164 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1
transform 1 0 30452 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1
transform 1 0 31188 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1
transform 1 0 31740 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1
transform 1 0 32476 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1
transform 1 0 82432 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1
transform 1 0 82156 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__CLK
timestamp 1
transform 1 0 86664 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__D
timestamp 1
transform 1 0 84088 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__Q
timestamp 1
transform 1 0 86480 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__CLK
timestamp 1
transform 1 0 88872 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__D
timestamp 1
transform -1 0 86112 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__Q
timestamp 1
transform -1 0 88872 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__CLK
timestamp 1
transform 1 0 88780 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__D
timestamp 1
transform -1 0 87032 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__Q
timestamp 1
transform 1 0 88504 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__CLK
timestamp 1
transform 1 0 88964 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__Q
timestamp 1
transform -1 0 88964 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__CLK
timestamp 1
transform 1 0 90804 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__Q
timestamp 1
transform 1 0 90620 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__CLK
timestamp 1
transform 1 0 91908 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__Q
timestamp 1
transform -1 0 91448 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__CLK
timestamp 1
transform 1 0 93196 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__CLK
timestamp 1
transform -1 0 95956 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__CLK
timestamp 1
transform 1 0 83628 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__CLK
timestamp 1
transform 1 0 86664 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__CLK
timestamp 1
transform 1 0 90528 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__CLK
timestamp 1
transform 1 0 91816 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__CLK
timestamp 1
transform 1 0 88780 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__CLK
timestamp 1
transform 1 0 88504 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__CLK
timestamp 1
transform 1 0 87216 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__CLK
timestamp 1
transform 1 0 83812 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__CLK
timestamp 1
transform 1 0 73416 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__CLK
timestamp 1
transform 1 0 19596 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__Q
timestamp 1
transform -1 0 21988 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__CLK
timestamp 1
transform 1 0 21528 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__Q
timestamp 1
transform -1 0 23736 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__CLK
timestamp 1
transform 1 0 22264 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__Q
timestamp 1
transform -1 0 24564 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__CLK
timestamp 1
transform 1 0 24840 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__Q
timestamp 1
transform -1 0 24840 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__CLK
timestamp 1
transform 1 0 26680 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__Q
timestamp 1
transform -1 0 26680 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__CLK
timestamp 1
transform -1 0 27232 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__Q
timestamp 1
transform -1 0 27600 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__CLK
timestamp 1
transform 1 0 81972 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__D
timestamp 1
transform -1 0 81972 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__Q
timestamp 1
transform -1 0 84456 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__CLK
timestamp 1
transform 1 0 85008 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__D
timestamp 1
transform -1 0 82984 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__Q
timestamp 1
transform -1 0 85008 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1
transform -1 0 56028 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 1
transform 1 0 57868 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_A
timestamp 1
transform -1 0 104512 0 1 90304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_X
timestamp 1
transform -1 0 106352 0 -1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_A
timestamp 1
transform 1 0 94208 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_X
timestamp 1
transform -1 0 96692 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_A
timestamp 1
transform 1 0 7268 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_X
timestamp 1
transform 1 0 7452 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_A
timestamp 1
transform 1 0 46460 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_X
timestamp 1
transform 1 0 46644 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload0_A
timestamp 1
transform 1 0 6900 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload1_A
timestamp 1
transform 1 0 44620 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout83_A
timestamp 1
transform 1 0 75440 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout83_X
timestamp 1
transform 1 0 75256 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout84_X
timestamp 1
transform -1 0 78292 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout111_A
timestamp 1
transform 1 0 89056 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout112_A
timestamp 1
transform 1 0 90160 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout112_X
timestamp 1
transform 1 0 90712 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_A
timestamp 1
transform -1 0 90528 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_X
timestamp 1
transform -1 0 90712 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1
transform -1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_X
timestamp 1
transform -1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1
transform -1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_X
timestamp 1
transform 1 0 2300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1
transform -1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_X
timestamp 1
transform -1 0 1932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1
transform -1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_X
timestamp 1
transform -1 0 1932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1
transform -1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_X
timestamp 1
transform -1 0 1932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1
transform -1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_X
timestamp 1
transform 1 0 1748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1
transform -1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_X
timestamp 1
transform 1 0 1748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1
transform -1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_X
timestamp 1
transform -1 0 1932 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1
transform -1 0 2116 0 -1 89216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_X
timestamp 1
transform 1 0 1748 0 -1 89216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1
transform -1 0 1564 0 -1 80512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_X
timestamp 1
transform -1 0 2484 0 1 80512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1
transform -1 0 1840 0 -1 104448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1
transform -1 0 1840 0 1 105536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1
transform -1 0 1840 0 1 106624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1
transform -1 0 1840 0 -1 108800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1
transform -1 0 1840 0 -1 109888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1
transform -1 0 1840 0 1 110976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1
transform -1 0 2024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_X
timestamp 1
transform 1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1
transform -1 0 1840 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1
transform -1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_X
timestamp 1
transform -1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1
transform -1 0 37444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1
transform -1 0 38732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1
transform -1 0 40020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1
transform -1 0 41308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1
transform -1 0 41952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1
transform -1 0 43240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1
transform -1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_X
timestamp 1
transform 1 0 1748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1
transform -1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_X
timestamp 1
transform -1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1
transform -1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_X
timestamp 1
transform -1 0 1932 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1
transform -1 0 2300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_X
timestamp 1
transform 1 0 1748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1
transform -1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1
transform -1 0 32936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1
transform -1 0 34224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1
transform -1 0 35512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1
transform -1 0 36156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1
transform -1 0 2116 0 -1 81600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_X
timestamp 1
transform 1 0 1748 0 -1 81600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1
transform -1 0 2116 0 1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_X
timestamp 1
transform 1 0 1748 0 1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1
transform -1 0 2116 0 1 81600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_X
timestamp 1
transform -1 0 1932 0 1 81600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1
transform -1 0 2116 0 -1 82688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_X
timestamp 1
transform 1 0 1748 0 -1 82688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1
transform -1 0 2116 0 -1 83776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_X
timestamp 1
transform 1 0 1748 0 -1 83776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1
transform -1 0 2116 0 -1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_X
timestamp 1
transform 1 0 1748 0 -1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1
transform -1 0 2116 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_X
timestamp 1
transform -1 0 1932 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1
transform -1 0 2116 0 -1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_X
timestamp 1
transform 1 0 1748 0 -1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1
transform -1 0 2116 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_X
timestamp 1
transform -1 0 1932 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1
transform -1 0 2116 0 1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_X
timestamp 1
transform 1 0 1748 0 1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1
transform -1 0 2116 0 -1 87040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_X
timestamp 1
transform 1 0 1748 0 -1 87040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1
transform -1 0 2116 0 1 83776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_X
timestamp 1
transform -1 0 1932 0 1 83776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1
transform -1 0 2116 0 1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_X
timestamp 1
transform -1 0 1932 0 1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1
transform -1 0 2116 0 -1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_X
timestamp 1
transform 1 0 1748 0 -1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1
transform -1 0 2116 0 1 87040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_X
timestamp 1
transform -1 0 1932 0 1 87040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1
transform -1 0 2116 0 -1 88128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_X
timestamp 1
transform 1 0 1748 0 -1 88128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1
transform -1 0 108284 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_X
timestamp 1
transform 1 0 107916 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew85_X
timestamp 1
transform -1 0 92368 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew87_X
timestamp 1
transform -1 0 92000 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew91_X
timestamp 1
transform -1 0 90344 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew94_X
timestamp 1
transform -1 0 91816 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew97_X
timestamp 1
transform 1 0 89976 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew98_X
timestamp 1
transform 1 0 92736 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew99_X
timestamp 1
transform -1 0 92920 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew100_X
timestamp 1
transform -1 0 91264 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew101_X
timestamp 1
transform 1 0 92184 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew104_X
timestamp 1
transform -1 0 87400 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew106_X
timestamp 1
transform -1 0 85928 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[0]
timestamp 1
transform -1 0 23644 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[1]
timestamp 1
transform -1 0 24840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[2]
timestamp 1
transform -1 0 7636 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[3]
timestamp 1
transform -1 0 7636 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[4]
timestamp 1
transform -1 0 7636 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[5]
timestamp 1
transform -1 0 7636 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[6]
timestamp 1
transform -1 0 7636 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[7]
timestamp 1
transform -1 0 7636 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[2]
timestamp 1
transform -1 0 104512 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[3]
timestamp 1
transform -1 0 104512 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[4]
timestamp 1
transform -1 0 104512 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[5]
timestamp 1
transform -1 0 90712 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[6]
timestamp 1
transform -1 0 90896 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[7]
timestamp 1
transform -1 0 91080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_clk0
timestamp 1
transform -1 0 16284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_clk1
timestamp 1
transform 1 0 96232 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_csb0
timestamp 1
transform -1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_din0[0]
timestamp 1
transform -1 0 26036 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_din0[1]
timestamp 1
transform -1 0 27140 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_din0[2]
timestamp 1
transform -1 0 28336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_din0[3]
timestamp 1
transform -1 0 29716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_din0[4]
timestamp 1
transform -1 0 30636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[0]
timestamp 1
transform -1 0 36248 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[1]
timestamp 1
transform -1 0 38824 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[2]
timestamp 1
transform -1 0 41308 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[3]
timestamp 1
transform -1 0 43792 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[4]
timestamp 1
transform -1 0 46276 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[5]
timestamp 1
transform -1 0 48760 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[6]
timestamp 1
transform 1 0 51060 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[7]
timestamp 1
transform 1 0 53544 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[8]
timestamp 1
transform 1 0 56120 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[9]
timestamp 1
transform 1 0 58604 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[10]
timestamp 1
transform 1 0 61088 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[11]
timestamp 1
transform 1 0 63572 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[12]
timestamp 1
transform 1 0 66056 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[13]
timestamp 1
transform 1 0 68540 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[14]
timestamp 1
transform 1 0 71024 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[15]
timestamp 1
transform 1 0 73508 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr0[0]
timestamp 1
transform -1 0 25024 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr0[1]
timestamp 1
transform -1 0 24840 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[0]
timestamp 1
transform -1 0 87492 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[1]
timestamp 1
transform -1 0 86388 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[2]
timestamp 1
transform -1 0 104512 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[3]
timestamp 1
transform -1 0 104512 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[4]
timestamp 1
transform -1 0 104512 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_clk0
timestamp 1
transform 1 0 16100 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_clk1
timestamp 1
transform -1 0 96048 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[0]
timestamp 1
transform -1 0 27784 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[1]
timestamp 1
transform -1 0 27416 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[2]
timestamp 1
transform -1 0 28336 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[3]
timestamp 1
transform -1 0 29716 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[4]
timestamp 1
transform -1 0 30636 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[5]
timestamp 1
transform -1 0 32476 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[6]
timestamp 1
transform -1 0 32660 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[7]
timestamp 1
transform -1 0 34132 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[8]
timestamp 1
transform -1 0 34868 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[9]
timestamp 1
transform -1 0 36524 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[10]
timestamp 1
transform -1 0 37168 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[11]
timestamp 1
transform -1 0 38824 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[12]
timestamp 1
transform -1 0 39744 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[13]
timestamp 1
transform -1 0 41400 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[14]
timestamp 1
transform -1 0 42320 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[15]
timestamp 1
transform -1 0 43976 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_dout1[0]
timestamp 1
transform -1 0 36248 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output52_A
timestamp 1
transform 1 0 1656 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output53_A
timestamp 1
transform 1 0 108100 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1
transform 1 0 108100 0 -1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output55_A
timestamp 1
transform -1 0 108284 0 1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1
transform 1 0 108100 0 -1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output59_A
timestamp 1
transform 1 0 1656 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output60_A
timestamp 1
transform -1 0 1840 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output61_A
timestamp 1
transform 1 0 1656 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output62_A
timestamp 1
transform 1 0 1656 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output63_A
timestamp 1
transform -1 0 1840 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1
transform -1 0 108284 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output65_A
timestamp 1
transform 1 0 108100 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 1
transform 1 0 108100 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output67_A
timestamp 1
transform -1 0 108284 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire68_X
timestamp 1
transform -1 0 61088 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire69_X
timestamp 1
transform -1 0 58604 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire70_X
timestamp 1
transform -1 0 56212 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire71_X
timestamp 1
transform -1 0 54004 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire72_X
timestamp 1
transform -1 0 48116 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire73_X
timestamp 1
transform -1 0 45632 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire74_X
timestamp 1
transform -1 0 43332 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire75_X
timestamp 1
transform -1 0 41032 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire76_X
timestamp 1
transform -1 0 38548 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire77_X
timestamp 1
transform -1 0 74612 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire78_X
timestamp 1
transform -1 0 72588 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire79_X
timestamp 1
transform -1 0 70196 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire80_X
timestamp 1
transform -1 0 67988 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire81_X
timestamp 1
transform -1 0 65412 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire82_X
timestamp 1
transform -1 0 63572 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform 1 0 56028 0 1 71808
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1
transform 1 0 104328 0 -1 91392
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1
transform 1 0 94392 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1
transform -1 0 7636 0 1 59840
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1
transform 1 0 44620 0 -1 72896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 1
transform 1 0 7084 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  clkload1
timestamp 1
transform 1 0 43976 0 -1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 1
transform 1 0 74520 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout84
timestamp 1
transform 1 0 77556 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout111
timestamp 1
transform -1 0 89056 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout112
timestamp 1
transform -1 0 90160 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout113
timestamp 1
transform -1 0 89608 0 1 68544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636968456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636968456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636968456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636968456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636968456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_321
timestamp 1
transform 1 0 30636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_329
timestamp 1
transform 1 0 31372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_343
timestamp 1
transform 1 0 32660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_349
timestamp 1
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_357
timestamp 1
transform 1 0 33948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_365
timestamp 1
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_371
timestamp 1
transform 1 0 35236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_377
timestamp 1
transform 1 0 35788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_398
timestamp 1
transform 1 0 37720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_406
timestamp 1
transform 1 0 38456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_426
timestamp 1
transform 1 0 40296 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_434
timestamp 1
transform 1 0 41032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_440
timestamp 1
transform 1 0 41584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_449
timestamp 1
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_455
timestamp 1
transform 1 0 42964 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1636968456
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1636968456
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1636968456
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1636968456
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1636968456
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1636968456
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1636968456
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1636968456
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1636968456
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1636968456
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1636968456
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_617
timestamp 1636968456
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_629
timestamp 1636968456
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1636968456
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1636968456
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1636968456
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_685
timestamp 1636968456
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1636968456
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1636968456
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1636968456
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1636968456
transform 1 0 69276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1636968456
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1636968456
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1636968456
transform 1 0 73324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_797
timestamp 1636968456
transform 1 0 74428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 1
transform 1 0 75532 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1636968456
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1636968456
transform 1 0 77004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1
transform 1 0 78108 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1636968456
transform 1 0 78476 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1636968456
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1636968456
transform 1 0 81052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1636968456
transform 1 0 82156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 1
transform 1 0 83260 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1636968456
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1636968456
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1636968456
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1636968456
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1636968456
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1636968456
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1636968456
transform 1 0 91356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1636968456
transform 1 0 92460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1009
timestamp 1636968456
transform 1 0 93932 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1021
timestamp 1636968456
transform 1 0 95036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1037
timestamp 1636968456
transform 1 0 96508 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1049
timestamp 1636968456
transform 1 0 97612 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1061
timestamp 1
transform 1 0 98716 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1636968456
transform 1 0 99084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1636968456
transform 1 0 100188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1636968456
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1105
timestamp 1636968456
transform 1 0 102764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1121
timestamp 1636968456
transform 1 0 104236 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1133
timestamp 1636968456
transform 1 0 105340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1149
timestamp 1636968456
transform 1 0 106812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1161
timestamp 1
transform 1 0 107916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1167
timestamp 1
transform 1 0 108468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636968456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636968456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636968456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636968456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636968456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636968456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636968456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636968456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636968456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636968456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636968456
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636968456
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636968456
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636968456
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636968456
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636968456
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636968456
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636968456
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636968456
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636968456
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636968456
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636968456
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636968456
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636968456
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1636968456
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1636968456
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1636968456
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1636968456
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1636968456
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1636968456
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1636968456
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1636968456
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1636968456
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1636968456
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1636968456
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1636968456
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1636968456
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1636968456
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1636968456
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1636968456
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 1
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1636968456
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1636968456
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1636968456
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1636968456
transform 1 0 81788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 1
transform 1 0 82892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1636968456
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1636968456
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1636968456
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1636968456
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1636968456
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1636968456
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1636968456
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1636968456
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1636968456
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1636968456
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1636968456
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1045
timestamp 1636968456
transform 1 0 97244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1057
timestamp 1
transform 1 0 98348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1636968456
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1636968456
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1636968456
transform 1 0 101292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1636968456
transform 1 0 102396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1
transform 1 0 103500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1636968456
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1636968456
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1636968456
transform 1 0 106444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1157
timestamp 1
transform 1 0 107548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1165
timestamp 1
transform 1 0 108284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636968456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636968456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636968456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636968456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636968456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636968456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636968456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636968456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636968456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636968456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636968456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636968456
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636968456
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636968456
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636968456
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636968456
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636968456
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636968456
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636968456
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636968456
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636968456
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636968456
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636968456
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636968456
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1636968456
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1636968456
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1636968456
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1636968456
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1636968456
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1636968456
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1636968456
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1636968456
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1636968456
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1636968456
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1636968456
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1636968456
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1636968456
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1636968456
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1636968456
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1636968456
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1636968456
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1636968456
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1636968456
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1636968456
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1636968456
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1636968456
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1636968456
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1636968456
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1636968456
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1636968456
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1636968456
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1636968456
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1636968456
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1636968456
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1636968456
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1636968456
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1636968456
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1636968456
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1636968456
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1636968456
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1636968456
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1636968456
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1636968456
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1161
timestamp 1
transform 1 0 107916 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1167
timestamp 1
transform 1 0 108468 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636968456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636968456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636968456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636968456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636968456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636968456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636968456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636968456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636968456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636968456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636968456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636968456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636968456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636968456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636968456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636968456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636968456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636968456
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636968456
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636968456
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636968456
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636968456
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636968456
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636968456
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636968456
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636968456
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636968456
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636968456
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636968456
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636968456
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636968456
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636968456
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636968456
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636968456
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1636968456
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1636968456
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1636968456
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636968456
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636968456
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1636968456
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1636968456
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1636968456
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1636968456
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1636968456
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1636968456
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1636968456
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1636968456
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1636968456
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1636968456
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1636968456
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1636968456
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1636968456
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1636968456
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1636968456
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1636968456
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1636968456
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1636968456
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1636968456
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1636968456
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1636968456
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1636968456
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1636968456
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1636968456
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1636968456
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1636968456
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1636968456
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1636968456
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1636968456
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1157
timestamp 1
transform 1 0 107548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1165
timestamp 1
transform 1 0 108284 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636968456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636968456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636968456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636968456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636968456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636968456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636968456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636968456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636968456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636968456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636968456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636968456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636968456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636968456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636968456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636968456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636968456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636968456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636968456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636968456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1636968456
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1636968456
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636968456
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636968456
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1636968456
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1636968456
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636968456
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636968456
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1636968456
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1636968456
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636968456
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636968456
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1636968456
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1636968456
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636968456
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636968456
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1636968456
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1636968456
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636968456
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636968456
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1636968456
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1636968456
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636968456
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636968456
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1636968456
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1636968456
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1636968456
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1636968456
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1636968456
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1636968456
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1636968456
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1636968456
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1636968456
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1636968456
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1636968456
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1636968456
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1636968456
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1636968456
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1636968456
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1636968456
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1636968456
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1636968456
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1636968456
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1636968456
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1636968456
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1636968456
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1636968456
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1636968456
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1636968456
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1636968456
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1636968456
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1161
timestamp 1
transform 1 0 107916 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1167
timestamp 1
transform 1 0 108468 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_11
timestamp 1636968456
transform 1 0 2116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_23
timestamp 1636968456
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1636968456
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636968456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636968456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636968456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636968456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636968456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636968456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636968456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636968456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636968456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636968456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636968456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636968456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636968456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636968456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636968456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636968456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636968456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636968456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636968456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636968456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636968456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636968456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636968456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636968456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1636968456
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1636968456
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1636968456
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1636968456
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1636968456
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1636968456
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1636968456
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1636968456
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1636968456
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1636968456
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1636968456
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1636968456
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1636968456
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1636968456
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1636968456
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1636968456
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1636968456
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1636968456
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1636968456
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1636968456
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1636968456
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1636968456
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1636968456
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1636968456
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1636968456
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1636968456
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1636968456
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1636968456
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1636968456
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1636968456
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1636968456
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1636968456
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1636968456
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1636968456
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1636968456
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1636968456
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1636968456
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1636968456
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1636968456
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1636968456
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1636968456
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1636968456
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1636968456
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1636968456
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1636968456
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1636968456
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1636968456
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1636968456
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1636968456
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1636968456
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1636968456
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1157
timestamp 1
transform 1 0 107548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1165
timestamp 1
transform 1 0 108284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_10
timestamp 1636968456
transform 1 0 2024 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 1
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636968456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636968456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636968456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636968456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636968456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636968456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636968456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636968456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636968456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636968456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636968456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636968456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636968456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636968456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636968456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636968456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636968456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636968456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636968456
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636968456
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636968456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636968456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636968456
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1636968456
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636968456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636968456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1636968456
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1636968456
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1636968456
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1636968456
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1636968456
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1636968456
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1636968456
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1636968456
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1636968456
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1636968456
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1636968456
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1636968456
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1636968456
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1636968456
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1636968456
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1636968456
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1636968456
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1636968456
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1636968456
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1636968456
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1636968456
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1636968456
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1636968456
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1636968456
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1636968456
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1636968456
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1636968456
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1636968456
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1636968456
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1636968456
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1636968456
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1636968456
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1636968456
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1636968456
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1636968456
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1636968456
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1636968456
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1636968456
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1636968456
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1636968456
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1636968456
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1636968456
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1636968456
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1636968456
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1636968456
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1636968456
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1636968456
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1636968456
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1636968456
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1636968456
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1636968456
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1161
timestamp 1
transform 1 0 107916 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1167
timestamp 1
transform 1 0 108468 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_11
timestamp 1636968456
transform 1 0 2116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_23
timestamp 1636968456
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1636968456
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636968456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636968456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636968456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636968456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636968456
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636968456
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636968456
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636968456
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636968456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636968456
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636968456
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636968456
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636968456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636968456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636968456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636968456
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636968456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636968456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636968456
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636968456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636968456
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636968456
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636968456
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636968456
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636968456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636968456
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1636968456
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1636968456
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1636968456
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1636968456
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1636968456
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1636968456
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1636968456
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1636968456
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1636968456
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1636968456
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1636968456
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1636968456
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1636968456
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1636968456
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1636968456
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1636968456
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1636968456
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1636968456
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1636968456
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1636968456
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1636968456
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1636968456
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1636968456
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1636968456
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1636968456
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1636968456
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1636968456
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1636968456
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1636968456
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1636968456
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1636968456
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1636968456
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1636968456
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1636968456
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1636968456
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1636968456
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1636968456
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1636968456
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1636968456
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1636968456
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1636968456
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1636968456
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1636968456
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1636968456
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1636968456
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1636968456
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1636968456
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1636968456
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1636968456
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1636968456
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1636968456
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1636968456
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1636968456
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1157
timestamp 1
transform 1 0 107548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1165
timestamp 1
transform 1 0 108284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636968456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636968456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636968456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636968456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636968456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636968456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636968456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636968456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636968456
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636968456
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636968456
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636968456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636968456
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636968456
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636968456
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636968456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636968456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636968456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636968456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636968456
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636968456
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636968456
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636968456
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636968456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636968456
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1636968456
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1636968456
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636968456
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636968456
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1636968456
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1636968456
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1636968456
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1636968456
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1636968456
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1636968456
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1636968456
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1636968456
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1636968456
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1636968456
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1636968456
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1636968456
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1636968456
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1636968456
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1636968456
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1636968456
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1636968456
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1636968456
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1636968456
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1636968456
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1636968456
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1636968456
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1636968456
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1636968456
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1636968456
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1636968456
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1636968456
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1636968456
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1636968456
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1636968456
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1636968456
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1636968456
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1636968456
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1636968456
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1636968456
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1636968456
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1636968456
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1636968456
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1636968456
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1636968456
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1636968456
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1636968456
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1636968456
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1636968456
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1636968456
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1636968456
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1636968456
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1636968456
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1636968456
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1636968456
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1636968456
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1161
timestamp 1
transform 1 0 107916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1167
timestamp 1
transform 1 0 108468 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_11
timestamp 1636968456
transform 1 0 2116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_29
timestamp 1636968456
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_41
timestamp 1636968456
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636968456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636968456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp 1
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_85
timestamp 1636968456
transform 1 0 8924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_97
timestamp 1636968456
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636968456
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636968456
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp 1
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_141
timestamp 1636968456
transform 1 0 14076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_153
timestamp 1
transform 1 0 15180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636968456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636968456
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1636968456
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_209
timestamp 1636968456
transform 1 0 20332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636968456
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_237
timestamp 1
transform 1 0 22908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_245
timestamp 1
transform 1 0 23644 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_251
timestamp 1
transform 1 0 24196 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_253
timestamp 1
transform 1 0 24380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_258
timestamp 1
transform 1 0 24840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_266
timestamp 1
transform 1 0 25576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_271
timestamp 1
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_283
timestamp 1
transform 1 0 27140 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_291
timestamp 1
transform 1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_296
timestamp 1636968456
transform 1 0 28336 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_311
timestamp 1
transform 1 0 29716 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_321
timestamp 1636968456
transform 1 0 30636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636968456
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1636968456
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp 1
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_365
timestamp 1636968456
transform 1 0 34684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_377
timestamp 1636968456
transform 1 0 35788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636968456
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1636968456
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_417
timestamp 1
transform 1 0 39468 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_421
timestamp 1636968456
transform 1 0 39836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_433
timestamp 1636968456
transform 1 0 40940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1636968456
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1636968456
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_473
timestamp 1
transform 1 0 44620 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_477
timestamp 1636968456
transform 1 0 44988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_489
timestamp 1636968456
transform 1 0 46092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1636968456
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1636968456
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_529
timestamp 1
transform 1 0 49772 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_533
timestamp 1636968456
transform 1 0 50140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_545
timestamp 1636968456
transform 1 0 51244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_557
timestamp 1
transform 1 0 52348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1636968456
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1636968456
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_585
timestamp 1
transform 1 0 54924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_589
timestamp 1636968456
transform 1 0 55292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_601
timestamp 1636968456
transform 1 0 56396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_613
timestamp 1
transform 1 0 57500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1636968456
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1636968456
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_641
timestamp 1
transform 1 0 60076 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_645
timestamp 1636968456
transform 1 0 60444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_657
timestamp 1636968456
transform 1 0 61548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_669
timestamp 1
transform 1 0 62652 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1636968456
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1636968456
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_697
timestamp 1
transform 1 0 65228 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_701
timestamp 1636968456
transform 1 0 65596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_713
timestamp 1636968456
transform 1 0 66700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_725
timestamp 1
transform 1 0 67804 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1636968456
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1636968456
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_753
timestamp 1
transform 1 0 70380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_757
timestamp 1636968456
transform 1 0 70748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_769
timestamp 1636968456
transform 1 0 71852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_781
timestamp 1
transform 1 0 72956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1636968456
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1636968456
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_809
timestamp 1
transform 1 0 75532 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_813
timestamp 1636968456
transform 1 0 75900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_825
timestamp 1636968456
transform 1 0 77004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_837
timestamp 1
transform 1 0 78108 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1636968456
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1636968456
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_865
timestamp 1
transform 1 0 80684 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_869
timestamp 1636968456
transform 1 0 81052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_881
timestamp 1636968456
transform 1 0 82156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_893
timestamp 1
transform 1 0 83260 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1636968456
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1636968456
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_921
timestamp 1
transform 1 0 85836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_925
timestamp 1636968456
transform 1 0 86204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_937
timestamp 1636968456
transform 1 0 87308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_949
timestamp 1
transform 1 0 88412 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1636968456
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_965
timestamp 1
transform 1 0 89884 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_971
timestamp 1
transform 1 0 90436 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_978
timestamp 1
transform 1 0 91080 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_981
timestamp 1636968456
transform 1 0 91356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_993
timestamp 1636968456
transform 1 0 92460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1005
timestamp 1
transform 1 0 93564 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1636968456
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1636968456
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1033
timestamp 1
transform 1 0 96140 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1037
timestamp 1636968456
transform 1 0 96508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1049
timestamp 1636968456
transform 1 0 97612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1061
timestamp 1
transform 1 0 98716 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1636968456
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1636968456
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1089
timestamp 1
transform 1 0 101292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1093
timestamp 1636968456
transform 1 0 101660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1105
timestamp 1636968456
transform 1 0 102764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1117
timestamp 1
transform 1 0 103868 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1636968456
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1636968456
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1145
timestamp 1
transform 1 0 106444 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1149
timestamp 1636968456
transform 1 0 106812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1161
timestamp 1
transform 1 0 107916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1167
timestamp 1
transform 1 0 108468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_13
timestamp 1636968456
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636968456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636968456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636968456
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 1
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1122
timestamp 1636968456
transform 1 0 104328 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1134
timestamp 1636968456
transform 1 0 105432 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1146
timestamp 1
transform 1 0 106536 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1148
timestamp 1636968456
transform 1 0 106720 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1160
timestamp 1
transform 1 0 107824 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636968456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636968456
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636968456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1122
timestamp 1636968456
transform 1 0 104328 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1134
timestamp 1636968456
transform 1 0 105432 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1146
timestamp 1636968456
transform 1 0 106536 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1158
timestamp 1
transform 1 0 107640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1166
timestamp 1
transform 1 0 108376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_11
timestamp 1636968456
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636968456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636968456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636968456
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_65
timestamp 1
transform 1 0 7084 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1122
timestamp 1636968456
transform 1 0 104328 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1134
timestamp 1636968456
transform 1 0 105432 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1146
timestamp 1
transform 1 0 106536 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1148
timestamp 1636968456
transform 1 0 106720 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1160
timestamp 1
transform 1 0 107824 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636968456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636968456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636968456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636968456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_69
timestamp 1
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1122
timestamp 1636968456
transform 1 0 104328 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1134
timestamp 1636968456
transform 1 0 105432 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1146
timestamp 1636968456
transform 1 0 106536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1158
timestamp 1
transform 1 0 107640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1166
timestamp 1
transform 1 0 108376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_11
timestamp 1636968456
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636968456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636968456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636968456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1
transform 1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1122
timestamp 1636968456
transform 1 0 104328 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1134
timestamp 1636968456
transform 1 0 105432 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1146
timestamp 1
transform 1 0 106536 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1148
timestamp 1636968456
transform 1 0 106720 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1160
timestamp 1
transform 1 0 107824 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_11
timestamp 1636968456
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1636968456
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1636968456
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636968456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1122
timestamp 1636968456
transform 1 0 104328 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1134
timestamp 1636968456
transform 1 0 105432 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1146
timestamp 1636968456
transform 1 0 106536 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1158
timestamp 1
transform 1 0 107640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1166
timestamp 1
transform 1 0 108376 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_11
timestamp 1636968456
transform 1 0 2116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636968456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636968456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636968456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_65
timestamp 1
transform 1 0 7084 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1122
timestamp 1636968456
transform 1 0 104328 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1134
timestamp 1636968456
transform 1 0 105432 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1146
timestamp 1
transform 1 0 106536 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1148
timestamp 1636968456
transform 1 0 106720 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1160
timestamp 1
transform 1 0 107824 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1636968456
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1636968456
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1636968456
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636968456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1122
timestamp 1636968456
transform 1 0 104328 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1134
timestamp 1636968456
transform 1 0 105432 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1146
timestamp 1636968456
transform 1 0 106536 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1158
timestamp 1
transform 1 0 107640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1166
timestamp 1
transform 1 0 108376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636968456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636968456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636968456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636968456
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636968456
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_65
timestamp 1
transform 1 0 7084 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1122
timestamp 1636968456
transform 1 0 104328 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1134
timestamp 1636968456
transform 1 0 105432 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1146
timestamp 1
transform 1 0 106536 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1148
timestamp 1636968456
transform 1 0 106720 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1160
timestamp 1
transform 1 0 107824 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_11
timestamp 1636968456
transform 1 0 2116 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_23
timestamp 1636968456
transform 1 0 3220 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_35
timestamp 1636968456
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636968456
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1122
timestamp 1636968456
transform 1 0 104328 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1134
timestamp 1636968456
transform 1 0 105432 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1146
timestamp 1636968456
transform 1 0 106536 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1158
timestamp 1
transform 1 0 107640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1166
timestamp 1
transform 1 0 108376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_11
timestamp 1636968456
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636968456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636968456
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636968456
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_65
timestamp 1
transform 1 0 7084 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1122
timestamp 1636968456
transform 1 0 104328 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1134
timestamp 1636968456
transform 1 0 105432 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1146
timestamp 1
transform 1 0 106536 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1148
timestamp 1636968456
transform 1 0 106720 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1160
timestamp 1
transform 1 0 107824 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_11
timestamp 1636968456
transform 1 0 2116 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_23
timestamp 1636968456
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_35
timestamp 1636968456
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636968456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1122
timestamp 1636968456
transform 1 0 104328 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1134
timestamp 1636968456
transform 1 0 105432 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1146
timestamp 1636968456
transform 1 0 106536 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_1158
timestamp 1
transform 1 0 107640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_1166
timestamp 1
transform 1 0 108376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636968456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636968456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636968456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636968456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636968456
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_65
timestamp 1
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1122
timestamp 1636968456
transform 1 0 104328 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1134
timestamp 1636968456
transform 1 0 105432 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1146
timestamp 1
transform 1 0 106536 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1148
timestamp 1636968456
transform 1 0 106720 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_1160
timestamp 1
transform 1 0 107824 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636968456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636968456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636968456
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636968456
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1122
timestamp 1636968456
transform 1 0 104328 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1134
timestamp 1636968456
transform 1 0 105432 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1146
timestamp 1636968456
transform 1 0 106536 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_1158
timestamp 1
transform 1 0 107640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_1166
timestamp 1
transform 1 0 108376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636968456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636968456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636968456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636968456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636968456
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1122
timestamp 1636968456
transform 1 0 104328 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1134
timestamp 1636968456
transform 1 0 105432 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1146
timestamp 1
transform 1 0 106536 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1148
timestamp 1636968456
transform 1 0 106720 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_1160
timestamp 1
transform 1 0 107824 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636968456
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1636968456
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1636968456
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636968456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1122
timestamp 1636968456
transform 1 0 104328 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1134
timestamp 1636968456
transform 1 0 105432 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1146
timestamp 1636968456
transform 1 0 106536 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_1158
timestamp 1
transform 1 0 107640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_1166
timestamp 1
transform 1 0 108376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636968456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636968456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636968456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636968456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636968456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_65
timestamp 1
transform 1 0 7084 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1122
timestamp 1636968456
transform 1 0 104328 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1134
timestamp 1636968456
transform 1 0 105432 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1146
timestamp 1
transform 1 0 106536 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1148
timestamp 1636968456
transform 1 0 106720 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_1160
timestamp 1
transform 1 0 107824 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636968456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636968456
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636968456
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636968456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1122
timestamp 1636968456
transform 1 0 104328 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1134
timestamp 1636968456
transform 1 0 105432 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1146
timestamp 1636968456
transform 1 0 106536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_1158
timestamp 1
transform 1 0 107640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_1166
timestamp 1
transform 1 0 108376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636968456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636968456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636968456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636968456
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_65
timestamp 1
transform 1 0 7084 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1122
timestamp 1636968456
transform 1 0 104328 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1134
timestamp 1636968456
transform 1 0 105432 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1146
timestamp 1
transform 1 0 106536 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1148
timestamp 1636968456
transform 1 0 106720 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_1160
timestamp 1
transform 1 0 107824 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636968456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636968456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636968456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636968456
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636968456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1122
timestamp 1636968456
transform 1 0 104328 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1134
timestamp 1636968456
transform 1 0 105432 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1146
timestamp 1636968456
transform 1 0 106536 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_1158
timestamp 1
transform 1 0 107640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_1166
timestamp 1
transform 1 0 108376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636968456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636968456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636968456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636968456
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636968456
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_65
timestamp 1
transform 1 0 7084 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1122
timestamp 1636968456
transform 1 0 104328 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1134
timestamp 1636968456
transform 1 0 105432 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1146
timestamp 1
transform 1 0 106536 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1148
timestamp 1636968456
transform 1 0 106720 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_1160
timestamp 1
transform 1 0 107824 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636968456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636968456
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636968456
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1636968456
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636968456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_69
timestamp 1
transform 1 0 7452 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1122
timestamp 1636968456
transform 1 0 104328 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1134
timestamp 1636968456
transform 1 0 105432 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1146
timestamp 1636968456
transform 1 0 106536 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_1158
timestamp 1
transform 1 0 107640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_1166
timestamp 1
transform 1 0 108376 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636968456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636968456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636968456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636968456
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636968456
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_65
timestamp 1
transform 1 0 7084 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1122
timestamp 1636968456
transform 1 0 104328 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1134
timestamp 1636968456
transform 1 0 105432 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1146
timestamp 1
transform 1 0 106536 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1148
timestamp 1636968456
transform 1 0 106720 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_1160
timestamp 1
transform 1 0 107824 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636968456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636968456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636968456
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1636968456
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636968456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1122
timestamp 1636968456
transform 1 0 104328 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1134
timestamp 1636968456
transform 1 0 105432 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1146
timestamp 1636968456
transform 1 0 106536 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_1158
timestamp 1
transform 1 0 107640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_1166
timestamp 1
transform 1 0 108376 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636968456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636968456
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636968456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1636968456
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1636968456
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_65
timestamp 1
transform 1 0 7084 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1122
timestamp 1636968456
transform 1 0 104328 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1134
timestamp 1636968456
transform 1 0 105432 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1146
timestamp 1
transform 1 0 106536 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1148
timestamp 1636968456
transform 1 0 106720 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_1160
timestamp 1
transform 1 0 107824 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636968456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636968456
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1636968456
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1636968456
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636968456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_69
timestamp 1
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1122
timestamp 1636968456
transform 1 0 104328 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1134
timestamp 1636968456
transform 1 0 105432 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1146
timestamp 1636968456
transform 1 0 106536 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_1158
timestamp 1
transform 1 0 107640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_1166
timestamp 1
transform 1 0 108376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636968456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636968456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636968456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1636968456
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1636968456
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_65
timestamp 1
transform 1 0 7084 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1122
timestamp 1636968456
transform 1 0 104328 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1134
timestamp 1636968456
transform 1 0 105432 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1146
timestamp 1
transform 1 0 106536 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1148
timestamp 1636968456
transform 1 0 106720 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_1160
timestamp 1
transform 1 0 107824 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1636968456
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1636968456
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1636968456
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1636968456
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636968456
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_69
timestamp 1
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1124
timestamp 1636968456
transform 1 0 104512 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1136
timestamp 1636968456
transform 1 0 105616 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1148
timestamp 1636968456
transform 1 0 106720 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_1160
timestamp 1
transform 1 0 107824 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636968456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636968456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636968456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636968456
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636968456
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_65
timestamp 1
transform 1 0 7084 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1122
timestamp 1636968456
transform 1 0 104328 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1134
timestamp 1636968456
transform 1 0 105432 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1146
timestamp 1
transform 1 0 106536 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1148
timestamp 1636968456
transform 1 0 106720 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_1160
timestamp 1
transform 1 0 107824 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636968456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636968456
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636968456
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1636968456
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636968456
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_69
timestamp 1
transform 1 0 7452 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1124
timestamp 1636968456
transform 1 0 104512 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1136
timestamp 1636968456
transform 1 0 105616 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1148
timestamp 1636968456
transform 1 0 106720 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_1160
timestamp 1
transform 1 0 107824 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636968456
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636968456
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636968456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636968456
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1636968456
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_65
timestamp 1
transform 1 0 7084 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1122
timestamp 1636968456
transform 1 0 104328 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1134
timestamp 1636968456
transform 1 0 105432 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1146
timestamp 1
transform 1 0 106536 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1148
timestamp 1636968456
transform 1 0 106720 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_1160
timestamp 1
transform 1 0 107824 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636968456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636968456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1636968456
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1636968456
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636968456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1122
timestamp 1636968456
transform 1 0 104328 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1134
timestamp 1636968456
transform 1 0 105432 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1146
timestamp 1636968456
transform 1 0 106536 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_1158
timestamp 1
transform 1 0 107640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_1166
timestamp 1
transform 1 0 108376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636968456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636968456
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636968456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636968456
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636968456
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_65
timestamp 1
transform 1 0 7084 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1124
timestamp 1636968456
transform 1 0 104512 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_1136
timestamp 1
transform 1 0 105616 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_1144
timestamp 1
transform 1 0 106352 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1148
timestamp 1636968456
transform 1 0 106720 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_1160
timestamp 1
transform 1 0 107824 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636968456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636968456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636968456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636968456
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636968456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_69
timestamp 1
transform 1 0 7452 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1122
timestamp 1636968456
transform 1 0 104328 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1134
timestamp 1636968456
transform 1 0 105432 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1146
timestamp 1636968456
transform 1 0 106536 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_1158
timestamp 1
transform 1 0 107640 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_1166
timestamp 1
transform 1 0 108376 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636968456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636968456
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636968456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636968456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636968456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_65
timestamp 1
transform 1 0 7084 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1122
timestamp 1636968456
transform 1 0 104328 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1134
timestamp 1636968456
transform 1 0 105432 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1146
timestamp 1
transform 1 0 106536 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1148
timestamp 1636968456
transform 1 0 106720 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_1160
timestamp 1
transform 1 0 107824 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636968456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636968456
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636968456
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636968456
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636968456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_69
timestamp 1
transform 1 0 7452 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1122
timestamp 1636968456
transform 1 0 104328 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1134
timestamp 1636968456
transform 1 0 105432 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1146
timestamp 1636968456
transform 1 0 106536 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_1158
timestamp 1
transform 1 0 107640 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_1166
timestamp 1
transform 1 0 108376 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636968456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636968456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636968456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636968456
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1636968456
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_65
timestamp 1
transform 1 0 7084 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1122
timestamp 1636968456
transform 1 0 104328 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1134
timestamp 1636968456
transform 1 0 105432 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1146
timestamp 1
transform 1 0 106536 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1148
timestamp 1636968456
transform 1 0 106720 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1160
timestamp 1
transform 1 0 107824 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636968456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636968456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1636968456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1636968456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636968456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_69
timestamp 1
transform 1 0 7452 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1122
timestamp 1636968456
transform 1 0 104328 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1134
timestamp 1636968456
transform 1 0 105432 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1146
timestamp 1636968456
transform 1 0 106536 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_1158
timestamp 1
transform 1 0 107640 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_1166
timestamp 1
transform 1 0 108376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636968456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636968456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636968456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636968456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1636968456
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_65
timestamp 1
transform 1 0 7084 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1122
timestamp 1636968456
transform 1 0 104328 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1134
timestamp 1636968456
transform 1 0 105432 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1146
timestamp 1
transform 1 0 106536 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1148
timestamp 1636968456
transform 1 0 106720 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_1160
timestamp 1
transform 1 0 107824 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636968456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1636968456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1636968456
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1636968456
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1636968456
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_69
timestamp 1
transform 1 0 7452 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1122
timestamp 1636968456
transform 1 0 104328 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1134
timestamp 1636968456
transform 1 0 105432 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1146
timestamp 1636968456
transform 1 0 106536 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_1158
timestamp 1
transform 1 0 107640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_1166
timestamp 1
transform 1 0 108376 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1636968456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1636968456
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636968456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1636968456
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1636968456
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_65
timestamp 1
transform 1 0 7084 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1122
timestamp 1636968456
transform 1 0 104328 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1134
timestamp 1636968456
transform 1 0 105432 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1146
timestamp 1
transform 1 0 106536 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1148
timestamp 1636968456
transform 1 0 106720 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_1160
timestamp 1
transform 1 0 107824 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636968456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636968456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1636968456
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1636968456
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1636968456
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_69
timestamp 1
transform 1 0 7452 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1122
timestamp 1636968456
transform 1 0 104328 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1134
timestamp 1636968456
transform 1 0 105432 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1146
timestamp 1636968456
transform 1 0 106536 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_1158
timestamp 1
transform 1 0 107640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_1166
timestamp 1
transform 1 0 108376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636968456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636968456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636968456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1636968456
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1636968456
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_65
timestamp 1
transform 1 0 7084 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1122
timestamp 1636968456
transform 1 0 104328 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1134
timestamp 1636968456
transform 1 0 105432 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1146
timestamp 1
transform 1 0 106536 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1148
timestamp 1636968456
transform 1 0 106720 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_1160
timestamp 1
transform 1 0 107824 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636968456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636968456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636968456
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1636968456
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1636968456
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_69
timestamp 1
transform 1 0 7452 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1122
timestamp 1636968456
transform 1 0 104328 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1134
timestamp 1636968456
transform 1 0 105432 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1146
timestamp 1636968456
transform 1 0 106536 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_1158
timestamp 1
transform 1 0 107640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_1166
timestamp 1
transform 1 0 108376 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636968456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636968456
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1636968456
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1636968456
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1636968456
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_65
timestamp 1
transform 1 0 7084 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1122
timestamp 1636968456
transform 1 0 104328 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1134
timestamp 1636968456
transform 1 0 105432 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1146
timestamp 1
transform 1 0 106536 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1148
timestamp 1636968456
transform 1 0 106720 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_1160
timestamp 1
transform 1 0 107824 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1636968456
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1636968456
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1636968456
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1636968456
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1636968456
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_69
timestamp 1
transform 1 0 7452 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1122
timestamp 1636968456
transform 1 0 104328 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1134
timestamp 1636968456
transform 1 0 105432 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1146
timestamp 1636968456
transform 1 0 106536 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_1158
timestamp 1
transform 1 0 107640 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_1166
timestamp 1
transform 1 0 108376 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636968456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636968456
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636968456
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1636968456
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1636968456
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_65
timestamp 1
transform 1 0 7084 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1122
timestamp 1636968456
transform 1 0 104328 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1134
timestamp 1636968456
transform 1 0 105432 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1146
timestamp 1
transform 1 0 106536 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1148
timestamp 1636968456
transform 1 0 106720 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_1160
timestamp 1
transform 1 0 107824 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1636968456
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1636968456
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1636968456
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1636968456
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1636968456
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_69
timestamp 1
transform 1 0 7452 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1122
timestamp 1636968456
transform 1 0 104328 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1134
timestamp 1636968456
transform 1 0 105432 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1146
timestamp 1636968456
transform 1 0 106536 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_1158
timestamp 1
transform 1 0 107640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_1166
timestamp 1
transform 1 0 108376 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636968456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636968456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636968456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1636968456
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1636968456
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_65
timestamp 1
transform 1 0 7084 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1122
timestamp 1636968456
transform 1 0 104328 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1134
timestamp 1636968456
transform 1 0 105432 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1146
timestamp 1
transform 1 0 106536 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1148
timestamp 1636968456
transform 1 0 106720 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_1160
timestamp 1
transform 1 0 107824 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636968456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636968456
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1636968456
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1636968456
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1636968456
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_69
timestamp 1
transform 1 0 7452 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1122
timestamp 1636968456
transform 1 0 104328 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1134
timestamp 1636968456
transform 1 0 105432 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1146
timestamp 1636968456
transform 1 0 106536 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1158
timestamp 1
transform 1 0 107640 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_1166
timestamp 1
transform 1 0 108376 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1636968456
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1636968456
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636968456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1636968456
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1636968456
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_65
timestamp 1
transform 1 0 7084 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1122
timestamp 1636968456
transform 1 0 104328 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1134
timestamp 1636968456
transform 1 0 105432 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1146
timestamp 1
transform 1 0 106536 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1148
timestamp 1636968456
transform 1 0 106720 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_1160
timestamp 1
transform 1 0 107824 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1636968456
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1636968456
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1636968456
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1636968456
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1636968456
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1122
timestamp 1636968456
transform 1 0 104328 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1134
timestamp 1636968456
transform 1 0 105432 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1146
timestamp 1636968456
transform 1 0 106536 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1158
timestamp 1
transform 1 0 107640 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1166
timestamp 1
transform 1 0 108376 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636968456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636968456
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1636968456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1636968456
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1636968456
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_65
timestamp 1
transform 1 0 7084 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1122
timestamp 1636968456
transform 1 0 104328 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1134
timestamp 1636968456
transform 1 0 105432 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1146
timestamp 1
transform 1 0 106536 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1148
timestamp 1636968456
transform 1 0 106720 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1160
timestamp 1
transform 1 0 107824 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636968456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636968456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1636968456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1636968456
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1636968456
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1122
timestamp 1636968456
transform 1 0 104328 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1134
timestamp 1636968456
transform 1 0 105432 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1146
timestamp 1636968456
transform 1 0 106536 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1158
timestamp 1
transform 1 0 107640 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1166
timestamp 1
transform 1 0 108376 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1636968456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1636968456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1636968456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1636968456
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1636968456
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_65
timestamp 1
transform 1 0 7084 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1122
timestamp 1636968456
transform 1 0 104328 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1134
timestamp 1636968456
transform 1 0 105432 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1146
timestamp 1
transform 1 0 106536 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1148
timestamp 1636968456
transform 1 0 106720 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_1160
timestamp 1
transform 1 0 107824 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1636968456
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1636968456
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1636968456
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1636968456
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1636968456
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_69
timestamp 1
transform 1 0 7452 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1122
timestamp 1636968456
transform 1 0 104328 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1134
timestamp 1636968456
transform 1 0 105432 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1146
timestamp 1636968456
transform 1 0 106536 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_1158
timestamp 1
transform 1 0 107640 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_1166
timestamp 1
transform 1 0 108376 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1636968456
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1636968456
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1636968456
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1636968456
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1636968456
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_65
timestamp 1
transform 1 0 7084 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1122
timestamp 1636968456
transform 1 0 104328 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1134
timestamp 1636968456
transform 1 0 105432 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_1146
timestamp 1
transform 1 0 106536 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1148
timestamp 1636968456
transform 1 0 106720 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_1160
timestamp 1
transform 1 0 107824 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1636968456
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1636968456
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1636968456
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1636968456
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1636968456
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1122
timestamp 1636968456
transform 1 0 104328 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1134
timestamp 1636968456
transform 1 0 105432 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1146
timestamp 1636968456
transform 1 0 106536 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_1158
timestamp 1
transform 1 0 107640 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_1166
timestamp 1
transform 1 0 108376 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636968456
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636968456
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636968456
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1636968456
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1636968456
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_65
timestamp 1
transform 1 0 7084 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1122
timestamp 1636968456
transform 1 0 104328 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1134
timestamp 1636968456
transform 1 0 105432 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_1146
timestamp 1
transform 1 0 106536 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1148
timestamp 1636968456
transform 1 0 106720 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_1160
timestamp 1
transform 1 0 107824 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636968456
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636968456
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636968456
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1636968456
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1636968456
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1122
timestamp 1636968456
transform 1 0 104328 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1134
timestamp 1636968456
transform 1 0 105432 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1146
timestamp 1636968456
transform 1 0 106536 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_1158
timestamp 1
transform 1 0 107640 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_1166
timestamp 1
transform 1 0 108376 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1636968456
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1636968456
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636968456
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1636968456
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1636968456
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_65
timestamp 1
transform 1 0 7084 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1122
timestamp 1636968456
transform 1 0 104328 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1134
timestamp 1636968456
transform 1 0 105432 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_1146
timestamp 1
transform 1 0 106536 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1148
timestamp 1636968456
transform 1 0 106720 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_1160
timestamp 1
transform 1 0 107824 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636968456
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636968456
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1636968456
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1636968456
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1636968456
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_69
timestamp 1
transform 1 0 7452 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1122
timestamp 1636968456
transform 1 0 104328 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1134
timestamp 1636968456
transform 1 0 105432 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1146
timestamp 1636968456
transform 1 0 106536 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_1158
timestamp 1
transform 1 0 107640 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_1166
timestamp 1
transform 1 0 108376 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1636968456
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1636968456
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636968456
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1636968456
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1636968456
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_65
timestamp 1
transform 1 0 7084 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1122
timestamp 1636968456
transform 1 0 104328 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1134
timestamp 1636968456
transform 1 0 105432 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_1146
timestamp 1
transform 1 0 106536 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1148
timestamp 1636968456
transform 1 0 106720 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_1160
timestamp 1
transform 1 0 107824 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636968456
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636968456
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636968456
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1636968456
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1636968456
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_69
timestamp 1
transform 1 0 7452 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1122
timestamp 1636968456
transform 1 0 104328 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1134
timestamp 1636968456
transform 1 0 105432 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1146
timestamp 1636968456
transform 1 0 106536 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_1158
timestamp 1
transform 1 0 107640 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_1166
timestamp 1
transform 1 0 108376 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636968456
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636968456
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636968456
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1636968456
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1636968456
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_65
timestamp 1
transform 1 0 7084 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1122
timestamp 1636968456
transform 1 0 104328 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1134
timestamp 1636968456
transform 1 0 105432 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1146
timestamp 1
transform 1 0 106536 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1148
timestamp 1636968456
transform 1 0 106720 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_1160
timestamp 1
transform 1 0 107824 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636968456
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1636968456
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1636968456
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1636968456
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1636968456
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_69
timestamp 1
transform 1 0 7452 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1122
timestamp 1636968456
transform 1 0 104328 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1134
timestamp 1636968456
transform 1 0 105432 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1146
timestamp 1636968456
transform 1 0 106536 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_1158
timestamp 1
transform 1 0 107640 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_1166
timestamp 1
transform 1 0 108376 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636968456
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636968456
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1636968456
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1636968456
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1636968456
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_65
timestamp 1
transform 1 0 7084 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1122
timestamp 1636968456
transform 1 0 104328 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1134
timestamp 1636968456
transform 1 0 105432 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_1146
timestamp 1
transform 1 0 106536 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1148
timestamp 1636968456
transform 1 0 106720 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_1160
timestamp 1
transform 1 0 107824 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1636968456
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1636968456
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1636968456
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1636968456
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1636968456
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_69
timestamp 1
transform 1 0 7452 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1122
timestamp 1636968456
transform 1 0 104328 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1134
timestamp 1636968456
transform 1 0 105432 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1146
timestamp 1636968456
transform 1 0 106536 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_1158
timestamp 1
transform 1 0 107640 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_1166
timestamp 1
transform 1 0 108376 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636968456
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636968456
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1636968456
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1636968456
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1636968456
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_65
timestamp 1
transform 1 0 7084 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1122
timestamp 1636968456
transform 1 0 104328 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1134
timestamp 1636968456
transform 1 0 105432 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_1146
timestamp 1
transform 1 0 106536 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1148
timestamp 1636968456
transform 1 0 106720 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_1160
timestamp 1
transform 1 0 107824 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636968456
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636968456
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1636968456
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1636968456
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1636968456
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_69
timestamp 1
transform 1 0 7452 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1122
timestamp 1636968456
transform 1 0 104328 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1134
timestamp 1636968456
transform 1 0 105432 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1146
timestamp 1636968456
transform 1 0 106536 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_1158
timestamp 1
transform 1 0 107640 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_1166
timestamp 1
transform 1 0 108376 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636968456
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636968456
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1636968456
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1636968456
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1636968456
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_65
timestamp 1
transform 1 0 7084 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1122
timestamp 1636968456
transform 1 0 104328 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1134
timestamp 1636968456
transform 1 0 105432 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_1146
timestamp 1
transform 1 0 106536 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1148
timestamp 1636968456
transform 1 0 106720 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_1160
timestamp 1
transform 1 0 107824 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1636968456
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1636968456
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1636968456
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1636968456
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1636968456
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_69
timestamp 1
transform 1 0 7452 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1122
timestamp 1636968456
transform 1 0 104328 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1134
timestamp 1636968456
transform 1 0 105432 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1146
timestamp 1636968456
transform 1 0 106536 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_1158
timestamp 1
transform 1 0 107640 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_1166
timestamp 1
transform 1 0 108376 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1636968456
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1636968456
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1636968456
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1636968456
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1636968456
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_65
timestamp 1
transform 1 0 7084 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1122
timestamp 1636968456
transform 1 0 104328 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1134
timestamp 1636968456
transform 1 0 105432 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_1146
timestamp 1
transform 1 0 106536 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1148
timestamp 1636968456
transform 1 0 106720 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_1160
timestamp 1
transform 1 0 107824 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636968456
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636968456
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1636968456
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1636968456
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1636968456
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_69
timestamp 1
transform 1 0 7452 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1122
timestamp 1636968456
transform 1 0 104328 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1134
timestamp 1636968456
transform 1 0 105432 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1146
timestamp 1636968456
transform 1 0 106536 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_1158
timestamp 1
transform 1 0 107640 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_1166
timestamp 1
transform 1 0 108376 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636968456
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1636968456
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1636968456
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1636968456
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1636968456
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_65
timestamp 1
transform 1 0 7084 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1122
timestamp 1636968456
transform 1 0 104328 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1134
timestamp 1636968456
transform 1 0 105432 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_1146
timestamp 1
transform 1 0 106536 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1148
timestamp 1636968456
transform 1 0 106720 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_1160
timestamp 1
transform 1 0 107824 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1636968456
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1636968456
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1636968456
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1636968456
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1636968456
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_69
timestamp 1
transform 1 0 7452 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1122
timestamp 1636968456
transform 1 0 104328 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1134
timestamp 1636968456
transform 1 0 105432 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1146
timestamp 1636968456
transform 1 0 106536 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_1158
timestamp 1
transform 1 0 107640 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_1166
timestamp 1
transform 1 0 108376 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1636968456
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1636968456
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1636968456
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1636968456
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1636968456
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_65
timestamp 1
transform 1 0 7084 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1122
timestamp 1636968456
transform 1 0 104328 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1134
timestamp 1636968456
transform 1 0 105432 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_1146
timestamp 1
transform 1 0 106536 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1148
timestamp 1636968456
transform 1 0 106720 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_1160
timestamp 1
transform 1 0 107824 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1636968456
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1636968456
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1636968456
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1636968456
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1636968456
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_69
timestamp 1
transform 1 0 7452 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1122
timestamp 1636968456
transform 1 0 104328 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1134
timestamp 1636968456
transform 1 0 105432 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1146
timestamp 1636968456
transform 1 0 106536 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_1158
timestamp 1
transform 1 0 107640 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_1166
timestamp 1
transform 1 0 108376 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1636968456
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1636968456
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1636968456
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1636968456
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1636968456
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_65
timestamp 1
transform 1 0 7084 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1122
timestamp 1636968456
transform 1 0 104328 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1134
timestamp 1636968456
transform 1 0 105432 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_1146
timestamp 1
transform 1 0 106536 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1148
timestamp 1636968456
transform 1 0 106720 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_1160
timestamp 1
transform 1 0 107824 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1636968456
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1636968456
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1636968456
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1636968456
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1636968456
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_69
timestamp 1
transform 1 0 7452 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1122
timestamp 1636968456
transform 1 0 104328 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1134
timestamp 1636968456
transform 1 0 105432 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1146
timestamp 1636968456
transform 1 0 106536 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_1158
timestamp 1
transform 1 0 107640 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_1166
timestamp 1
transform 1 0 108376 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1636968456
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1636968456
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1636968456
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1636968456
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1636968456
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_65
timestamp 1
transform 1 0 7084 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1122
timestamp 1636968456
transform 1 0 104328 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1134
timestamp 1636968456
transform 1 0 105432 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_1146
timestamp 1
transform 1 0 106536 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1148
timestamp 1636968456
transform 1 0 106720 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_1160
timestamp 1
transform 1 0 107824 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1636968456
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1636968456
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1636968456
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1636968456
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1636968456
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_69
timestamp 1
transform 1 0 7452 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1122
timestamp 1636968456
transform 1 0 104328 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1134
timestamp 1636968456
transform 1 0 105432 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1146
timestamp 1636968456
transform 1 0 106536 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_1158
timestamp 1
transform 1 0 107640 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_1166
timestamp 1
transform 1 0 108376 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1636968456
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1636968456
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1636968456
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1636968456
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1636968456
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_65
timestamp 1
transform 1 0 7084 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1122
timestamp 1636968456
transform 1 0 104328 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1134
timestamp 1636968456
transform 1 0 105432 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_1146
timestamp 1
transform 1 0 106536 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1148
timestamp 1636968456
transform 1 0 106720 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_1160
timestamp 1
transform 1 0 107824 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1636968456
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1636968456
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1636968456
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1636968456
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1636968456
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_69
timestamp 1
transform 1 0 7452 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1122
timestamp 1636968456
transform 1 0 104328 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1134
timestamp 1636968456
transform 1 0 105432 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1146
timestamp 1636968456
transform 1 0 106536 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_1158
timestamp 1
transform 1 0 107640 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_1166
timestamp 1
transform 1 0 108376 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1636968456
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1636968456
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1636968456
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1636968456
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1636968456
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_65
timestamp 1
transform 1 0 7084 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1122
timestamp 1636968456
transform 1 0 104328 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1134
timestamp 1636968456
transform 1 0 105432 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_1146
timestamp 1
transform 1 0 106536 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1148
timestamp 1636968456
transform 1 0 106720 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_1160
timestamp 1
transform 1 0 107824 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1636968456
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1636968456
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1636968456
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1636968456
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1636968456
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_69
timestamp 1
transform 1 0 7452 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1122
timestamp 1636968456
transform 1 0 104328 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1134
timestamp 1636968456
transform 1 0 105432 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1146
timestamp 1636968456
transform 1 0 106536 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_1158
timestamp 1
transform 1 0 107640 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_1166
timestamp 1
transform 1 0 108376 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1636968456
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1636968456
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1636968456
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1636968456
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1636968456
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_65
timestamp 1
transform 1 0 7084 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1122
timestamp 1636968456
transform 1 0 104328 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1134
timestamp 1636968456
transform 1 0 105432 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_1146
timestamp 1
transform 1 0 106536 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1148
timestamp 1636968456
transform 1 0 106720 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_1160
timestamp 1
transform 1 0 107824 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1636968456
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1636968456
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1636968456
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1636968456
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1636968456
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_69
timestamp 1
transform 1 0 7452 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1122
timestamp 1636968456
transform 1 0 104328 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1134
timestamp 1636968456
transform 1 0 105432 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1146
timestamp 1636968456
transform 1 0 106536 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_1158
timestamp 1
transform 1 0 107640 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_1166
timestamp 1
transform 1 0 108376 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1636968456
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1636968456
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1636968456
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1636968456
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1636968456
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_65
timestamp 1
transform 1 0 7084 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1122
timestamp 1636968456
transform 1 0 104328 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1134
timestamp 1636968456
transform 1 0 105432 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_1146
timestamp 1
transform 1 0 106536 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1148
timestamp 1636968456
transform 1 0 106720 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_1160
timestamp 1
transform 1 0 107824 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1636968456
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1636968456
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1636968456
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1636968456
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1636968456
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_69
timestamp 1
transform 1 0 7452 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1122
timestamp 1636968456
transform 1 0 104328 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1134
timestamp 1636968456
transform 1 0 105432 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1146
timestamp 1636968456
transform 1 0 106536 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_1158
timestamp 1
transform 1 0 107640 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_1166
timestamp 1
transform 1 0 108376 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1636968456
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1636968456
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1636968456
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1636968456
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1636968456
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_65
timestamp 1
transform 1 0 7084 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1122
timestamp 1636968456
transform 1 0 104328 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1134
timestamp 1636968456
transform 1 0 105432 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_1146
timestamp 1
transform 1 0 106536 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1148
timestamp 1636968456
transform 1 0 106720 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_1160
timestamp 1
transform 1 0 107824 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1636968456
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1636968456
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_27
timestamp 1636968456
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_39
timestamp 1636968456
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1636968456
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_69
timestamp 1
transform 1 0 7452 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1122
timestamp 1636968456
transform 1 0 104328 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1134
timestamp 1636968456
transform 1 0 105432 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1146
timestamp 1636968456
transform 1 0 106536 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_1158
timestamp 1
transform 1 0 107640 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_1166
timestamp 1
transform 1 0 108376 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_3
timestamp 1636968456
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_15
timestamp 1636968456
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1636968456
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1636968456
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1636968456
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_65
timestamp 1
transform 1 0 7084 0 1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1122
timestamp 1636968456
transform 1 0 104328 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1134
timestamp 1636968456
transform 1 0 105432 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_1146
timestamp 1
transform 1 0 106536 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1148
timestamp 1636968456
transform 1 0 106720 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_1160
timestamp 1
transform 1 0 107824 0 1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1636968456
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1636968456
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_27
timestamp 1636968456
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_39
timestamp 1636968456
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_51
timestamp 1
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1636968456
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_69
timestamp 1
transform 1 0 7452 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1122
timestamp 1636968456
transform 1 0 104328 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1134
timestamp 1636968456
transform 1 0 105432 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1146
timestamp 1636968456
transform 1 0 106536 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_1158
timestamp 1
transform 1 0 107640 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_103_1166
timestamp 1
transform 1 0 108376 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_3
timestamp 1636968456
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_15
timestamp 1636968456
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1636968456
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1636968456
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1636968456
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_65
timestamp 1
transform 1 0 7084 0 1 58752
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1122
timestamp 1636968456
transform 1 0 104328 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1134
timestamp 1636968456
transform 1 0 105432 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_1146
timestamp 1
transform 1 0 106536 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1148
timestamp 1636968456
transform 1 0 106720 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_1160
timestamp 1
transform 1 0 107824 0 1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_105_3
timestamp 1636968456
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_15
timestamp 1636968456
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_27
timestamp 1636968456
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_39
timestamp 1636968456
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_105_57
timestamp 1
transform 1 0 6348 0 -1 59840
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1122
timestamp 1636968456
transform 1 0 104328 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1134
timestamp 1636968456
transform 1 0 105432 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1146
timestamp 1636968456
transform 1 0 106536 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_1158
timestamp 1
transform 1 0 107640 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_1166
timestamp 1
transform 1 0 108376 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1636968456
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1636968456
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1636968456
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_41
timestamp 1
transform 1 0 4876 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_49
timestamp 1
transform 1 0 5612 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1125
timestamp 1636968456
transform 1 0 104604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_1137
timestamp 1
transform 1 0 105708 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_1145
timestamp 1
transform 1 0 106444 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1148
timestamp 1636968456
transform 1 0 106720 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_1160
timestamp 1
transform 1 0 107824 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_107_3
timestamp 1636968456
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_15
timestamp 1636968456
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_27
timestamp 1636968456
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_39
timestamp 1636968456
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_51
timestamp 1
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_57
timestamp 1
transform 1 0 6348 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_65
timestamp 1
transform 1 0 7084 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1122
timestamp 1636968456
transform 1 0 104328 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1134
timestamp 1636968456
transform 1 0 105432 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1146
timestamp 1636968456
transform 1 0 106536 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_1158
timestamp 1
transform 1 0 107640 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_1166
timestamp 1
transform 1 0 108376 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1636968456
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1636968456
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1636968456
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_41
timestamp 1636968456
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_53
timestamp 1636968456
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_65
timestamp 1
transform 1 0 7084 0 1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1122
timestamp 1636968456
transform 1 0 104328 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1134
timestamp 1636968456
transform 1 0 105432 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_1146
timestamp 1
transform 1 0 106536 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1148
timestamp 1636968456
transform 1 0 106720 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_1160
timestamp 1
transform 1 0 107824 0 1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_109_3
timestamp 1636968456
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_15
timestamp 1636968456
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_27
timestamp 1636968456
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_39
timestamp 1636968456
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_51
timestamp 1
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_57
timestamp 1636968456
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_69
timestamp 1
transform 1 0 7452 0 -1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1122
timestamp 1636968456
transform 1 0 104328 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1134
timestamp 1636968456
transform 1 0 105432 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1146
timestamp 1636968456
transform 1 0 106536 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_1158
timestamp 1
transform 1 0 107640 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_1166
timestamp 1
transform 1 0 108376 0 -1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_110_3
timestamp 1636968456
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_15
timestamp 1636968456
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_29
timestamp 1636968456
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_41
timestamp 1636968456
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_53
timestamp 1636968456
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_65
timestamp 1
transform 1 0 7084 0 1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1122
timestamp 1636968456
transform 1 0 104328 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1134
timestamp 1636968456
transform 1 0 105432 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_1146
timestamp 1
transform 1 0 106536 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1148
timestamp 1636968456
transform 1 0 106720 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_1160
timestamp 1
transform 1 0 107824 0 1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1636968456
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1636968456
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_27
timestamp 1636968456
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_39
timestamp 1636968456
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_51
timestamp 1
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_57
timestamp 1636968456
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_69
timestamp 1
transform 1 0 7452 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1122
timestamp 1636968456
transform 1 0 104328 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1134
timestamp 1636968456
transform 1 0 105432 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1146
timestamp 1636968456
transform 1 0 106536 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_1158
timestamp 1
transform 1 0 107640 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_111_1166
timestamp 1
transform 1 0 108376 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_112_3
timestamp 1636968456
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_15
timestamp 1636968456
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1636968456
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_41
timestamp 1636968456
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_53
timestamp 1636968456
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_65
timestamp 1
transform 1 0 7084 0 1 63104
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1122
timestamp 1636968456
transform 1 0 104328 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1134
timestamp 1636968456
transform 1 0 105432 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_1146
timestamp 1
transform 1 0 106536 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1148
timestamp 1636968456
transform 1 0 106720 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_1160
timestamp 1
transform 1 0 107824 0 1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1636968456
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1636968456
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_27
timestamp 1636968456
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_39
timestamp 1636968456
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_57
timestamp 1636968456
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_113_69
timestamp 1
transform 1 0 7452 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1122
timestamp 1636968456
transform 1 0 104328 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1134
timestamp 1636968456
transform 1 0 105432 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1146
timestamp 1636968456
transform 1 0 106536 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_1158
timestamp 1
transform 1 0 107640 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_113_1166
timestamp 1
transform 1 0 108376 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_114_3
timestamp 1636968456
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_15
timestamp 1636968456
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1636968456
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_41
timestamp 1636968456
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_53
timestamp 1636968456
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_65
timestamp 1
transform 1 0 7084 0 1 64192
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1122
timestamp 1636968456
transform 1 0 104328 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1134
timestamp 1636968456
transform 1 0 105432 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_1146
timestamp 1
transform 1 0 106536 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1148
timestamp 1636968456
transform 1 0 106720 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_1160
timestamp 1
transform 1 0 107824 0 1 64192
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_115_3
timestamp 1636968456
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_15
timestamp 1636968456
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_27
timestamp 1636968456
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_39
timestamp 1636968456
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_51
timestamp 1
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_57
timestamp 1636968456
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_115_69
timestamp 1
transform 1 0 7452 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1122
timestamp 1636968456
transform 1 0 104328 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1134
timestamp 1636968456
transform 1 0 105432 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1146
timestamp 1636968456
transform 1 0 106536 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_1158
timestamp 1
transform 1 0 107640 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_115_1166
timestamp 1
transform 1 0 108376 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1636968456
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1636968456
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_29
timestamp 1636968456
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_41
timestamp 1636968456
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_53
timestamp 1636968456
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_65
timestamp 1
transform 1 0 7084 0 1 65280
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1122
timestamp 1636968456
transform 1 0 104328 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1134
timestamp 1636968456
transform 1 0 105432 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_1146
timestamp 1
transform 1 0 106536 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1148
timestamp 1636968456
transform 1 0 106720 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_1160
timestamp 1
transform 1 0 107824 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_117_3
timestamp 1636968456
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_15
timestamp 1636968456
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_27
timestamp 1
transform 1 0 3588 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_29
timestamp 1636968456
transform 1 0 3772 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_41
timestamp 1636968456
transform 1 0 4876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_53
timestamp 1
transform 1 0 5980 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_57
timestamp 1636968456
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_69
timestamp 1636968456
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_81
timestamp 1
transform 1 0 8556 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_85
timestamp 1636968456
transform 1 0 8924 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_97
timestamp 1636968456
transform 1 0 10028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_109
timestamp 1
transform 1 0 11132 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_113
timestamp 1636968456
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_125
timestamp 1636968456
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_137
timestamp 1
transform 1 0 13708 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_141
timestamp 1636968456
transform 1 0 14076 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_153
timestamp 1636968456
transform 1 0 15180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_165
timestamp 1
transform 1 0 16284 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_169
timestamp 1636968456
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_181
timestamp 1636968456
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_193
timestamp 1
transform 1 0 18860 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_197
timestamp 1636968456
transform 1 0 19228 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_209
timestamp 1636968456
transform 1 0 20332 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_221
timestamp 1
transform 1 0 21436 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_225
timestamp 1636968456
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_237
timestamp 1636968456
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_249
timestamp 1
transform 1 0 24012 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_253
timestamp 1636968456
transform 1 0 24380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_265
timestamp 1636968456
transform 1 0 25484 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_277
timestamp 1
transform 1 0 26588 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_281
timestamp 1636968456
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_293
timestamp 1636968456
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_305
timestamp 1
transform 1 0 29164 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_309
timestamp 1636968456
transform 1 0 29532 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_321
timestamp 1636968456
transform 1 0 30636 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_333
timestamp 1
transform 1 0 31740 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_337
timestamp 1636968456
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_349
timestamp 1636968456
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_361
timestamp 1
transform 1 0 34316 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_365
timestamp 1636968456
transform 1 0 34684 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_377
timestamp 1
transform 1 0 35788 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_117_382
timestamp 1
transform 1 0 36248 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_390
timestamp 1
transform 1 0 36984 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_393
timestamp 1636968456
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_405
timestamp 1
transform 1 0 38364 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_117_410
timestamp 1
transform 1 0 38824 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_418
timestamp 1
transform 1 0 39560 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_421
timestamp 1636968456
transform 1 0 39836 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_117_433
timestamp 1
transform 1 0 40940 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_117_437
timestamp 1
transform 1 0 41308 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_117_445
timestamp 1
transform 1 0 42044 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_449
timestamp 1636968456
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_461
timestamp 1
transform 1 0 43516 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_464
timestamp 1636968456
transform 1 0 43792 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_477
timestamp 1636968456
transform 1 0 44988 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_491
timestamp 1636968456
transform 1 0 46276 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_503
timestamp 1
transform 1 0 47380 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_505
timestamp 1
transform 1 0 47564 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_117_513
timestamp 1
transform 1 0 48300 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_518
timestamp 1636968456
transform 1 0 48760 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_117_530
timestamp 1
transform 1 0 49864 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_117_533
timestamp 1
transform 1 0 50140 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_541
timestamp 1
transform 1 0 50876 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_545
timestamp 1636968456
transform 1 0 51244 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_557
timestamp 1
transform 1 0 52348 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_117_561
timestamp 1
transform 1 0 52716 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_117_569
timestamp 1
transform 1 0 53452 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_572
timestamp 1636968456
transform 1 0 53728 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_584
timestamp 1
transform 1 0 54832 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_117_589
timestamp 1
transform 1 0 55292 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_117_597
timestamp 1
transform 1 0 56028 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_600
timestamp 1636968456
transform 1 0 56304 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_612
timestamp 1
transform 1 0 57408 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_117_617
timestamp 1
transform 1 0 57868 0 -1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_117_627
timestamp 1636968456
transform 1 0 58788 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_639
timestamp 1
transform 1 0 59892 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_643
timestamp 1
transform 1 0 60260 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_117_645
timestamp 1
transform 1 0 60444 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_651
timestamp 1
transform 1 0 60996 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_654
timestamp 1636968456
transform 1 0 61272 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_666
timestamp 1
transform 1 0 62376 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_117_673
timestamp 1
transform 1 0 63020 0 -1 66368
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_117_681
timestamp 1636968456
transform 1 0 63756 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_693
timestamp 1
transform 1 0 64860 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_699
timestamp 1
transform 1 0 65412 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_701
timestamp 1
transform 1 0 65596 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_705
timestamp 1
transform 1 0 65964 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_708
timestamp 1636968456
transform 1 0 66240 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_720
timestamp 1
transform 1 0 67344 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_117_729
timestamp 1
transform 1 0 68172 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_117_735
timestamp 1636968456
transform 1 0 68724 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_747
timestamp 1
transform 1 0 69828 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_117_755
timestamp 1
transform 1 0 70564 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_117_757
timestamp 1
transform 1 0 70748 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_762
timestamp 1636968456
transform 1 0 71208 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_774
timestamp 1
transform 1 0 72312 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_782
timestamp 1
transform 1 0 73048 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_117_785
timestamp 1
transform 1 0 73324 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_789
timestamp 1636968456
transform 1 0 73692 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_801
timestamp 1
transform 1 0 74796 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_117_809
timestamp 1
transform 1 0 75532 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_813
timestamp 1636968456
transform 1 0 75900 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_825
timestamp 1636968456
transform 1 0 77004 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_837
timestamp 1
transform 1 0 78108 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_841
timestamp 1636968456
transform 1 0 78476 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_853
timestamp 1636968456
transform 1 0 79580 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_865
timestamp 1
transform 1 0 80684 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_869
timestamp 1636968456
transform 1 0 81052 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_881
timestamp 1636968456
transform 1 0 82156 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_893
timestamp 1
transform 1 0 83260 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_897
timestamp 1636968456
transform 1 0 83628 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_909
timestamp 1
transform 1 0 84732 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_913
timestamp 1
transform 1 0 85100 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_920
timestamp 1
transform 1 0 85744 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_117_992
timestamp 1636968456
transform 1 0 92368 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_1004
timestamp 1
transform 1 0 93472 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1009
timestamp 1
transform 1 0 93932 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1039
timestamp 1636968456
transform 1 0 96692 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1051
timestamp 1636968456
transform 1 0 97796 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1063
timestamp 1
transform 1 0 98900 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1065
timestamp 1636968456
transform 1 0 99084 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1077
timestamp 1636968456
transform 1 0 100188 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1089
timestamp 1
transform 1 0 101292 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1093
timestamp 1636968456
transform 1 0 101660 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1105
timestamp 1636968456
transform 1 0 102764 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1117
timestamp 1
transform 1 0 103868 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1121
timestamp 1636968456
transform 1 0 104236 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1133
timestamp 1636968456
transform 1 0 105340 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1145
timestamp 1
transform 1 0 106444 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1149
timestamp 1636968456
transform 1 0 106812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_1161
timestamp 1
transform 1 0 107916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1167
timestamp 1
transform 1 0 108468 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1636968456
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1636968456
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1636968456
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_41
timestamp 1636968456
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_53
timestamp 1636968456
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_65
timestamp 1636968456
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_85
timestamp 1636968456
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_97
timestamp 1636968456
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_109
timestamp 1636968456
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_121
timestamp 1636968456
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_141
timestamp 1636968456
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_153
timestamp 1636968456
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_165
timestamp 1636968456
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_177
timestamp 1636968456
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_189
timestamp 1
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_195
timestamp 1
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_197
timestamp 1636968456
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_209
timestamp 1636968456
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_221
timestamp 1636968456
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_233
timestamp 1636968456
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_245
timestamp 1
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_251
timestamp 1
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_253
timestamp 1636968456
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_265
timestamp 1636968456
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_277
timestamp 1636968456
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_289
timestamp 1636968456
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_301
timestamp 1
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_307
timestamp 1
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_309
timestamp 1636968456
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_321
timestamp 1636968456
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_333
timestamp 1636968456
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_345
timestamp 1636968456
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_357
timestamp 1
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_363
timestamp 1
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_365
timestamp 1636968456
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_377
timestamp 1636968456
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_389
timestamp 1636968456
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_401
timestamp 1636968456
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_413
timestamp 1
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_419
timestamp 1
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_421
timestamp 1636968456
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_433
timestamp 1636968456
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_445
timestamp 1636968456
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_457
timestamp 1636968456
transform 1 0 43148 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_469
timestamp 1
transform 1 0 44252 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_475
timestamp 1
transform 1 0 44804 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_477
timestamp 1636968456
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_489
timestamp 1636968456
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_501
timestamp 1636968456
transform 1 0 47196 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_513
timestamp 1636968456
transform 1 0 48300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_525
timestamp 1
transform 1 0 49404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_531
timestamp 1
transform 1 0 49956 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_533
timestamp 1636968456
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_545
timestamp 1636968456
transform 1 0 51244 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_557
timestamp 1636968456
transform 1 0 52348 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_569
timestamp 1636968456
transform 1 0 53452 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_581
timestamp 1
transform 1 0 54556 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_587
timestamp 1
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_589
timestamp 1636968456
transform 1 0 55292 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_601
timestamp 1636968456
transform 1 0 56396 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_613
timestamp 1636968456
transform 1 0 57500 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_625
timestamp 1636968456
transform 1 0 58604 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_637
timestamp 1
transform 1 0 59708 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_643
timestamp 1
transform 1 0 60260 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_645
timestamp 1636968456
transform 1 0 60444 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_657
timestamp 1636968456
transform 1 0 61548 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_669
timestamp 1636968456
transform 1 0 62652 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_681
timestamp 1636968456
transform 1 0 63756 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_693
timestamp 1
transform 1 0 64860 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_699
timestamp 1
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_701
timestamp 1636968456
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_713
timestamp 1636968456
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_725
timestamp 1636968456
transform 1 0 67804 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_737
timestamp 1636968456
transform 1 0 68908 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_749
timestamp 1
transform 1 0 70012 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_755
timestamp 1
transform 1 0 70564 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_757
timestamp 1636968456
transform 1 0 70748 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_769
timestamp 1636968456
transform 1 0 71852 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_781
timestamp 1636968456
transform 1 0 72956 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_793
timestamp 1636968456
transform 1 0 74060 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_805
timestamp 1
transform 1 0 75164 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_811
timestamp 1
transform 1 0 75716 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_813
timestamp 1636968456
transform 1 0 75900 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_825
timestamp 1636968456
transform 1 0 77004 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_837
timestamp 1636968456
transform 1 0 78108 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_849
timestamp 1636968456
transform 1 0 79212 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_861
timestamp 1
transform 1 0 80316 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_867
timestamp 1
transform 1 0 80868 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_869
timestamp 1636968456
transform 1 0 81052 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_881
timestamp 1636968456
transform 1 0 82156 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_893
timestamp 1
transform 1 0 83260 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_118_921
timestamp 1
transform 1 0 85836 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_118_925
timestamp 1
transform 1 0 86204 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_933
timestamp 1
transform 1 0 86940 0 1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_118_988
timestamp 1636968456
transform 1 0 92000 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1000
timestamp 1636968456
transform 1 0 93104 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1012
timestamp 1636968456
transform 1 0 94208 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1024
timestamp 1636968456
transform 1 0 95312 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1037
timestamp 1636968456
transform 1 0 96508 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1049
timestamp 1636968456
transform 1 0 97612 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1061
timestamp 1636968456
transform 1 0 98716 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1073
timestamp 1636968456
transform 1 0 99820 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1085
timestamp 1
transform 1 0 100924 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1091
timestamp 1
transform 1 0 101476 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1093
timestamp 1636968456
transform 1 0 101660 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1105
timestamp 1636968456
transform 1 0 102764 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1117
timestamp 1636968456
transform 1 0 103868 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1129
timestamp 1636968456
transform 1 0 104972 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1141
timestamp 1
transform 1 0 106076 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1147
timestamp 1
transform 1 0 106628 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1149
timestamp 1636968456
transform 1 0 106812 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1161
timestamp 1
transform 1 0 107916 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1167
timestamp 1
transform 1 0 108468 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_3
timestamp 1636968456
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_15
timestamp 1636968456
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_27
timestamp 1636968456
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_39
timestamp 1636968456
transform 1 0 4692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_51
timestamp 1
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_57
timestamp 1636968456
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_69
timestamp 1636968456
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_81
timestamp 1636968456
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_93
timestamp 1636968456
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_113
timestamp 1636968456
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_125
timestamp 1636968456
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_137
timestamp 1636968456
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_149
timestamp 1636968456
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_169
timestamp 1636968456
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_181
timestamp 1636968456
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_193
timestamp 1636968456
transform 1 0 18860 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_205
timestamp 1636968456
transform 1 0 19964 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_217
timestamp 1
transform 1 0 21068 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_223
timestamp 1
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_225
timestamp 1636968456
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_237
timestamp 1636968456
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_249
timestamp 1636968456
transform 1 0 24012 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_261
timestamp 1636968456
transform 1 0 25116 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_273
timestamp 1
transform 1 0 26220 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_279
timestamp 1
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_281
timestamp 1636968456
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_293
timestamp 1636968456
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_305
timestamp 1636968456
transform 1 0 29164 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_317
timestamp 1636968456
transform 1 0 30268 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_329
timestamp 1
transform 1 0 31372 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_335
timestamp 1
transform 1 0 31924 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_337
timestamp 1636968456
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_349
timestamp 1636968456
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_361
timestamp 1636968456
transform 1 0 34316 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_373
timestamp 1636968456
transform 1 0 35420 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_385
timestamp 1
transform 1 0 36524 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_391
timestamp 1
transform 1 0 37076 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_393
timestamp 1636968456
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_405
timestamp 1636968456
transform 1 0 38364 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_417
timestamp 1636968456
transform 1 0 39468 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_429
timestamp 1636968456
transform 1 0 40572 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_441
timestamp 1
transform 1 0 41676 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_447
timestamp 1
transform 1 0 42228 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_449
timestamp 1636968456
transform 1 0 42412 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_461
timestamp 1636968456
transform 1 0 43516 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_473
timestamp 1636968456
transform 1 0 44620 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_485
timestamp 1636968456
transform 1 0 45724 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_497
timestamp 1
transform 1 0 46828 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_503
timestamp 1
transform 1 0 47380 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_505
timestamp 1636968456
transform 1 0 47564 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_517
timestamp 1636968456
transform 1 0 48668 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_529
timestamp 1636968456
transform 1 0 49772 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_541
timestamp 1636968456
transform 1 0 50876 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_553
timestamp 1
transform 1 0 51980 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_559
timestamp 1
transform 1 0 52532 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_561
timestamp 1636968456
transform 1 0 52716 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_573
timestamp 1636968456
transform 1 0 53820 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_585
timestamp 1636968456
transform 1 0 54924 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_597
timestamp 1636968456
transform 1 0 56028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_609
timestamp 1
transform 1 0 57132 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_615
timestamp 1
transform 1 0 57684 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_617
timestamp 1636968456
transform 1 0 57868 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_629
timestamp 1636968456
transform 1 0 58972 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_641
timestamp 1636968456
transform 1 0 60076 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_653
timestamp 1636968456
transform 1 0 61180 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_665
timestamp 1
transform 1 0 62284 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_671
timestamp 1
transform 1 0 62836 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_673
timestamp 1636968456
transform 1 0 63020 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_685
timestamp 1636968456
transform 1 0 64124 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_697
timestamp 1636968456
transform 1 0 65228 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_709
timestamp 1636968456
transform 1 0 66332 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_721
timestamp 1
transform 1 0 67436 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_727
timestamp 1
transform 1 0 67988 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_729
timestamp 1636968456
transform 1 0 68172 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_741
timestamp 1636968456
transform 1 0 69276 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_753
timestamp 1636968456
transform 1 0 70380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_765
timestamp 1636968456
transform 1 0 71484 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_777
timestamp 1
transform 1 0 72588 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_783
timestamp 1
transform 1 0 73140 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_785
timestamp 1636968456
transform 1 0 73324 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_797
timestamp 1636968456
transform 1 0 74428 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_809
timestamp 1636968456
transform 1 0 75532 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_821
timestamp 1636968456
transform 1 0 76636 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_833
timestamp 1
transform 1 0 77740 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_839
timestamp 1
transform 1 0 78292 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_841
timestamp 1636968456
transform 1 0 78476 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_853
timestamp 1636968456
transform 1 0 79580 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_865
timestamp 1636968456
transform 1 0 80684 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_877
timestamp 1636968456
transform 1 0 81788 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_889
timestamp 1
transform 1 0 82892 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_895
timestamp 1
transform 1 0 83444 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_119_897
timestamp 1
transform 1 0 83628 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_901
timestamp 1
transform 1 0 83996 0 -1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_119_908
timestamp 1636968456
transform 1 0 84640 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_920
timestamp 1
transform 1 0 85744 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_119_928
timestamp 1
transform 1 0 86480 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_119_988
timestamp 1636968456
transform 1 0 92000 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_1000
timestamp 1
transform 1 0 93104 0 -1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1009
timestamp 1636968456
transform 1 0 93932 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1021
timestamp 1636968456
transform 1 0 95036 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1033
timestamp 1636968456
transform 1 0 96140 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1045
timestamp 1636968456
transform 1 0 97244 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1057
timestamp 1
transform 1 0 98348 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1063
timestamp 1
transform 1 0 98900 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1065
timestamp 1636968456
transform 1 0 99084 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1077
timestamp 1636968456
transform 1 0 100188 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1089
timestamp 1636968456
transform 1 0 101292 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1101
timestamp 1636968456
transform 1 0 102396 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1113
timestamp 1
transform 1 0 103500 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1119
timestamp 1
transform 1 0 104052 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1121
timestamp 1636968456
transform 1 0 104236 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1133
timestamp 1636968456
transform 1 0 105340 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1145
timestamp 1636968456
transform 1 0 106444 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_1157
timestamp 1
transform 1 0 107548 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_1165
timestamp 1
transform 1 0 108284 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_3
timestamp 1636968456
transform 1 0 1380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_15
timestamp 1636968456
transform 1 0 2484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1636968456
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_41
timestamp 1636968456
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_53
timestamp 1636968456
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_65
timestamp 1636968456
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_85
timestamp 1636968456
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_97
timestamp 1636968456
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_109
timestamp 1636968456
transform 1 0 11132 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_121
timestamp 1636968456
transform 1 0 12236 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_133
timestamp 1
transform 1 0 13340 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_139
timestamp 1
transform 1 0 13892 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_141
timestamp 1636968456
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_153
timestamp 1636968456
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_165
timestamp 1636968456
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_177
timestamp 1636968456
transform 1 0 17388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_189
timestamp 1
transform 1 0 18492 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_195
timestamp 1
transform 1 0 19044 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_197
timestamp 1636968456
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_209
timestamp 1636968456
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_221
timestamp 1636968456
transform 1 0 21436 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_233
timestamp 1636968456
transform 1 0 22540 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_245
timestamp 1
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_251
timestamp 1
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_253
timestamp 1636968456
transform 1 0 24380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_265
timestamp 1636968456
transform 1 0 25484 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_277
timestamp 1636968456
transform 1 0 26588 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_289
timestamp 1636968456
transform 1 0 27692 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_301
timestamp 1
transform 1 0 28796 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_307
timestamp 1
transform 1 0 29348 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_309
timestamp 1636968456
transform 1 0 29532 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_321
timestamp 1636968456
transform 1 0 30636 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_333
timestamp 1636968456
transform 1 0 31740 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_345
timestamp 1636968456
transform 1 0 32844 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_357
timestamp 1
transform 1 0 33948 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_363
timestamp 1
transform 1 0 34500 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_365
timestamp 1636968456
transform 1 0 34684 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_377
timestamp 1636968456
transform 1 0 35788 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_389
timestamp 1636968456
transform 1 0 36892 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_401
timestamp 1636968456
transform 1 0 37996 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_413
timestamp 1
transform 1 0 39100 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_419
timestamp 1
transform 1 0 39652 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_421
timestamp 1636968456
transform 1 0 39836 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_433
timestamp 1636968456
transform 1 0 40940 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_445
timestamp 1636968456
transform 1 0 42044 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_457
timestamp 1636968456
transform 1 0 43148 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_469
timestamp 1
transform 1 0 44252 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_475
timestamp 1
transform 1 0 44804 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_477
timestamp 1636968456
transform 1 0 44988 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_489
timestamp 1636968456
transform 1 0 46092 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_501
timestamp 1636968456
transform 1 0 47196 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_513
timestamp 1636968456
transform 1 0 48300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_525
timestamp 1
transform 1 0 49404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_531
timestamp 1
transform 1 0 49956 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_533
timestamp 1636968456
transform 1 0 50140 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_545
timestamp 1636968456
transform 1 0 51244 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_557
timestamp 1636968456
transform 1 0 52348 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_569
timestamp 1636968456
transform 1 0 53452 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_581
timestamp 1
transform 1 0 54556 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_587
timestamp 1
transform 1 0 55108 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_589
timestamp 1636968456
transform 1 0 55292 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_601
timestamp 1636968456
transform 1 0 56396 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_613
timestamp 1636968456
transform 1 0 57500 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_625
timestamp 1636968456
transform 1 0 58604 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_637
timestamp 1
transform 1 0 59708 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_643
timestamp 1
transform 1 0 60260 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_645
timestamp 1636968456
transform 1 0 60444 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_657
timestamp 1636968456
transform 1 0 61548 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_669
timestamp 1636968456
transform 1 0 62652 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_681
timestamp 1636968456
transform 1 0 63756 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_693
timestamp 1
transform 1 0 64860 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_699
timestamp 1
transform 1 0 65412 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_701
timestamp 1636968456
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_713
timestamp 1636968456
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_725
timestamp 1636968456
transform 1 0 67804 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_737
timestamp 1636968456
transform 1 0 68908 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_749
timestamp 1
transform 1 0 70012 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_755
timestamp 1
transform 1 0 70564 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_757
timestamp 1636968456
transform 1 0 70748 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_769
timestamp 1636968456
transform 1 0 71852 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_781
timestamp 1636968456
transform 1 0 72956 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_793
timestamp 1636968456
transform 1 0 74060 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_805
timestamp 1
transform 1 0 75164 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_811
timestamp 1
transform 1 0 75716 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_813
timestamp 1636968456
transform 1 0 75900 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_825
timestamp 1636968456
transform 1 0 77004 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_837
timestamp 1636968456
transform 1 0 78108 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_849
timestamp 1636968456
transform 1 0 79212 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_861
timestamp 1
transform 1 0 80316 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_867
timestamp 1
transform 1 0 80868 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_869
timestamp 1636968456
transform 1 0 81052 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_881
timestamp 1636968456
transform 1 0 82156 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_893
timestamp 1636968456
transform 1 0 83260 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_905
timestamp 1636968456
transform 1 0 84364 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_917
timestamp 1
transform 1 0 85468 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_923
timestamp 1
transform 1 0 86020 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_928
timestamp 1636968456
transform 1 0 86480 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_940
timestamp 1
transform 1 0 87584 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_948
timestamp 1
transform 1 0 88320 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_120_954
timestamp 1
transform 1 0 88872 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_958
timestamp 1
transform 1 0 89240 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_120_973
timestamp 1
transform 1 0 90620 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_120_979
timestamp 1
transform 1 0 91172 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_981
timestamp 1
transform 1 0 91356 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_989
timestamp 1
transform 1 0 92092 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_998
timestamp 1636968456
transform 1 0 92920 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1010
timestamp 1636968456
transform 1 0 94024 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1022
timestamp 1636968456
transform 1 0 95128 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_120_1034
timestamp 1
transform 1 0 96232 0 1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1037
timestamp 1636968456
transform 1 0 96508 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1049
timestamp 1636968456
transform 1 0 97612 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1061
timestamp 1636968456
transform 1 0 98716 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1073
timestamp 1636968456
transform 1 0 99820 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_1085
timestamp 1
transform 1 0 100924 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1091
timestamp 1
transform 1 0 101476 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1093
timestamp 1636968456
transform 1 0 101660 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1105
timestamp 1636968456
transform 1 0 102764 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1117
timestamp 1636968456
transform 1 0 103868 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1129
timestamp 1636968456
transform 1 0 104972 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_1141
timestamp 1
transform 1 0 106076 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1147
timestamp 1
transform 1 0 106628 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1149
timestamp 1636968456
transform 1 0 106812 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1636968456
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1636968456
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_27
timestamp 1636968456
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_39
timestamp 1636968456
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_51
timestamp 1
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_57
timestamp 1636968456
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_69
timestamp 1636968456
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_81
timestamp 1636968456
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_93
timestamp 1636968456
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_113
timestamp 1636968456
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_125
timestamp 1636968456
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_137
timestamp 1636968456
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_149
timestamp 1636968456
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_161
timestamp 1
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_167
timestamp 1
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_169
timestamp 1636968456
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_181
timestamp 1636968456
transform 1 0 17756 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_193
timestamp 1636968456
transform 1 0 18860 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_205
timestamp 1636968456
transform 1 0 19964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_217
timestamp 1
transform 1 0 21068 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_223
timestamp 1
transform 1 0 21620 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_225
timestamp 1636968456
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_237
timestamp 1636968456
transform 1 0 22908 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_249
timestamp 1636968456
transform 1 0 24012 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_261
timestamp 1636968456
transform 1 0 25116 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_273
timestamp 1
transform 1 0 26220 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_279
timestamp 1
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_281
timestamp 1636968456
transform 1 0 26956 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_293
timestamp 1636968456
transform 1 0 28060 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_305
timestamp 1636968456
transform 1 0 29164 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_317
timestamp 1636968456
transform 1 0 30268 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_329
timestamp 1
transform 1 0 31372 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_335
timestamp 1
transform 1 0 31924 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_337
timestamp 1636968456
transform 1 0 32108 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_349
timestamp 1636968456
transform 1 0 33212 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_361
timestamp 1636968456
transform 1 0 34316 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_373
timestamp 1636968456
transform 1 0 35420 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_385
timestamp 1
transform 1 0 36524 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_391
timestamp 1
transform 1 0 37076 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_393
timestamp 1636968456
transform 1 0 37260 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_405
timestamp 1636968456
transform 1 0 38364 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_417
timestamp 1636968456
transform 1 0 39468 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_429
timestamp 1636968456
transform 1 0 40572 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_441
timestamp 1
transform 1 0 41676 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_447
timestamp 1
transform 1 0 42228 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_449
timestamp 1636968456
transform 1 0 42412 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_461
timestamp 1636968456
transform 1 0 43516 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_473
timestamp 1636968456
transform 1 0 44620 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_485
timestamp 1636968456
transform 1 0 45724 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_497
timestamp 1
transform 1 0 46828 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_503
timestamp 1
transform 1 0 47380 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_505
timestamp 1636968456
transform 1 0 47564 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_517
timestamp 1636968456
transform 1 0 48668 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_529
timestamp 1636968456
transform 1 0 49772 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_541
timestamp 1636968456
transform 1 0 50876 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_553
timestamp 1
transform 1 0 51980 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_559
timestamp 1
transform 1 0 52532 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_561
timestamp 1636968456
transform 1 0 52716 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_573
timestamp 1636968456
transform 1 0 53820 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_585
timestamp 1636968456
transform 1 0 54924 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_597
timestamp 1636968456
transform 1 0 56028 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_609
timestamp 1
transform 1 0 57132 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_615
timestamp 1
transform 1 0 57684 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_617
timestamp 1636968456
transform 1 0 57868 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_629
timestamp 1636968456
transform 1 0 58972 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_641
timestamp 1636968456
transform 1 0 60076 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_653
timestamp 1636968456
transform 1 0 61180 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_665
timestamp 1
transform 1 0 62284 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_671
timestamp 1
transform 1 0 62836 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_673
timestamp 1636968456
transform 1 0 63020 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_685
timestamp 1636968456
transform 1 0 64124 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_697
timestamp 1636968456
transform 1 0 65228 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_709
timestamp 1636968456
transform 1 0 66332 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_721
timestamp 1
transform 1 0 67436 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_727
timestamp 1
transform 1 0 67988 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_729
timestamp 1636968456
transform 1 0 68172 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_741
timestamp 1636968456
transform 1 0 69276 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_753
timestamp 1636968456
transform 1 0 70380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_765
timestamp 1636968456
transform 1 0 71484 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_777
timestamp 1
transform 1 0 72588 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_783
timestamp 1
transform 1 0 73140 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_785
timestamp 1636968456
transform 1 0 73324 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_797
timestamp 1636968456
transform 1 0 74428 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_809
timestamp 1636968456
transform 1 0 75532 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_821
timestamp 1636968456
transform 1 0 76636 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_833
timestamp 1
transform 1 0 77740 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_839
timestamp 1
transform 1 0 78292 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_841
timestamp 1636968456
transform 1 0 78476 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_853
timestamp 1636968456
transform 1 0 79580 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_865
timestamp 1636968456
transform 1 0 80684 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_877
timestamp 1636968456
transform 1 0 81788 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_889
timestamp 1
transform 1 0 82892 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_895
timestamp 1
transform 1 0 83444 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_897
timestamp 1636968456
transform 1 0 83628 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_909
timestamp 1636968456
transform 1 0 84732 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_921
timestamp 1
transform 1 0 85836 0 -1 68544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_121_932
timestamp 1636968456
transform 1 0 86848 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_944
timestamp 1
transform 1 0 87952 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_121_953
timestamp 1
transform 1 0 88780 0 -1 68544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_121_958
timestamp 1636968456
transform 1 0 89240 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_970
timestamp 1636968456
transform 1 0 90344 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_982
timestamp 1636968456
transform 1 0 91448 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_994
timestamp 1636968456
transform 1 0 92552 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_121_1006
timestamp 1
transform 1 0 93656 0 -1 68544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1009
timestamp 1636968456
transform 1 0 93932 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1021
timestamp 1636968456
transform 1 0 95036 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1033
timestamp 1636968456
transform 1 0 96140 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1045
timestamp 1636968456
transform 1 0 97244 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_1057
timestamp 1
transform 1 0 98348 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1063
timestamp 1
transform 1 0 98900 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1065
timestamp 1636968456
transform 1 0 99084 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1077
timestamp 1636968456
transform 1 0 100188 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1089
timestamp 1636968456
transform 1 0 101292 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1101
timestamp 1636968456
transform 1 0 102396 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_1113
timestamp 1
transform 1 0 103500 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1119
timestamp 1
transform 1 0 104052 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1121
timestamp 1636968456
transform 1 0 104236 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1133
timestamp 1636968456
transform 1 0 105340 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1145
timestamp 1636968456
transform 1 0 106444 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_1157
timestamp 1
transform 1 0 107548 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_121_1165
timestamp 1
transform 1 0 108284 0 -1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_122_3
timestamp 1636968456
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_15
timestamp 1636968456
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1636968456
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_41
timestamp 1636968456
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_53
timestamp 1636968456
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_65
timestamp 1636968456
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_85
timestamp 1636968456
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_97
timestamp 1636968456
transform 1 0 10028 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_109
timestamp 1636968456
transform 1 0 11132 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_121
timestamp 1636968456
transform 1 0 12236 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_133
timestamp 1
transform 1 0 13340 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_139
timestamp 1
transform 1 0 13892 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_141
timestamp 1636968456
transform 1 0 14076 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_153
timestamp 1636968456
transform 1 0 15180 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_165
timestamp 1636968456
transform 1 0 16284 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_177
timestamp 1636968456
transform 1 0 17388 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_189
timestamp 1
transform 1 0 18492 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_195
timestamp 1
transform 1 0 19044 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_197
timestamp 1636968456
transform 1 0 19228 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_209
timestamp 1636968456
transform 1 0 20332 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_221
timestamp 1636968456
transform 1 0 21436 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_233
timestamp 1636968456
transform 1 0 22540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_245
timestamp 1
transform 1 0 23644 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_251
timestamp 1
transform 1 0 24196 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_253
timestamp 1636968456
transform 1 0 24380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_265
timestamp 1636968456
transform 1 0 25484 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_277
timestamp 1636968456
transform 1 0 26588 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_289
timestamp 1636968456
transform 1 0 27692 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_301
timestamp 1
transform 1 0 28796 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_307
timestamp 1
transform 1 0 29348 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_309
timestamp 1636968456
transform 1 0 29532 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_321
timestamp 1636968456
transform 1 0 30636 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_333
timestamp 1636968456
transform 1 0 31740 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_345
timestamp 1636968456
transform 1 0 32844 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_357
timestamp 1
transform 1 0 33948 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_363
timestamp 1
transform 1 0 34500 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_365
timestamp 1636968456
transform 1 0 34684 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_377
timestamp 1636968456
transform 1 0 35788 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_389
timestamp 1636968456
transform 1 0 36892 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_401
timestamp 1636968456
transform 1 0 37996 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_413
timestamp 1
transform 1 0 39100 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_419
timestamp 1
transform 1 0 39652 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_421
timestamp 1636968456
transform 1 0 39836 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_433
timestamp 1636968456
transform 1 0 40940 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_445
timestamp 1636968456
transform 1 0 42044 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_457
timestamp 1636968456
transform 1 0 43148 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_469
timestamp 1
transform 1 0 44252 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_475
timestamp 1
transform 1 0 44804 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_477
timestamp 1636968456
transform 1 0 44988 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_489
timestamp 1636968456
transform 1 0 46092 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_501
timestamp 1636968456
transform 1 0 47196 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_513
timestamp 1636968456
transform 1 0 48300 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_525
timestamp 1
transform 1 0 49404 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_531
timestamp 1
transform 1 0 49956 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_533
timestamp 1636968456
transform 1 0 50140 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_545
timestamp 1636968456
transform 1 0 51244 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_557
timestamp 1636968456
transform 1 0 52348 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_569
timestamp 1636968456
transform 1 0 53452 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_581
timestamp 1
transform 1 0 54556 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_587
timestamp 1
transform 1 0 55108 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_589
timestamp 1636968456
transform 1 0 55292 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_601
timestamp 1636968456
transform 1 0 56396 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_613
timestamp 1636968456
transform 1 0 57500 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_625
timestamp 1636968456
transform 1 0 58604 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_637
timestamp 1
transform 1 0 59708 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_643
timestamp 1
transform 1 0 60260 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_645
timestamp 1636968456
transform 1 0 60444 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_657
timestamp 1636968456
transform 1 0 61548 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_669
timestamp 1636968456
transform 1 0 62652 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_681
timestamp 1636968456
transform 1 0 63756 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_693
timestamp 1
transform 1 0 64860 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_699
timestamp 1
transform 1 0 65412 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_701
timestamp 1636968456
transform 1 0 65596 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_713
timestamp 1636968456
transform 1 0 66700 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_725
timestamp 1636968456
transform 1 0 67804 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_737
timestamp 1636968456
transform 1 0 68908 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_749
timestamp 1
transform 1 0 70012 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_755
timestamp 1
transform 1 0 70564 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_757
timestamp 1636968456
transform 1 0 70748 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_769
timestamp 1636968456
transform 1 0 71852 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_781
timestamp 1636968456
transform 1 0 72956 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_793
timestamp 1636968456
transform 1 0 74060 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_805
timestamp 1
transform 1 0 75164 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_811
timestamp 1
transform 1 0 75716 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_813
timestamp 1636968456
transform 1 0 75900 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_825
timestamp 1636968456
transform 1 0 77004 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_837
timestamp 1636968456
transform 1 0 78108 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_849
timestamp 1636968456
transform 1 0 79212 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_861
timestamp 1
transform 1 0 80316 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_867
timestamp 1
transform 1 0 80868 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_869
timestamp 1636968456
transform 1 0 81052 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_881
timestamp 1636968456
transform 1 0 82156 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_893
timestamp 1636968456
transform 1 0 83260 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_905
timestamp 1636968456
transform 1 0 84364 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_917
timestamp 1
transform 1 0 85468 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_923
timestamp 1
transform 1 0 86020 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_925
timestamp 1636968456
transform 1 0 86204 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_937
timestamp 1636968456
transform 1 0 87308 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_949
timestamp 1
transform 1 0 88412 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_976
timestamp 1
transform 1 0 90896 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_122_981
timestamp 1
transform 1 0 91356 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_989
timestamp 1
transform 1 0 92092 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_993
timestamp 1636968456
transform 1 0 92460 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1005
timestamp 1636968456
transform 1 0 93564 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1017
timestamp 1636968456
transform 1 0 94668 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1029
timestamp 1
transform 1 0 95772 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1035
timestamp 1
transform 1 0 96324 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1037
timestamp 1636968456
transform 1 0 96508 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1049
timestamp 1636968456
transform 1 0 97612 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1061
timestamp 1636968456
transform 1 0 98716 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1073
timestamp 1636968456
transform 1 0 99820 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1085
timestamp 1
transform 1 0 100924 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1091
timestamp 1
transform 1 0 101476 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1093
timestamp 1636968456
transform 1 0 101660 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1105
timestamp 1636968456
transform 1 0 102764 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1117
timestamp 1636968456
transform 1 0 103868 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1129
timestamp 1636968456
transform 1 0 104972 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1141
timestamp 1
transform 1 0 106076 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1147
timestamp 1
transform 1 0 106628 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1149
timestamp 1636968456
transform 1 0 106812 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1161
timestamp 1
transform 1 0 107916 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1167
timestamp 1
transform 1 0 108468 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1636968456
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1636968456
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_27
timestamp 1636968456
transform 1 0 3588 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_39
timestamp 1636968456
transform 1 0 4692 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_51
timestamp 1
transform 1 0 5796 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_57
timestamp 1636968456
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_69
timestamp 1636968456
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_81
timestamp 1636968456
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_93
timestamp 1636968456
transform 1 0 9660 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_105
timestamp 1
transform 1 0 10764 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_111
timestamp 1
transform 1 0 11316 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_113
timestamp 1636968456
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_125
timestamp 1636968456
transform 1 0 12604 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_137
timestamp 1636968456
transform 1 0 13708 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_149
timestamp 1636968456
transform 1 0 14812 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_161
timestamp 1
transform 1 0 15916 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_167
timestamp 1
transform 1 0 16468 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_169
timestamp 1636968456
transform 1 0 16652 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_181
timestamp 1636968456
transform 1 0 17756 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_193
timestamp 1636968456
transform 1 0 18860 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_205
timestamp 1636968456
transform 1 0 19964 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_217
timestamp 1
transform 1 0 21068 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_223
timestamp 1
transform 1 0 21620 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_225
timestamp 1636968456
transform 1 0 21804 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_237
timestamp 1636968456
transform 1 0 22908 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_249
timestamp 1636968456
transform 1 0 24012 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_261
timestamp 1636968456
transform 1 0 25116 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_273
timestamp 1
transform 1 0 26220 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_279
timestamp 1
transform 1 0 26772 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_281
timestamp 1636968456
transform 1 0 26956 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_293
timestamp 1636968456
transform 1 0 28060 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_305
timestamp 1636968456
transform 1 0 29164 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_317
timestamp 1636968456
transform 1 0 30268 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_329
timestamp 1
transform 1 0 31372 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_335
timestamp 1
transform 1 0 31924 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_337
timestamp 1636968456
transform 1 0 32108 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_349
timestamp 1636968456
transform 1 0 33212 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_361
timestamp 1636968456
transform 1 0 34316 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_373
timestamp 1636968456
transform 1 0 35420 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_385
timestamp 1
transform 1 0 36524 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_391
timestamp 1
transform 1 0 37076 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_393
timestamp 1636968456
transform 1 0 37260 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_405
timestamp 1636968456
transform 1 0 38364 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_417
timestamp 1636968456
transform 1 0 39468 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_429
timestamp 1636968456
transform 1 0 40572 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_441
timestamp 1
transform 1 0 41676 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_447
timestamp 1
transform 1 0 42228 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_449
timestamp 1636968456
transform 1 0 42412 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_461
timestamp 1636968456
transform 1 0 43516 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_473
timestamp 1636968456
transform 1 0 44620 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_485
timestamp 1636968456
transform 1 0 45724 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_497
timestamp 1
transform 1 0 46828 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_503
timestamp 1
transform 1 0 47380 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_505
timestamp 1636968456
transform 1 0 47564 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_517
timestamp 1636968456
transform 1 0 48668 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_529
timestamp 1636968456
transform 1 0 49772 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_541
timestamp 1636968456
transform 1 0 50876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_553
timestamp 1
transform 1 0 51980 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_559
timestamp 1
transform 1 0 52532 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_561
timestamp 1636968456
transform 1 0 52716 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_573
timestamp 1636968456
transform 1 0 53820 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_585
timestamp 1636968456
transform 1 0 54924 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_597
timestamp 1636968456
transform 1 0 56028 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_609
timestamp 1
transform 1 0 57132 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_615
timestamp 1
transform 1 0 57684 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_617
timestamp 1636968456
transform 1 0 57868 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_629
timestamp 1636968456
transform 1 0 58972 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_641
timestamp 1636968456
transform 1 0 60076 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_653
timestamp 1636968456
transform 1 0 61180 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_665
timestamp 1
transform 1 0 62284 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_671
timestamp 1
transform 1 0 62836 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_673
timestamp 1636968456
transform 1 0 63020 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_685
timestamp 1636968456
transform 1 0 64124 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_697
timestamp 1636968456
transform 1 0 65228 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_709
timestamp 1636968456
transform 1 0 66332 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_721
timestamp 1
transform 1 0 67436 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_727
timestamp 1
transform 1 0 67988 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_729
timestamp 1636968456
transform 1 0 68172 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_741
timestamp 1636968456
transform 1 0 69276 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_753
timestamp 1636968456
transform 1 0 70380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_765
timestamp 1636968456
transform 1 0 71484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_777
timestamp 1
transform 1 0 72588 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_783
timestamp 1
transform 1 0 73140 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_785
timestamp 1636968456
transform 1 0 73324 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_797
timestamp 1636968456
transform 1 0 74428 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_809
timestamp 1636968456
transform 1 0 75532 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_821
timestamp 1636968456
transform 1 0 76636 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_833
timestamp 1
transform 1 0 77740 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_839
timestamp 1
transform 1 0 78292 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_841
timestamp 1636968456
transform 1 0 78476 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_853
timestamp 1636968456
transform 1 0 79580 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_865
timestamp 1636968456
transform 1 0 80684 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_877
timestamp 1636968456
transform 1 0 81788 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_889
timestamp 1
transform 1 0 82892 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_895
timestamp 1
transform 1 0 83444 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_897
timestamp 1636968456
transform 1 0 83628 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_909
timestamp 1636968456
transform 1 0 84732 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_921
timestamp 1636968456
transform 1 0 85836 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_933
timestamp 1636968456
transform 1 0 86940 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_945
timestamp 1
transform 1 0 88044 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_951
timestamp 1
transform 1 0 88596 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_123_953
timestamp 1
transform 1 0 88780 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_958
timestamp 1636968456
transform 1 0 89240 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_970
timestamp 1636968456
transform 1 0 90344 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_982
timestamp 1636968456
transform 1 0 91448 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_994
timestamp 1636968456
transform 1 0 92552 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_1006
timestamp 1
transform 1 0 93656 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1009
timestamp 1636968456
transform 1 0 93932 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1021
timestamp 1636968456
transform 1 0 95036 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1033
timestamp 1636968456
transform 1 0 96140 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1045
timestamp 1636968456
transform 1 0 97244 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_1057
timestamp 1
transform 1 0 98348 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1063
timestamp 1
transform 1 0 98900 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1065
timestamp 1636968456
transform 1 0 99084 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1077
timestamp 1636968456
transform 1 0 100188 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1089
timestamp 1636968456
transform 1 0 101292 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1101
timestamp 1636968456
transform 1 0 102396 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_1113
timestamp 1
transform 1 0 103500 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1119
timestamp 1
transform 1 0 104052 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1121
timestamp 1636968456
transform 1 0 104236 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1133
timestamp 1636968456
transform 1 0 105340 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1145
timestamp 1636968456
transform 1 0 106444 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_1157
timestamp 1
transform 1 0 107548 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_123_1165
timestamp 1
transform 1 0 108284 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_124_3
timestamp 1636968456
transform 1 0 1380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_15
timestamp 1636968456
transform 1 0 2484 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 1
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_29
timestamp 1636968456
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_41
timestamp 1636968456
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_53
timestamp 1636968456
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_65
timestamp 1636968456
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_85
timestamp 1636968456
transform 1 0 8924 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_97
timestamp 1636968456
transform 1 0 10028 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_109
timestamp 1636968456
transform 1 0 11132 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_121
timestamp 1636968456
transform 1 0 12236 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_133
timestamp 1
transform 1 0 13340 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_139
timestamp 1
transform 1 0 13892 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_141
timestamp 1636968456
transform 1 0 14076 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_153
timestamp 1636968456
transform 1 0 15180 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_165
timestamp 1636968456
transform 1 0 16284 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_177
timestamp 1636968456
transform 1 0 17388 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_189
timestamp 1
transform 1 0 18492 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_195
timestamp 1
transform 1 0 19044 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_197
timestamp 1636968456
transform 1 0 19228 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_209
timestamp 1636968456
transform 1 0 20332 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_221
timestamp 1636968456
transform 1 0 21436 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_233
timestamp 1636968456
transform 1 0 22540 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_245
timestamp 1
transform 1 0 23644 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_251
timestamp 1
transform 1 0 24196 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_253
timestamp 1636968456
transform 1 0 24380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_265
timestamp 1636968456
transform 1 0 25484 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_277
timestamp 1636968456
transform 1 0 26588 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_289
timestamp 1636968456
transform 1 0 27692 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_301
timestamp 1
transform 1 0 28796 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_307
timestamp 1
transform 1 0 29348 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_309
timestamp 1636968456
transform 1 0 29532 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_321
timestamp 1636968456
transform 1 0 30636 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_333
timestamp 1636968456
transform 1 0 31740 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_345
timestamp 1636968456
transform 1 0 32844 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_357
timestamp 1
transform 1 0 33948 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_363
timestamp 1
transform 1 0 34500 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_365
timestamp 1636968456
transform 1 0 34684 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_377
timestamp 1636968456
transform 1 0 35788 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_389
timestamp 1636968456
transform 1 0 36892 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_401
timestamp 1636968456
transform 1 0 37996 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_413
timestamp 1
transform 1 0 39100 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_419
timestamp 1
transform 1 0 39652 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_421
timestamp 1636968456
transform 1 0 39836 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_433
timestamp 1636968456
transform 1 0 40940 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_445
timestamp 1636968456
transform 1 0 42044 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_457
timestamp 1636968456
transform 1 0 43148 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_469
timestamp 1
transform 1 0 44252 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_475
timestamp 1
transform 1 0 44804 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_477
timestamp 1636968456
transform 1 0 44988 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_489
timestamp 1636968456
transform 1 0 46092 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_501
timestamp 1636968456
transform 1 0 47196 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_513
timestamp 1636968456
transform 1 0 48300 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_525
timestamp 1
transform 1 0 49404 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_531
timestamp 1
transform 1 0 49956 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_533
timestamp 1636968456
transform 1 0 50140 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_545
timestamp 1636968456
transform 1 0 51244 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_557
timestamp 1636968456
transform 1 0 52348 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_569
timestamp 1636968456
transform 1 0 53452 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_581
timestamp 1
transform 1 0 54556 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_587
timestamp 1
transform 1 0 55108 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_589
timestamp 1636968456
transform 1 0 55292 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_601
timestamp 1636968456
transform 1 0 56396 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_613
timestamp 1636968456
transform 1 0 57500 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_625
timestamp 1636968456
transform 1 0 58604 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_637
timestamp 1
transform 1 0 59708 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_643
timestamp 1
transform 1 0 60260 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_645
timestamp 1636968456
transform 1 0 60444 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_657
timestamp 1636968456
transform 1 0 61548 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_669
timestamp 1636968456
transform 1 0 62652 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_681
timestamp 1636968456
transform 1 0 63756 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_693
timestamp 1
transform 1 0 64860 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_699
timestamp 1
transform 1 0 65412 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_701
timestamp 1636968456
transform 1 0 65596 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_713
timestamp 1636968456
transform 1 0 66700 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_725
timestamp 1636968456
transform 1 0 67804 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_737
timestamp 1636968456
transform 1 0 68908 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_749
timestamp 1
transform 1 0 70012 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_755
timestamp 1
transform 1 0 70564 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_757
timestamp 1636968456
transform 1 0 70748 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_769
timestamp 1636968456
transform 1 0 71852 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_781
timestamp 1636968456
transform 1 0 72956 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_793
timestamp 1636968456
transform 1 0 74060 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_805
timestamp 1
transform 1 0 75164 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_811
timestamp 1
transform 1 0 75716 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_813
timestamp 1636968456
transform 1 0 75900 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_825
timestamp 1636968456
transform 1 0 77004 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_837
timestamp 1636968456
transform 1 0 78108 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_849
timestamp 1636968456
transform 1 0 79212 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_861
timestamp 1
transform 1 0 80316 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_867
timestamp 1
transform 1 0 80868 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_869
timestamp 1636968456
transform 1 0 81052 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_881
timestamp 1636968456
transform 1 0 82156 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_893
timestamp 1636968456
transform 1 0 83260 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_905
timestamp 1636968456
transform 1 0 84364 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_917
timestamp 1
transform 1 0 85468 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_923
timestamp 1
transform 1 0 86020 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_925
timestamp 1636968456
transform 1 0 86204 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_937
timestamp 1636968456
transform 1 0 87308 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_949
timestamp 1636968456
transform 1 0 88412 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_961
timestamp 1636968456
transform 1 0 89516 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_973
timestamp 1
transform 1 0 90620 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_979
timestamp 1
transform 1 0 91172 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_981
timestamp 1636968456
transform 1 0 91356 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_993
timestamp 1636968456
transform 1 0 92460 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1005
timestamp 1636968456
transform 1 0 93564 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1017
timestamp 1636968456
transform 1 0 94668 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1029
timestamp 1
transform 1 0 95772 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1035
timestamp 1
transform 1 0 96324 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1037
timestamp 1636968456
transform 1 0 96508 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1049
timestamp 1636968456
transform 1 0 97612 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1061
timestamp 1636968456
transform 1 0 98716 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1073
timestamp 1636968456
transform 1 0 99820 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1085
timestamp 1
transform 1 0 100924 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1091
timestamp 1
transform 1 0 101476 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1093
timestamp 1636968456
transform 1 0 101660 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1105
timestamp 1636968456
transform 1 0 102764 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1117
timestamp 1636968456
transform 1 0 103868 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1129
timestamp 1636968456
transform 1 0 104972 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1141
timestamp 1
transform 1 0 106076 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1147
timestamp 1
transform 1 0 106628 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1149
timestamp 1636968456
transform 1 0 106812 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1161
timestamp 1
transform 1 0 107916 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1167
timestamp 1
transform 1 0 108468 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_3
timestamp 1636968456
transform 1 0 1380 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_15
timestamp 1636968456
transform 1 0 2484 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_27
timestamp 1636968456
transform 1 0 3588 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_39
timestamp 1636968456
transform 1 0 4692 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_51
timestamp 1
transform 1 0 5796 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_57
timestamp 1636968456
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_69
timestamp 1636968456
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_81
timestamp 1636968456
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_93
timestamp 1636968456
transform 1 0 9660 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_105
timestamp 1
transform 1 0 10764 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_111
timestamp 1
transform 1 0 11316 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_113
timestamp 1636968456
transform 1 0 11500 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_125
timestamp 1636968456
transform 1 0 12604 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_137
timestamp 1636968456
transform 1 0 13708 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_149
timestamp 1636968456
transform 1 0 14812 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_161
timestamp 1
transform 1 0 15916 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_167
timestamp 1
transform 1 0 16468 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_169
timestamp 1636968456
transform 1 0 16652 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_181
timestamp 1636968456
transform 1 0 17756 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_193
timestamp 1636968456
transform 1 0 18860 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_205
timestamp 1636968456
transform 1 0 19964 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_217
timestamp 1
transform 1 0 21068 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_223
timestamp 1
transform 1 0 21620 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_225
timestamp 1636968456
transform 1 0 21804 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_237
timestamp 1636968456
transform 1 0 22908 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_249
timestamp 1636968456
transform 1 0 24012 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_261
timestamp 1636968456
transform 1 0 25116 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_273
timestamp 1
transform 1 0 26220 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_279
timestamp 1
transform 1 0 26772 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_281
timestamp 1636968456
transform 1 0 26956 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_293
timestamp 1636968456
transform 1 0 28060 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_305
timestamp 1636968456
transform 1 0 29164 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_317
timestamp 1636968456
transform 1 0 30268 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_329
timestamp 1
transform 1 0 31372 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_335
timestamp 1
transform 1 0 31924 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_337
timestamp 1636968456
transform 1 0 32108 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_349
timestamp 1636968456
transform 1 0 33212 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_361
timestamp 1636968456
transform 1 0 34316 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_373
timestamp 1636968456
transform 1 0 35420 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_385
timestamp 1
transform 1 0 36524 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_391
timestamp 1
transform 1 0 37076 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_393
timestamp 1636968456
transform 1 0 37260 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_405
timestamp 1636968456
transform 1 0 38364 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_417
timestamp 1636968456
transform 1 0 39468 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_429
timestamp 1636968456
transform 1 0 40572 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_441
timestamp 1
transform 1 0 41676 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_447
timestamp 1
transform 1 0 42228 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_449
timestamp 1636968456
transform 1 0 42412 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_461
timestamp 1636968456
transform 1 0 43516 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_473
timestamp 1636968456
transform 1 0 44620 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_485
timestamp 1636968456
transform 1 0 45724 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_497
timestamp 1
transform 1 0 46828 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_503
timestamp 1
transform 1 0 47380 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_505
timestamp 1636968456
transform 1 0 47564 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_517
timestamp 1636968456
transform 1 0 48668 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_529
timestamp 1636968456
transform 1 0 49772 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_541
timestamp 1636968456
transform 1 0 50876 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_553
timestamp 1
transform 1 0 51980 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_559
timestamp 1
transform 1 0 52532 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_561
timestamp 1636968456
transform 1 0 52716 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_573
timestamp 1636968456
transform 1 0 53820 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_585
timestamp 1636968456
transform 1 0 54924 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_597
timestamp 1636968456
transform 1 0 56028 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_609
timestamp 1
transform 1 0 57132 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_615
timestamp 1
transform 1 0 57684 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_617
timestamp 1636968456
transform 1 0 57868 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_629
timestamp 1636968456
transform 1 0 58972 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_641
timestamp 1636968456
transform 1 0 60076 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_653
timestamp 1636968456
transform 1 0 61180 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_665
timestamp 1
transform 1 0 62284 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_671
timestamp 1
transform 1 0 62836 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_673
timestamp 1636968456
transform 1 0 63020 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_685
timestamp 1636968456
transform 1 0 64124 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_697
timestamp 1636968456
transform 1 0 65228 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_709
timestamp 1636968456
transform 1 0 66332 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_721
timestamp 1
transform 1 0 67436 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_727
timestamp 1
transform 1 0 67988 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_729
timestamp 1636968456
transform 1 0 68172 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_741
timestamp 1636968456
transform 1 0 69276 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_753
timestamp 1636968456
transform 1 0 70380 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_765
timestamp 1636968456
transform 1 0 71484 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_777
timestamp 1
transform 1 0 72588 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_783
timestamp 1
transform 1 0 73140 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_785
timestamp 1636968456
transform 1 0 73324 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_797
timestamp 1636968456
transform 1 0 74428 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_809
timestamp 1636968456
transform 1 0 75532 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_821
timestamp 1
transform 1 0 76636 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_125_838
timestamp 1
transform 1 0 78200 0 -1 70720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_125_841
timestamp 1636968456
transform 1 0 78476 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_853
timestamp 1636968456
transform 1 0 79580 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_865
timestamp 1636968456
transform 1 0 80684 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_877
timestamp 1636968456
transform 1 0 81788 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_889
timestamp 1
transform 1 0 82892 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_895
timestamp 1
transform 1 0 83444 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_897
timestamp 1636968456
transform 1 0 83628 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_909
timestamp 1636968456
transform 1 0 84732 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_921
timestamp 1636968456
transform 1 0 85836 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_933
timestamp 1636968456
transform 1 0 86940 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_945
timestamp 1
transform 1 0 88044 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_951
timestamp 1
transform 1 0 88596 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_953
timestamp 1636968456
transform 1 0 88780 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_965
timestamp 1636968456
transform 1 0 89884 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_977
timestamp 1636968456
transform 1 0 90988 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_989
timestamp 1636968456
transform 1 0 92092 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1001
timestamp 1
transform 1 0 93196 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1007
timestamp 1
transform 1 0 93748 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1009
timestamp 1636968456
transform 1 0 93932 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1021
timestamp 1636968456
transform 1 0 95036 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1033
timestamp 1636968456
transform 1 0 96140 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1045
timestamp 1636968456
transform 1 0 97244 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1057
timestamp 1
transform 1 0 98348 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1063
timestamp 1
transform 1 0 98900 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1065
timestamp 1636968456
transform 1 0 99084 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1077
timestamp 1636968456
transform 1 0 100188 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1089
timestamp 1636968456
transform 1 0 101292 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1101
timestamp 1636968456
transform 1 0 102396 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1113
timestamp 1
transform 1 0 103500 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1119
timestamp 1
transform 1 0 104052 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1121
timestamp 1636968456
transform 1 0 104236 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1133
timestamp 1636968456
transform 1 0 105340 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1145
timestamp 1636968456
transform 1 0 106444 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_1157
timestamp 1
transform 1 0 107548 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_125_1165
timestamp 1
transform 1 0 108284 0 -1 70720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_126_3
timestamp 1636968456
transform 1 0 1380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_15
timestamp 1636968456
transform 1 0 2484 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 1
transform 1 0 3588 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_29
timestamp 1636968456
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_41
timestamp 1636968456
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_53
timestamp 1636968456
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_65
timestamp 1636968456
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_85
timestamp 1636968456
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_97
timestamp 1636968456
transform 1 0 10028 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_109
timestamp 1636968456
transform 1 0 11132 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_121
timestamp 1636968456
transform 1 0 12236 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_133
timestamp 1
transform 1 0 13340 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_139
timestamp 1
transform 1 0 13892 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_141
timestamp 1636968456
transform 1 0 14076 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_153
timestamp 1636968456
transform 1 0 15180 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_165
timestamp 1636968456
transform 1 0 16284 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_177
timestamp 1636968456
transform 1 0 17388 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_189
timestamp 1
transform 1 0 18492 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_195
timestamp 1
transform 1 0 19044 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_197
timestamp 1636968456
transform 1 0 19228 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_209
timestamp 1636968456
transform 1 0 20332 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_221
timestamp 1636968456
transform 1 0 21436 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_233
timestamp 1636968456
transform 1 0 22540 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_245
timestamp 1
transform 1 0 23644 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_251
timestamp 1
transform 1 0 24196 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_253
timestamp 1636968456
transform 1 0 24380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_265
timestamp 1636968456
transform 1 0 25484 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_277
timestamp 1636968456
transform 1 0 26588 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_289
timestamp 1636968456
transform 1 0 27692 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_301
timestamp 1
transform 1 0 28796 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_307
timestamp 1
transform 1 0 29348 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_309
timestamp 1636968456
transform 1 0 29532 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_321
timestamp 1636968456
transform 1 0 30636 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_333
timestamp 1636968456
transform 1 0 31740 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_345
timestamp 1636968456
transform 1 0 32844 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_357
timestamp 1
transform 1 0 33948 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_363
timestamp 1
transform 1 0 34500 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_365
timestamp 1636968456
transform 1 0 34684 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_377
timestamp 1636968456
transform 1 0 35788 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_389
timestamp 1636968456
transform 1 0 36892 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_401
timestamp 1636968456
transform 1 0 37996 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_413
timestamp 1
transform 1 0 39100 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_419
timestamp 1
transform 1 0 39652 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_421
timestamp 1636968456
transform 1 0 39836 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_433
timestamp 1636968456
transform 1 0 40940 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_445
timestamp 1636968456
transform 1 0 42044 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_457
timestamp 1636968456
transform 1 0 43148 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_469
timestamp 1
transform 1 0 44252 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_475
timestamp 1
transform 1 0 44804 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_477
timestamp 1636968456
transform 1 0 44988 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_489
timestamp 1636968456
transform 1 0 46092 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_501
timestamp 1636968456
transform 1 0 47196 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_513
timestamp 1636968456
transform 1 0 48300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_525
timestamp 1
transform 1 0 49404 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_531
timestamp 1
transform 1 0 49956 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_533
timestamp 1636968456
transform 1 0 50140 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_545
timestamp 1636968456
transform 1 0 51244 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_557
timestamp 1636968456
transform 1 0 52348 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_569
timestamp 1636968456
transform 1 0 53452 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_581
timestamp 1
transform 1 0 54556 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_587
timestamp 1
transform 1 0 55108 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_589
timestamp 1636968456
transform 1 0 55292 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_601
timestamp 1636968456
transform 1 0 56396 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_613
timestamp 1636968456
transform 1 0 57500 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_625
timestamp 1636968456
transform 1 0 58604 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_637
timestamp 1
transform 1 0 59708 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_643
timestamp 1
transform 1 0 60260 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_645
timestamp 1636968456
transform 1 0 60444 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_657
timestamp 1636968456
transform 1 0 61548 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_669
timestamp 1636968456
transform 1 0 62652 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_681
timestamp 1636968456
transform 1 0 63756 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_693
timestamp 1
transform 1 0 64860 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_699
timestamp 1
transform 1 0 65412 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_701
timestamp 1636968456
transform 1 0 65596 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_713
timestamp 1636968456
transform 1 0 66700 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_725
timestamp 1636968456
transform 1 0 67804 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_737
timestamp 1636968456
transform 1 0 68908 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_749
timestamp 1
transform 1 0 70012 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_755
timestamp 1
transform 1 0 70564 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_757
timestamp 1636968456
transform 1 0 70748 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_769
timestamp 1636968456
transform 1 0 71852 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_781
timestamp 1636968456
transform 1 0 72956 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_793
timestamp 1636968456
transform 1 0 74060 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_805
timestamp 1
transform 1 0 75164 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_811
timestamp 1
transform 1 0 75716 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_813
timestamp 1636968456
transform 1 0 75900 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_825
timestamp 1
transform 1 0 77004 0 1 70720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_126_839
timestamp 1636968456
transform 1 0 78292 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_851
timestamp 1636968456
transform 1 0 79396 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_863
timestamp 1
transform 1 0 80500 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_126_867
timestamp 1
transform 1 0 80868 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_869
timestamp 1636968456
transform 1 0 81052 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_881
timestamp 1636968456
transform 1 0 82156 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_893
timestamp 1636968456
transform 1 0 83260 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_905
timestamp 1636968456
transform 1 0 84364 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_917
timestamp 1
transform 1 0 85468 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_923
timestamp 1
transform 1 0 86020 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_925
timestamp 1636968456
transform 1 0 86204 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_937
timestamp 1
transform 1 0 87308 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_126_946
timestamp 1
transform 1 0 88136 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_126_974
timestamp 1
transform 1 0 90712 0 1 70720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_126_981
timestamp 1636968456
transform 1 0 91356 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_993
timestamp 1636968456
transform 1 0 92460 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1005
timestamp 1636968456
transform 1 0 93564 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1017
timestamp 1636968456
transform 1 0 94668 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_1029
timestamp 1
transform 1 0 95772 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1035
timestamp 1
transform 1 0 96324 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1037
timestamp 1636968456
transform 1 0 96508 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1049
timestamp 1636968456
transform 1 0 97612 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1061
timestamp 1636968456
transform 1 0 98716 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1073
timestamp 1636968456
transform 1 0 99820 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_1085
timestamp 1
transform 1 0 100924 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1091
timestamp 1
transform 1 0 101476 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1093
timestamp 1636968456
transform 1 0 101660 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1105
timestamp 1636968456
transform 1 0 102764 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1117
timestamp 1636968456
transform 1 0 103868 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1129
timestamp 1636968456
transform 1 0 104972 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_1141
timestamp 1
transform 1 0 106076 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1147
timestamp 1
transform 1 0 106628 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1149
timestamp 1636968456
transform 1 0 106812 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_1161
timestamp 1
transform 1 0 107916 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1167
timestamp 1
transform 1 0 108468 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_3
timestamp 1636968456
transform 1 0 1380 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_15
timestamp 1636968456
transform 1 0 2484 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_27
timestamp 1636968456
transform 1 0 3588 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_39
timestamp 1636968456
transform 1 0 4692 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_51
timestamp 1
transform 1 0 5796 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_57
timestamp 1636968456
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_69
timestamp 1636968456
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_81
timestamp 1636968456
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_93
timestamp 1636968456
transform 1 0 9660 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_105
timestamp 1
transform 1 0 10764 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_111
timestamp 1
transform 1 0 11316 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_113
timestamp 1636968456
transform 1 0 11500 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_125
timestamp 1636968456
transform 1 0 12604 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_137
timestamp 1636968456
transform 1 0 13708 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_149
timestamp 1636968456
transform 1 0 14812 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_161
timestamp 1
transform 1 0 15916 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_167
timestamp 1
transform 1 0 16468 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_169
timestamp 1636968456
transform 1 0 16652 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_181
timestamp 1636968456
transform 1 0 17756 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_193
timestamp 1636968456
transform 1 0 18860 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_205
timestamp 1636968456
transform 1 0 19964 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_217
timestamp 1
transform 1 0 21068 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_223
timestamp 1
transform 1 0 21620 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_225
timestamp 1636968456
transform 1 0 21804 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_237
timestamp 1636968456
transform 1 0 22908 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_249
timestamp 1636968456
transform 1 0 24012 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_261
timestamp 1636968456
transform 1 0 25116 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_273
timestamp 1
transform 1 0 26220 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_279
timestamp 1
transform 1 0 26772 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_281
timestamp 1636968456
transform 1 0 26956 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_293
timestamp 1636968456
transform 1 0 28060 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_305
timestamp 1636968456
transform 1 0 29164 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_317
timestamp 1636968456
transform 1 0 30268 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_329
timestamp 1
transform 1 0 31372 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_335
timestamp 1
transform 1 0 31924 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_337
timestamp 1636968456
transform 1 0 32108 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_349
timestamp 1636968456
transform 1 0 33212 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_361
timestamp 1636968456
transform 1 0 34316 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_373
timestamp 1636968456
transform 1 0 35420 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_385
timestamp 1
transform 1 0 36524 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_391
timestamp 1
transform 1 0 37076 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_393
timestamp 1636968456
transform 1 0 37260 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_405
timestamp 1636968456
transform 1 0 38364 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_417
timestamp 1636968456
transform 1 0 39468 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_429
timestamp 1636968456
transform 1 0 40572 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_441
timestamp 1
transform 1 0 41676 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_447
timestamp 1
transform 1 0 42228 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_449
timestamp 1636968456
transform 1 0 42412 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_461
timestamp 1636968456
transform 1 0 43516 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_473
timestamp 1636968456
transform 1 0 44620 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_485
timestamp 1636968456
transform 1 0 45724 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_497
timestamp 1
transform 1 0 46828 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_503
timestamp 1
transform 1 0 47380 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_505
timestamp 1636968456
transform 1 0 47564 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_517
timestamp 1636968456
transform 1 0 48668 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_529
timestamp 1636968456
transform 1 0 49772 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_541
timestamp 1636968456
transform 1 0 50876 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_553
timestamp 1
transform 1 0 51980 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_559
timestamp 1
transform 1 0 52532 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_561
timestamp 1636968456
transform 1 0 52716 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_573
timestamp 1636968456
transform 1 0 53820 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_585
timestamp 1636968456
transform 1 0 54924 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_597
timestamp 1636968456
transform 1 0 56028 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_609
timestamp 1
transform 1 0 57132 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_615
timestamp 1
transform 1 0 57684 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_617
timestamp 1636968456
transform 1 0 57868 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_629
timestamp 1636968456
transform 1 0 58972 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_641
timestamp 1636968456
transform 1 0 60076 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_653
timestamp 1636968456
transform 1 0 61180 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_665
timestamp 1
transform 1 0 62284 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_671
timestamp 1
transform 1 0 62836 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_673
timestamp 1636968456
transform 1 0 63020 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_685
timestamp 1636968456
transform 1 0 64124 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_697
timestamp 1636968456
transform 1 0 65228 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_709
timestamp 1636968456
transform 1 0 66332 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_721
timestamp 1
transform 1 0 67436 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_727
timestamp 1
transform 1 0 67988 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_729
timestamp 1636968456
transform 1 0 68172 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_741
timestamp 1636968456
transform 1 0 69276 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_753
timestamp 1636968456
transform 1 0 70380 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_765
timestamp 1636968456
transform 1 0 71484 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_777
timestamp 1
transform 1 0 72588 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_783
timestamp 1
transform 1 0 73140 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_785
timestamp 1636968456
transform 1 0 73324 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_797
timestamp 1636968456
transform 1 0 74428 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_809
timestamp 1636968456
transform 1 0 75532 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_821
timestamp 1636968456
transform 1 0 76636 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_833
timestamp 1
transform 1 0 77740 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_839
timestamp 1
transform 1 0 78292 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_841
timestamp 1636968456
transform 1 0 78476 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_853
timestamp 1636968456
transform 1 0 79580 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_865
timestamp 1636968456
transform 1 0 80684 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_877
timestamp 1636968456
transform 1 0 81788 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_889
timestamp 1
transform 1 0 82892 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_895
timestamp 1
transform 1 0 83444 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_897
timestamp 1636968456
transform 1 0 83628 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_909
timestamp 1636968456
transform 1 0 84732 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_921
timestamp 1636968456
transform 1 0 85836 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_933
timestamp 1636968456
transform 1 0 86940 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_945
timestamp 1
transform 1 0 88044 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_951
timestamp 1
transform 1 0 88596 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_953
timestamp 1636968456
transform 1 0 88780 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_965
timestamp 1
transform 1 0 89884 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_973
timestamp 1
transform 1 0 90620 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_127_977
timestamp 1
transform 1 0 90988 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_985
timestamp 1
transform 1 0 91724 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_992
timestamp 1636968456
transform 1 0 92368 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_1004
timestamp 1
transform 1 0 93472 0 -1 71808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1009
timestamp 1636968456
transform 1 0 93932 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1021
timestamp 1636968456
transform 1 0 95036 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1033
timestamp 1636968456
transform 1 0 96140 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1045
timestamp 1636968456
transform 1 0 97244 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_1057
timestamp 1
transform 1 0 98348 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1063
timestamp 1
transform 1 0 98900 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1065
timestamp 1636968456
transform 1 0 99084 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1077
timestamp 1636968456
transform 1 0 100188 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1089
timestamp 1636968456
transform 1 0 101292 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1101
timestamp 1636968456
transform 1 0 102396 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_1113
timestamp 1
transform 1 0 103500 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1119
timestamp 1
transform 1 0 104052 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1121
timestamp 1636968456
transform 1 0 104236 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1133
timestamp 1636968456
transform 1 0 105340 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1145
timestamp 1636968456
transform 1 0 106444 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_1157
timestamp 1
transform 1 0 107548 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_127_1165
timestamp 1
transform 1 0 108284 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_128_3
timestamp 1636968456
transform 1 0 1380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_15
timestamp 1636968456
transform 1 0 2484 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 1
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_29
timestamp 1636968456
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_41
timestamp 1636968456
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_53
timestamp 1636968456
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_65
timestamp 1636968456
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_85
timestamp 1636968456
transform 1 0 8924 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_97
timestamp 1636968456
transform 1 0 10028 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_109
timestamp 1636968456
transform 1 0 11132 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_121
timestamp 1636968456
transform 1 0 12236 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_133
timestamp 1
transform 1 0 13340 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_139
timestamp 1
transform 1 0 13892 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_141
timestamp 1636968456
transform 1 0 14076 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_153
timestamp 1636968456
transform 1 0 15180 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_165
timestamp 1636968456
transform 1 0 16284 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_177
timestamp 1636968456
transform 1 0 17388 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_189
timestamp 1
transform 1 0 18492 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_195
timestamp 1
transform 1 0 19044 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_197
timestamp 1636968456
transform 1 0 19228 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_209
timestamp 1636968456
transform 1 0 20332 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_221
timestamp 1636968456
transform 1 0 21436 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_233
timestamp 1636968456
transform 1 0 22540 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_245
timestamp 1
transform 1 0 23644 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_251
timestamp 1
transform 1 0 24196 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_253
timestamp 1636968456
transform 1 0 24380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_265
timestamp 1636968456
transform 1 0 25484 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_277
timestamp 1636968456
transform 1 0 26588 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_289
timestamp 1636968456
transform 1 0 27692 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_301
timestamp 1
transform 1 0 28796 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_307
timestamp 1
transform 1 0 29348 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_309
timestamp 1636968456
transform 1 0 29532 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_321
timestamp 1636968456
transform 1 0 30636 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_333
timestamp 1636968456
transform 1 0 31740 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_345
timestamp 1636968456
transform 1 0 32844 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_357
timestamp 1
transform 1 0 33948 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_363
timestamp 1
transform 1 0 34500 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_365
timestamp 1636968456
transform 1 0 34684 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_377
timestamp 1636968456
transform 1 0 35788 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_389
timestamp 1636968456
transform 1 0 36892 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_401
timestamp 1636968456
transform 1 0 37996 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_413
timestamp 1
transform 1 0 39100 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_419
timestamp 1
transform 1 0 39652 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_421
timestamp 1636968456
transform 1 0 39836 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_433
timestamp 1636968456
transform 1 0 40940 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_445
timestamp 1636968456
transform 1 0 42044 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_457
timestamp 1636968456
transform 1 0 43148 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_128_469
timestamp 1
transform 1 0 44252 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_128_475
timestamp 1
transform 1 0 44804 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_477
timestamp 1636968456
transform 1 0 44988 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_489
timestamp 1636968456
transform 1 0 46092 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_501
timestamp 1636968456
transform 1 0 47196 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_513
timestamp 1636968456
transform 1 0 48300 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_525
timestamp 1
transform 1 0 49404 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_531
timestamp 1
transform 1 0 49956 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_533
timestamp 1636968456
transform 1 0 50140 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_545
timestamp 1636968456
transform 1 0 51244 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_557
timestamp 1636968456
transform 1 0 52348 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_569
timestamp 1636968456
transform 1 0 53452 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_581
timestamp 1
transform 1 0 54556 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_587
timestamp 1
transform 1 0 55108 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_128_589
timestamp 1
transform 1 0 55292 0 1 71808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_128_619
timestamp 1636968456
transform 1 0 58052 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_631
timestamp 1636968456
transform 1 0 59156 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_643
timestamp 1
transform 1 0 60260 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_645
timestamp 1636968456
transform 1 0 60444 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_657
timestamp 1636968456
transform 1 0 61548 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_669
timestamp 1636968456
transform 1 0 62652 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_681
timestamp 1636968456
transform 1 0 63756 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_693
timestamp 1
transform 1 0 64860 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_699
timestamp 1
transform 1 0 65412 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_701
timestamp 1636968456
transform 1 0 65596 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_713
timestamp 1636968456
transform 1 0 66700 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_725
timestamp 1636968456
transform 1 0 67804 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_737
timestamp 1636968456
transform 1 0 68908 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_749
timestamp 1
transform 1 0 70012 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_755
timestamp 1
transform 1 0 70564 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_757
timestamp 1636968456
transform 1 0 70748 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_769
timestamp 1636968456
transform 1 0 71852 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_781
timestamp 1636968456
transform 1 0 72956 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_798
timestamp 1636968456
transform 1 0 74520 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_128_810
timestamp 1
transform 1 0 75624 0 1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_128_813
timestamp 1636968456
transform 1 0 75900 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_825
timestamp 1636968456
transform 1 0 77004 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_837
timestamp 1636968456
transform 1 0 78108 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_849
timestamp 1636968456
transform 1 0 79212 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_861
timestamp 1
transform 1 0 80316 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_867
timestamp 1
transform 1 0 80868 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_869
timestamp 1636968456
transform 1 0 81052 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_881
timestamp 1636968456
transform 1 0 82156 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_893
timestamp 1636968456
transform 1 0 83260 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_905
timestamp 1636968456
transform 1 0 84364 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_917
timestamp 1
transform 1 0 85468 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_923
timestamp 1
transform 1 0 86020 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_925
timestamp 1636968456
transform 1 0 86204 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_937
timestamp 1636968456
transform 1 0 87308 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_949
timestamp 1636968456
transform 1 0 88412 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_961
timestamp 1
transform 1 0 89516 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_128_969
timestamp 1
transform 1 0 90252 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_128_975
timestamp 1
transform 1 0 90804 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_128_979
timestamp 1
transform 1 0 91172 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_128_981
timestamp 1
transform 1 0 91356 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_128_991
timestamp 1
transform 1 0 92276 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_998
timestamp 1636968456
transform 1 0 92920 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1010
timestamp 1636968456
transform 1 0 94024 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1022
timestamp 1636968456
transform 1 0 95128 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_128_1034
timestamp 1
transform 1 0 96232 0 1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1037
timestamp 1636968456
transform 1 0 96508 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1049
timestamp 1636968456
transform 1 0 97612 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1061
timestamp 1636968456
transform 1 0 98716 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1073
timestamp 1636968456
transform 1 0 99820 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_1085
timestamp 1
transform 1 0 100924 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1091
timestamp 1
transform 1 0 101476 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1093
timestamp 1636968456
transform 1 0 101660 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1105
timestamp 1636968456
transform 1 0 102764 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1117
timestamp 1636968456
transform 1 0 103868 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1129
timestamp 1636968456
transform 1 0 104972 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_1141
timestamp 1
transform 1 0 106076 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1147
timestamp 1
transform 1 0 106628 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1149
timestamp 1636968456
transform 1 0 106812 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_1161
timestamp 1
transform 1 0 107916 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1167
timestamp 1
transform 1 0 108468 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_11
timestamp 1636968456
transform 1 0 2116 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_23
timestamp 1636968456
transform 1 0 3220 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_35
timestamp 1636968456
transform 1 0 4324 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_47
timestamp 1
transform 1 0 5428 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_129_55
timestamp 1
transform 1 0 6164 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_57
timestamp 1636968456
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_69
timestamp 1636968456
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_81
timestamp 1636968456
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_93
timestamp 1636968456
transform 1 0 9660 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_105
timestamp 1
transform 1 0 10764 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_111
timestamp 1
transform 1 0 11316 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_113
timestamp 1636968456
transform 1 0 11500 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_125
timestamp 1636968456
transform 1 0 12604 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_137
timestamp 1636968456
transform 1 0 13708 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_149
timestamp 1636968456
transform 1 0 14812 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_161
timestamp 1
transform 1 0 15916 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_167
timestamp 1
transform 1 0 16468 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_169
timestamp 1636968456
transform 1 0 16652 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_181
timestamp 1636968456
transform 1 0 17756 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_193
timestamp 1636968456
transform 1 0 18860 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_205
timestamp 1636968456
transform 1 0 19964 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_217
timestamp 1
transform 1 0 21068 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_223
timestamp 1
transform 1 0 21620 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_225
timestamp 1636968456
transform 1 0 21804 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_237
timestamp 1636968456
transform 1 0 22908 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_249
timestamp 1636968456
transform 1 0 24012 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_261
timestamp 1636968456
transform 1 0 25116 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_273
timestamp 1
transform 1 0 26220 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_279
timestamp 1
transform 1 0 26772 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_281
timestamp 1636968456
transform 1 0 26956 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_293
timestamp 1636968456
transform 1 0 28060 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_305
timestamp 1636968456
transform 1 0 29164 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_317
timestamp 1636968456
transform 1 0 30268 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_329
timestamp 1
transform 1 0 31372 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_335
timestamp 1
transform 1 0 31924 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_337
timestamp 1636968456
transform 1 0 32108 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_349
timestamp 1636968456
transform 1 0 33212 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_361
timestamp 1636968456
transform 1 0 34316 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_373
timestamp 1636968456
transform 1 0 35420 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_385
timestamp 1
transform 1 0 36524 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_391
timestamp 1
transform 1 0 37076 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_393
timestamp 1636968456
transform 1 0 37260 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_405
timestamp 1636968456
transform 1 0 38364 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_417
timestamp 1636968456
transform 1 0 39468 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_429
timestamp 1636968456
transform 1 0 40572 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_441
timestamp 1
transform 1 0 41676 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_447
timestamp 1
transform 1 0 42228 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_449
timestamp 1636968456
transform 1 0 42412 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_129_461
timestamp 1
transform 1 0 43516 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_465
timestamp 1
transform 1 0 43884 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_129_497
timestamp 1
transform 1 0 46828 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_503
timestamp 1
transform 1 0 47380 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_505
timestamp 1636968456
transform 1 0 47564 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_517
timestamp 1636968456
transform 1 0 48668 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_529
timestamp 1636968456
transform 1 0 49772 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_541
timestamp 1636968456
transform 1 0 50876 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_553
timestamp 1
transform 1 0 51980 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_559
timestamp 1
transform 1 0 52532 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_561
timestamp 1636968456
transform 1 0 52716 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_573
timestamp 1636968456
transform 1 0 53820 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_585
timestamp 1636968456
transform 1 0 54924 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_597
timestamp 1636968456
transform 1 0 56028 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_609
timestamp 1
transform 1 0 57132 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_615
timestamp 1
transform 1 0 57684 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_617
timestamp 1636968456
transform 1 0 57868 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_629
timestamp 1636968456
transform 1 0 58972 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_641
timestamp 1636968456
transform 1 0 60076 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_653
timestamp 1636968456
transform 1 0 61180 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_665
timestamp 1
transform 1 0 62284 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_671
timestamp 1
transform 1 0 62836 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_673
timestamp 1636968456
transform 1 0 63020 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_685
timestamp 1636968456
transform 1 0 64124 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_697
timestamp 1636968456
transform 1 0 65228 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_709
timestamp 1636968456
transform 1 0 66332 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_721
timestamp 1
transform 1 0 67436 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_727
timestamp 1
transform 1 0 67988 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_729
timestamp 1636968456
transform 1 0 68172 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_741
timestamp 1636968456
transform 1 0 69276 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_753
timestamp 1636968456
transform 1 0 70380 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_765
timestamp 1636968456
transform 1 0 71484 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_777
timestamp 1
transform 1 0 72588 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_783
timestamp 1
transform 1 0 73140 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_129_785
timestamp 1
transform 1 0 73324 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_808
timestamp 1636968456
transform 1 0 75440 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_820
timestamp 1636968456
transform 1 0 76544 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_832
timestamp 1
transform 1 0 77648 0 -1 72896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_129_841
timestamp 1636968456
transform 1 0 78476 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_853
timestamp 1636968456
transform 1 0 79580 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_865
timestamp 1636968456
transform 1 0 80684 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_877
timestamp 1636968456
transform 1 0 81788 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_889
timestamp 1
transform 1 0 82892 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_895
timestamp 1
transform 1 0 83444 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_897
timestamp 1636968456
transform 1 0 83628 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_909
timestamp 1636968456
transform 1 0 84732 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_921
timestamp 1636968456
transform 1 0 85836 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_933
timestamp 1636968456
transform 1 0 86940 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_945
timestamp 1
transform 1 0 88044 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_951
timestamp 1
transform 1 0 88596 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_953
timestamp 1636968456
transform 1 0 88780 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_965
timestamp 1636968456
transform 1 0 89884 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_977
timestamp 1636968456
transform 1 0 90988 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_989
timestamp 1636968456
transform 1 0 92092 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_1001
timestamp 1
transform 1 0 93196 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1007
timestamp 1
transform 1 0 93748 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1009
timestamp 1636968456
transform 1 0 93932 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1021
timestamp 1636968456
transform 1 0 95036 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1033
timestamp 1636968456
transform 1 0 96140 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1045
timestamp 1636968456
transform 1 0 97244 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_1057
timestamp 1
transform 1 0 98348 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1063
timestamp 1
transform 1 0 98900 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1065
timestamp 1636968456
transform 1 0 99084 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1077
timestamp 1636968456
transform 1 0 100188 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1089
timestamp 1636968456
transform 1 0 101292 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1101
timestamp 1636968456
transform 1 0 102396 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_1113
timestamp 1
transform 1 0 103500 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1119
timestamp 1
transform 1 0 104052 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1121
timestamp 1636968456
transform 1 0 104236 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1133
timestamp 1636968456
transform 1 0 105340 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1145
timestamp 1636968456
transform 1 0 106444 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_1157
timestamp 1
transform 1 0 107548 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_129_1165
timestamp 1
transform 1 0 108284 0 -1 72896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_130_8
timestamp 1636968456
transform 1 0 1840 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_20
timestamp 1
transform 1 0 2944 0 1 72896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_130_29
timestamp 1636968456
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_41
timestamp 1636968456
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_53
timestamp 1636968456
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_65
timestamp 1636968456
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_85
timestamp 1636968456
transform 1 0 8924 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_97
timestamp 1636968456
transform 1 0 10028 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_109
timestamp 1636968456
transform 1 0 11132 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_121
timestamp 1636968456
transform 1 0 12236 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_133
timestamp 1
transform 1 0 13340 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_139
timestamp 1
transform 1 0 13892 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_141
timestamp 1636968456
transform 1 0 14076 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_153
timestamp 1636968456
transform 1 0 15180 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_165
timestamp 1636968456
transform 1 0 16284 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_177
timestamp 1636968456
transform 1 0 17388 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_189
timestamp 1
transform 1 0 18492 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_195
timestamp 1
transform 1 0 19044 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_197
timestamp 1636968456
transform 1 0 19228 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_209
timestamp 1636968456
transform 1 0 20332 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_221
timestamp 1636968456
transform 1 0 21436 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_233
timestamp 1636968456
transform 1 0 22540 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_245
timestamp 1
transform 1 0 23644 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_251
timestamp 1
transform 1 0 24196 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_253
timestamp 1636968456
transform 1 0 24380 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_265
timestamp 1636968456
transform 1 0 25484 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_277
timestamp 1636968456
transform 1 0 26588 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_289
timestamp 1636968456
transform 1 0 27692 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_301
timestamp 1
transform 1 0 28796 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_307
timestamp 1
transform 1 0 29348 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_309
timestamp 1636968456
transform 1 0 29532 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_321
timestamp 1636968456
transform 1 0 30636 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_333
timestamp 1636968456
transform 1 0 31740 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_345
timestamp 1636968456
transform 1 0 32844 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_357
timestamp 1
transform 1 0 33948 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_363
timestamp 1
transform 1 0 34500 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_365
timestamp 1636968456
transform 1 0 34684 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_377
timestamp 1636968456
transform 1 0 35788 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_389
timestamp 1636968456
transform 1 0 36892 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_401
timestamp 1636968456
transform 1 0 37996 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_413
timestamp 1
transform 1 0 39100 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_419
timestamp 1
transform 1 0 39652 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_421
timestamp 1636968456
transform 1 0 39836 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_433
timestamp 1636968456
transform 1 0 40940 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_445
timestamp 1636968456
transform 1 0 42044 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_457
timestamp 1636968456
transform 1 0 43148 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_469
timestamp 1
transform 1 0 44252 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_475
timestamp 1
transform 1 0 44804 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_477
timestamp 1636968456
transform 1 0 44988 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_489
timestamp 1636968456
transform 1 0 46092 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_501
timestamp 1636968456
transform 1 0 47196 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_513
timestamp 1636968456
transform 1 0 48300 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_525
timestamp 1
transform 1 0 49404 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_531
timestamp 1
transform 1 0 49956 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_533
timestamp 1636968456
transform 1 0 50140 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_545
timestamp 1636968456
transform 1 0 51244 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_557
timestamp 1636968456
transform 1 0 52348 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_569
timestamp 1636968456
transform 1 0 53452 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_581
timestamp 1
transform 1 0 54556 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_587
timestamp 1
transform 1 0 55108 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_589
timestamp 1636968456
transform 1 0 55292 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_601
timestamp 1636968456
transform 1 0 56396 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_613
timestamp 1636968456
transform 1 0 57500 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_625
timestamp 1636968456
transform 1 0 58604 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_637
timestamp 1
transform 1 0 59708 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_643
timestamp 1
transform 1 0 60260 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_645
timestamp 1636968456
transform 1 0 60444 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_657
timestamp 1636968456
transform 1 0 61548 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_669
timestamp 1636968456
transform 1 0 62652 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_681
timestamp 1636968456
transform 1 0 63756 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_693
timestamp 1
transform 1 0 64860 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_699
timestamp 1
transform 1 0 65412 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_701
timestamp 1636968456
transform 1 0 65596 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_713
timestamp 1636968456
transform 1 0 66700 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_725
timestamp 1636968456
transform 1 0 67804 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_737
timestamp 1636968456
transform 1 0 68908 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_749
timestamp 1
transform 1 0 70012 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_755
timestamp 1
transform 1 0 70564 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_757
timestamp 1636968456
transform 1 0 70748 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_769
timestamp 1636968456
transform 1 0 71852 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_781
timestamp 1636968456
transform 1 0 72956 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_793
timestamp 1636968456
transform 1 0 74060 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_805
timestamp 1
transform 1 0 75164 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_811
timestamp 1
transform 1 0 75716 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_813
timestamp 1636968456
transform 1 0 75900 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_825
timestamp 1636968456
transform 1 0 77004 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_837
timestamp 1636968456
transform 1 0 78108 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_849
timestamp 1636968456
transform 1 0 79212 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_861
timestamp 1
transform 1 0 80316 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_867
timestamp 1
transform 1 0 80868 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_869
timestamp 1636968456
transform 1 0 81052 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_881
timestamp 1636968456
transform 1 0 82156 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_893
timestamp 1636968456
transform 1 0 83260 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_905
timestamp 1636968456
transform 1 0 84364 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_917
timestamp 1
transform 1 0 85468 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_923
timestamp 1
transform 1 0 86020 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_925
timestamp 1636968456
transform 1 0 86204 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_937
timestamp 1636968456
transform 1 0 87308 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_949
timestamp 1636968456
transform 1 0 88412 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_961
timestamp 1
transform 1 0 89516 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_130_970
timestamp 1
transform 1 0 90344 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_130_978
timestamp 1
transform 1 0 91080 0 1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_130_981
timestamp 1636968456
transform 1 0 91356 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_993
timestamp 1636968456
transform 1 0 92460 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1005
timestamp 1636968456
transform 1 0 93564 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1017
timestamp 1636968456
transform 1 0 94668 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_1029
timestamp 1
transform 1 0 95772 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1035
timestamp 1
transform 1 0 96324 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1037
timestamp 1636968456
transform 1 0 96508 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1049
timestamp 1636968456
transform 1 0 97612 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1061
timestamp 1636968456
transform 1 0 98716 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1073
timestamp 1636968456
transform 1 0 99820 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_1085
timestamp 1
transform 1 0 100924 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1091
timestamp 1
transform 1 0 101476 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1093
timestamp 1636968456
transform 1 0 101660 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1105
timestamp 1636968456
transform 1 0 102764 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1117
timestamp 1636968456
transform 1 0 103868 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1129
timestamp 1636968456
transform 1 0 104972 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_1141
timestamp 1
transform 1 0 106076 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1147
timestamp 1
transform 1 0 106628 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1149
timestamp 1636968456
transform 1 0 106812 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_130_1161
timestamp 1
transform 1 0 107916 0 1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_131_8
timestamp 1636968456
transform 1 0 1840 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_20
timestamp 1636968456
transform 1 0 2944 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_32
timestamp 1636968456
transform 1 0 4048 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_44
timestamp 1636968456
transform 1 0 5152 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_57
timestamp 1636968456
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_69
timestamp 1636968456
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_81
timestamp 1636968456
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_93
timestamp 1636968456
transform 1 0 9660 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_105
timestamp 1
transform 1 0 10764 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_111
timestamp 1
transform 1 0 11316 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_113
timestamp 1636968456
transform 1 0 11500 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_125
timestamp 1636968456
transform 1 0 12604 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_137
timestamp 1636968456
transform 1 0 13708 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_149
timestamp 1636968456
transform 1 0 14812 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_161
timestamp 1
transform 1 0 15916 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_167
timestamp 1
transform 1 0 16468 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_169
timestamp 1636968456
transform 1 0 16652 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_181
timestamp 1636968456
transform 1 0 17756 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_193
timestamp 1636968456
transform 1 0 18860 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_205
timestamp 1636968456
transform 1 0 19964 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_217
timestamp 1
transform 1 0 21068 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_223
timestamp 1
transform 1 0 21620 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_225
timestamp 1636968456
transform 1 0 21804 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_237
timestamp 1636968456
transform 1 0 22908 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_249
timestamp 1636968456
transform 1 0 24012 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_261
timestamp 1636968456
transform 1 0 25116 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_273
timestamp 1
transform 1 0 26220 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_279
timestamp 1
transform 1 0 26772 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_281
timestamp 1636968456
transform 1 0 26956 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_293
timestamp 1636968456
transform 1 0 28060 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_305
timestamp 1636968456
transform 1 0 29164 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_317
timestamp 1636968456
transform 1 0 30268 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_329
timestamp 1
transform 1 0 31372 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_335
timestamp 1
transform 1 0 31924 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_337
timestamp 1636968456
transform 1 0 32108 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_349
timestamp 1636968456
transform 1 0 33212 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_361
timestamp 1636968456
transform 1 0 34316 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_373
timestamp 1636968456
transform 1 0 35420 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_385
timestamp 1
transform 1 0 36524 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_391
timestamp 1
transform 1 0 37076 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_393
timestamp 1636968456
transform 1 0 37260 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_405
timestamp 1636968456
transform 1 0 38364 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_417
timestamp 1636968456
transform 1 0 39468 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_429
timestamp 1636968456
transform 1 0 40572 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_441
timestamp 1
transform 1 0 41676 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_447
timestamp 1
transform 1 0 42228 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_449
timestamp 1636968456
transform 1 0 42412 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_461
timestamp 1636968456
transform 1 0 43516 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_473
timestamp 1636968456
transform 1 0 44620 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_485
timestamp 1636968456
transform 1 0 45724 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_497
timestamp 1
transform 1 0 46828 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_503
timestamp 1
transform 1 0 47380 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_505
timestamp 1636968456
transform 1 0 47564 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_517
timestamp 1636968456
transform 1 0 48668 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_529
timestamp 1636968456
transform 1 0 49772 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_541
timestamp 1636968456
transform 1 0 50876 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_553
timestamp 1
transform 1 0 51980 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_559
timestamp 1
transform 1 0 52532 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_561
timestamp 1636968456
transform 1 0 52716 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_573
timestamp 1636968456
transform 1 0 53820 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_585
timestamp 1636968456
transform 1 0 54924 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_597
timestamp 1636968456
transform 1 0 56028 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_609
timestamp 1
transform 1 0 57132 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_615
timestamp 1
transform 1 0 57684 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_617
timestamp 1636968456
transform 1 0 57868 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_629
timestamp 1636968456
transform 1 0 58972 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_641
timestamp 1636968456
transform 1 0 60076 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_653
timestamp 1636968456
transform 1 0 61180 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_665
timestamp 1
transform 1 0 62284 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_671
timestamp 1
transform 1 0 62836 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_673
timestamp 1636968456
transform 1 0 63020 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_685
timestamp 1636968456
transform 1 0 64124 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_697
timestamp 1636968456
transform 1 0 65228 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_709
timestamp 1636968456
transform 1 0 66332 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_721
timestamp 1
transform 1 0 67436 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_727
timestamp 1
transform 1 0 67988 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_729
timestamp 1636968456
transform 1 0 68172 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_741
timestamp 1636968456
transform 1 0 69276 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_753
timestamp 1636968456
transform 1 0 70380 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_765
timestamp 1636968456
transform 1 0 71484 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_777
timestamp 1
transform 1 0 72588 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_783
timestamp 1
transform 1 0 73140 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_785
timestamp 1636968456
transform 1 0 73324 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_797
timestamp 1636968456
transform 1 0 74428 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_809
timestamp 1636968456
transform 1 0 75532 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_821
timestamp 1636968456
transform 1 0 76636 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_833
timestamp 1
transform 1 0 77740 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_839
timestamp 1
transform 1 0 78292 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_841
timestamp 1636968456
transform 1 0 78476 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_853
timestamp 1636968456
transform 1 0 79580 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_865
timestamp 1636968456
transform 1 0 80684 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_877
timestamp 1636968456
transform 1 0 81788 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_889
timestamp 1
transform 1 0 82892 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_895
timestamp 1
transform 1 0 83444 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_897
timestamp 1636968456
transform 1 0 83628 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_909
timestamp 1636968456
transform 1 0 84732 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_921
timestamp 1636968456
transform 1 0 85836 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_933
timestamp 1636968456
transform 1 0 86940 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_945
timestamp 1
transform 1 0 88044 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_951
timestamp 1
transform 1 0 88596 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_953
timestamp 1636968456
transform 1 0 88780 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_965
timestamp 1636968456
transform 1 0 89884 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_977
timestamp 1636968456
transform 1 0 90988 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_989
timestamp 1636968456
transform 1 0 92092 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_1001
timestamp 1
transform 1 0 93196 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_1007
timestamp 1
transform 1 0 93748 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1009
timestamp 1636968456
transform 1 0 93932 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1021
timestamp 1636968456
transform 1 0 95036 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1033
timestamp 1636968456
transform 1 0 96140 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1045
timestamp 1636968456
transform 1 0 97244 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_1057
timestamp 1
transform 1 0 98348 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_1063
timestamp 1
transform 1 0 98900 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1065
timestamp 1636968456
transform 1 0 99084 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1077
timestamp 1636968456
transform 1 0 100188 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1089
timestamp 1636968456
transform 1 0 101292 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1101
timestamp 1636968456
transform 1 0 102396 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_1113
timestamp 1
transform 1 0 103500 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_1119
timestamp 1
transform 1 0 104052 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1121
timestamp 1636968456
transform 1 0 104236 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1133
timestamp 1636968456
transform 1 0 105340 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1145
timestamp 1636968456
transform 1 0 106444 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_1157
timestamp 1
transform 1 0 107548 0 -1 73984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_132_8
timestamp 1636968456
transform 1 0 1840 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_20
timestamp 1
transform 1 0 2944 0 1 73984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_132_29
timestamp 1636968456
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_41
timestamp 1636968456
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_53
timestamp 1636968456
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_65
timestamp 1636968456
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1
transform 1 0 8188 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_85
timestamp 1636968456
transform 1 0 8924 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_97
timestamp 1636968456
transform 1 0 10028 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_109
timestamp 1636968456
transform 1 0 11132 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_121
timestamp 1636968456
transform 1 0 12236 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_133
timestamp 1
transform 1 0 13340 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_139
timestamp 1
transform 1 0 13892 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_141
timestamp 1636968456
transform 1 0 14076 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_153
timestamp 1636968456
transform 1 0 15180 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_165
timestamp 1636968456
transform 1 0 16284 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_177
timestamp 1636968456
transform 1 0 17388 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_189
timestamp 1
transform 1 0 18492 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_195
timestamp 1
transform 1 0 19044 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_197
timestamp 1636968456
transform 1 0 19228 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_209
timestamp 1636968456
transform 1 0 20332 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_221
timestamp 1636968456
transform 1 0 21436 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_233
timestamp 1636968456
transform 1 0 22540 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_245
timestamp 1
transform 1 0 23644 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_251
timestamp 1
transform 1 0 24196 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_253
timestamp 1636968456
transform 1 0 24380 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_265
timestamp 1636968456
transform 1 0 25484 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_277
timestamp 1636968456
transform 1 0 26588 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_289
timestamp 1636968456
transform 1 0 27692 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_301
timestamp 1
transform 1 0 28796 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_307
timestamp 1
transform 1 0 29348 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_309
timestamp 1636968456
transform 1 0 29532 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_321
timestamp 1636968456
transform 1 0 30636 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_333
timestamp 1636968456
transform 1 0 31740 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_345
timestamp 1636968456
transform 1 0 32844 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_357
timestamp 1
transform 1 0 33948 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_363
timestamp 1
transform 1 0 34500 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_365
timestamp 1636968456
transform 1 0 34684 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_377
timestamp 1636968456
transform 1 0 35788 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_389
timestamp 1636968456
transform 1 0 36892 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_401
timestamp 1636968456
transform 1 0 37996 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_413
timestamp 1
transform 1 0 39100 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_419
timestamp 1
transform 1 0 39652 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_421
timestamp 1636968456
transform 1 0 39836 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_433
timestamp 1636968456
transform 1 0 40940 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_445
timestamp 1636968456
transform 1 0 42044 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_457
timestamp 1636968456
transform 1 0 43148 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_469
timestamp 1
transform 1 0 44252 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_475
timestamp 1
transform 1 0 44804 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_477
timestamp 1636968456
transform 1 0 44988 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_489
timestamp 1636968456
transform 1 0 46092 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_501
timestamp 1636968456
transform 1 0 47196 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_513
timestamp 1636968456
transform 1 0 48300 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_525
timestamp 1
transform 1 0 49404 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_531
timestamp 1
transform 1 0 49956 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_533
timestamp 1636968456
transform 1 0 50140 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_545
timestamp 1636968456
transform 1 0 51244 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_557
timestamp 1636968456
transform 1 0 52348 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_569
timestamp 1636968456
transform 1 0 53452 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_581
timestamp 1
transform 1 0 54556 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_587
timestamp 1
transform 1 0 55108 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_589
timestamp 1636968456
transform 1 0 55292 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_601
timestamp 1636968456
transform 1 0 56396 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_613
timestamp 1636968456
transform 1 0 57500 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_625
timestamp 1636968456
transform 1 0 58604 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_637
timestamp 1
transform 1 0 59708 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_643
timestamp 1
transform 1 0 60260 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_645
timestamp 1636968456
transform 1 0 60444 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_657
timestamp 1636968456
transform 1 0 61548 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_669
timestamp 1636968456
transform 1 0 62652 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_681
timestamp 1636968456
transform 1 0 63756 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_693
timestamp 1
transform 1 0 64860 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_699
timestamp 1
transform 1 0 65412 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_701
timestamp 1636968456
transform 1 0 65596 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_713
timestamp 1636968456
transform 1 0 66700 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_725
timestamp 1636968456
transform 1 0 67804 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_737
timestamp 1636968456
transform 1 0 68908 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_749
timestamp 1
transform 1 0 70012 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_755
timestamp 1
transform 1 0 70564 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_757
timestamp 1636968456
transform 1 0 70748 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_769
timestamp 1636968456
transform 1 0 71852 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_781
timestamp 1636968456
transform 1 0 72956 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_793
timestamp 1636968456
transform 1 0 74060 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_805
timestamp 1
transform 1 0 75164 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_811
timestamp 1
transform 1 0 75716 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_813
timestamp 1636968456
transform 1 0 75900 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_825
timestamp 1636968456
transform 1 0 77004 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_837
timestamp 1636968456
transform 1 0 78108 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_849
timestamp 1636968456
transform 1 0 79212 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_861
timestamp 1
transform 1 0 80316 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_867
timestamp 1
transform 1 0 80868 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_869
timestamp 1636968456
transform 1 0 81052 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_881
timestamp 1636968456
transform 1 0 82156 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_893
timestamp 1636968456
transform 1 0 83260 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_905
timestamp 1636968456
transform 1 0 84364 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_917
timestamp 1
transform 1 0 85468 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_923
timestamp 1
transform 1 0 86020 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_925
timestamp 1636968456
transform 1 0 86204 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_937
timestamp 1636968456
transform 1 0 87308 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_949
timestamp 1636968456
transform 1 0 88412 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_961
timestamp 1636968456
transform 1 0 89516 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_973
timestamp 1
transform 1 0 90620 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_979
timestamp 1
transform 1 0 91172 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_981
timestamp 1636968456
transform 1 0 91356 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_993
timestamp 1636968456
transform 1 0 92460 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1005
timestamp 1636968456
transform 1 0 93564 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1017
timestamp 1636968456
transform 1 0 94668 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_1029
timestamp 1
transform 1 0 95772 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1035
timestamp 1
transform 1 0 96324 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1037
timestamp 1636968456
transform 1 0 96508 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1049
timestamp 1636968456
transform 1 0 97612 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1061
timestamp 1636968456
transform 1 0 98716 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1073
timestamp 1636968456
transform 1 0 99820 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_1085
timestamp 1
transform 1 0 100924 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1091
timestamp 1
transform 1 0 101476 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1093
timestamp 1636968456
transform 1 0 101660 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1105
timestamp 1636968456
transform 1 0 102764 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1117
timestamp 1636968456
transform 1 0 103868 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1129
timestamp 1636968456
transform 1 0 104972 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_1141
timestamp 1
transform 1 0 106076 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1147
timestamp 1
transform 1 0 106628 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1149
timestamp 1636968456
transform 1 0 106812 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_132_1161
timestamp 1
transform 1 0 107916 0 1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_133_3
timestamp 1636968456
transform 1 0 1380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_15
timestamp 1636968456
transform 1 0 2484 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_27
timestamp 1636968456
transform 1 0 3588 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_39
timestamp 1636968456
transform 1 0 4692 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_51
timestamp 1
transform 1 0 5796 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_133_55
timestamp 1
transform 1 0 6164 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_57
timestamp 1636968456
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_69
timestamp 1636968456
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_81
timestamp 1636968456
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_93
timestamp 1636968456
transform 1 0 9660 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_105
timestamp 1
transform 1 0 10764 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_111
timestamp 1
transform 1 0 11316 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_113
timestamp 1636968456
transform 1 0 11500 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_125
timestamp 1636968456
transform 1 0 12604 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_137
timestamp 1636968456
transform 1 0 13708 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_149
timestamp 1636968456
transform 1 0 14812 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_161
timestamp 1
transform 1 0 15916 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_167
timestamp 1
transform 1 0 16468 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_169
timestamp 1636968456
transform 1 0 16652 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_181
timestamp 1636968456
transform 1 0 17756 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_193
timestamp 1636968456
transform 1 0 18860 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_205
timestamp 1636968456
transform 1 0 19964 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_217
timestamp 1
transform 1 0 21068 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_223
timestamp 1
transform 1 0 21620 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_225
timestamp 1636968456
transform 1 0 21804 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_237
timestamp 1636968456
transform 1 0 22908 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_249
timestamp 1636968456
transform 1 0 24012 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_261
timestamp 1636968456
transform 1 0 25116 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_273
timestamp 1
transform 1 0 26220 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_279
timestamp 1
transform 1 0 26772 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_281
timestamp 1636968456
transform 1 0 26956 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_293
timestamp 1636968456
transform 1 0 28060 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_305
timestamp 1636968456
transform 1 0 29164 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_317
timestamp 1636968456
transform 1 0 30268 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_329
timestamp 1
transform 1 0 31372 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_335
timestamp 1
transform 1 0 31924 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_337
timestamp 1636968456
transform 1 0 32108 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_349
timestamp 1636968456
transform 1 0 33212 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_361
timestamp 1636968456
transform 1 0 34316 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_373
timestamp 1636968456
transform 1 0 35420 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_385
timestamp 1
transform 1 0 36524 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_391
timestamp 1
transform 1 0 37076 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_393
timestamp 1636968456
transform 1 0 37260 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_405
timestamp 1636968456
transform 1 0 38364 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_417
timestamp 1636968456
transform 1 0 39468 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_429
timestamp 1636968456
transform 1 0 40572 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_441
timestamp 1
transform 1 0 41676 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_447
timestamp 1
transform 1 0 42228 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_449
timestamp 1636968456
transform 1 0 42412 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_461
timestamp 1636968456
transform 1 0 43516 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_473
timestamp 1636968456
transform 1 0 44620 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_485
timestamp 1636968456
transform 1 0 45724 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_497
timestamp 1
transform 1 0 46828 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_503
timestamp 1
transform 1 0 47380 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_505
timestamp 1636968456
transform 1 0 47564 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_517
timestamp 1636968456
transform 1 0 48668 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_529
timestamp 1636968456
transform 1 0 49772 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_541
timestamp 1636968456
transform 1 0 50876 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_553
timestamp 1
transform 1 0 51980 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_559
timestamp 1
transform 1 0 52532 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_561
timestamp 1636968456
transform 1 0 52716 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_573
timestamp 1636968456
transform 1 0 53820 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_585
timestamp 1636968456
transform 1 0 54924 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_597
timestamp 1636968456
transform 1 0 56028 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_609
timestamp 1
transform 1 0 57132 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_615
timestamp 1
transform 1 0 57684 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_617
timestamp 1636968456
transform 1 0 57868 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_629
timestamp 1636968456
transform 1 0 58972 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_641
timestamp 1636968456
transform 1 0 60076 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_653
timestamp 1636968456
transform 1 0 61180 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_665
timestamp 1
transform 1 0 62284 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_671
timestamp 1
transform 1 0 62836 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_673
timestamp 1636968456
transform 1 0 63020 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_685
timestamp 1636968456
transform 1 0 64124 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_697
timestamp 1636968456
transform 1 0 65228 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_709
timestamp 1636968456
transform 1 0 66332 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_721
timestamp 1
transform 1 0 67436 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_727
timestamp 1
transform 1 0 67988 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_729
timestamp 1636968456
transform 1 0 68172 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_741
timestamp 1636968456
transform 1 0 69276 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_753
timestamp 1636968456
transform 1 0 70380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_765
timestamp 1636968456
transform 1 0 71484 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_777
timestamp 1
transform 1 0 72588 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_783
timestamp 1
transform 1 0 73140 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_785
timestamp 1636968456
transform 1 0 73324 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_797
timestamp 1636968456
transform 1 0 74428 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_809
timestamp 1636968456
transform 1 0 75532 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_821
timestamp 1636968456
transform 1 0 76636 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_833
timestamp 1
transform 1 0 77740 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_839
timestamp 1
transform 1 0 78292 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_841
timestamp 1636968456
transform 1 0 78476 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_853
timestamp 1636968456
transform 1 0 79580 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_865
timestamp 1636968456
transform 1 0 80684 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_877
timestamp 1
transform 1 0 81788 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_883
timestamp 1
transform 1 0 82340 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_133_886
timestamp 1
transform 1 0 82616 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_133_894
timestamp 1
transform 1 0 83352 0 -1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_133_897
timestamp 1636968456
transform 1 0 83628 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_909
timestamp 1636968456
transform 1 0 84732 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_921
timestamp 1636968456
transform 1 0 85836 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_933
timestamp 1636968456
transform 1 0 86940 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_945
timestamp 1
transform 1 0 88044 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_951
timestamp 1
transform 1 0 88596 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_953
timestamp 1636968456
transform 1 0 88780 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_965
timestamp 1636968456
transform 1 0 89884 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_977
timestamp 1636968456
transform 1 0 90988 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_989
timestamp 1636968456
transform 1 0 92092 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_1001
timestamp 1
transform 1 0 93196 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_1007
timestamp 1
transform 1 0 93748 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1009
timestamp 1636968456
transform 1 0 93932 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1021
timestamp 1636968456
transform 1 0 95036 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1033
timestamp 1636968456
transform 1 0 96140 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1045
timestamp 1636968456
transform 1 0 97244 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_1057
timestamp 1
transform 1 0 98348 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_1063
timestamp 1
transform 1 0 98900 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1065
timestamp 1636968456
transform 1 0 99084 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1077
timestamp 1636968456
transform 1 0 100188 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1089
timestamp 1636968456
transform 1 0 101292 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1101
timestamp 1636968456
transform 1 0 102396 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_1113
timestamp 1
transform 1 0 103500 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_1119
timestamp 1
transform 1 0 104052 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1121
timestamp 1636968456
transform 1 0 104236 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1133
timestamp 1636968456
transform 1 0 105340 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1145
timestamp 1636968456
transform 1 0 106444 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_1157
timestamp 1
transform 1 0 107548 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_133_1165
timestamp 1
transform 1 0 108284 0 -1 75072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_134_8
timestamp 1636968456
transform 1 0 1840 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_20
timestamp 1
transform 1 0 2944 0 1 75072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_134_29
timestamp 1636968456
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_41
timestamp 1636968456
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_53
timestamp 1636968456
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_65
timestamp 1636968456
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_85
timestamp 1636968456
transform 1 0 8924 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_97
timestamp 1636968456
transform 1 0 10028 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_109
timestamp 1636968456
transform 1 0 11132 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_121
timestamp 1636968456
transform 1 0 12236 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_133
timestamp 1
transform 1 0 13340 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_139
timestamp 1
transform 1 0 13892 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_141
timestamp 1636968456
transform 1 0 14076 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_153
timestamp 1636968456
transform 1 0 15180 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_165
timestamp 1636968456
transform 1 0 16284 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_177
timestamp 1636968456
transform 1 0 17388 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_189
timestamp 1
transform 1 0 18492 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_195
timestamp 1
transform 1 0 19044 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_197
timestamp 1636968456
transform 1 0 19228 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_209
timestamp 1636968456
transform 1 0 20332 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_221
timestamp 1636968456
transform 1 0 21436 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_233
timestamp 1636968456
transform 1 0 22540 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_245
timestamp 1
transform 1 0 23644 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_251
timestamp 1
transform 1 0 24196 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_253
timestamp 1636968456
transform 1 0 24380 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_265
timestamp 1636968456
transform 1 0 25484 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_277
timestamp 1636968456
transform 1 0 26588 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_289
timestamp 1636968456
transform 1 0 27692 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_301
timestamp 1
transform 1 0 28796 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_307
timestamp 1
transform 1 0 29348 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_309
timestamp 1636968456
transform 1 0 29532 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_321
timestamp 1636968456
transform 1 0 30636 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_333
timestamp 1636968456
transform 1 0 31740 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_345
timestamp 1636968456
transform 1 0 32844 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_357
timestamp 1
transform 1 0 33948 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_363
timestamp 1
transform 1 0 34500 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_365
timestamp 1636968456
transform 1 0 34684 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_377
timestamp 1636968456
transform 1 0 35788 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_389
timestamp 1636968456
transform 1 0 36892 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_401
timestamp 1636968456
transform 1 0 37996 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_413
timestamp 1
transform 1 0 39100 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_419
timestamp 1
transform 1 0 39652 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_421
timestamp 1636968456
transform 1 0 39836 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_433
timestamp 1636968456
transform 1 0 40940 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_445
timestamp 1636968456
transform 1 0 42044 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_457
timestamp 1636968456
transform 1 0 43148 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_469
timestamp 1
transform 1 0 44252 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_475
timestamp 1
transform 1 0 44804 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_477
timestamp 1636968456
transform 1 0 44988 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_489
timestamp 1636968456
transform 1 0 46092 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_501
timestamp 1636968456
transform 1 0 47196 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_513
timestamp 1636968456
transform 1 0 48300 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_525
timestamp 1
transform 1 0 49404 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_531
timestamp 1
transform 1 0 49956 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_533
timestamp 1636968456
transform 1 0 50140 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_545
timestamp 1636968456
transform 1 0 51244 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_557
timestamp 1636968456
transform 1 0 52348 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_569
timestamp 1636968456
transform 1 0 53452 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_581
timestamp 1
transform 1 0 54556 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_587
timestamp 1
transform 1 0 55108 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_589
timestamp 1636968456
transform 1 0 55292 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_601
timestamp 1636968456
transform 1 0 56396 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_613
timestamp 1636968456
transform 1 0 57500 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_625
timestamp 1636968456
transform 1 0 58604 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_637
timestamp 1
transform 1 0 59708 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_643
timestamp 1
transform 1 0 60260 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_645
timestamp 1636968456
transform 1 0 60444 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_657
timestamp 1636968456
transform 1 0 61548 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_669
timestamp 1636968456
transform 1 0 62652 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_681
timestamp 1636968456
transform 1 0 63756 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_693
timestamp 1
transform 1 0 64860 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_699
timestamp 1
transform 1 0 65412 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_701
timestamp 1636968456
transform 1 0 65596 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_713
timestamp 1636968456
transform 1 0 66700 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_725
timestamp 1636968456
transform 1 0 67804 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_737
timestamp 1636968456
transform 1 0 68908 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_749
timestamp 1
transform 1 0 70012 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_755
timestamp 1
transform 1 0 70564 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_757
timestamp 1636968456
transform 1 0 70748 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_769
timestamp 1636968456
transform 1 0 71852 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_781
timestamp 1636968456
transform 1 0 72956 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_793
timestamp 1636968456
transform 1 0 74060 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_805
timestamp 1
transform 1 0 75164 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_811
timestamp 1
transform 1 0 75716 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_813
timestamp 1636968456
transform 1 0 75900 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_825
timestamp 1636968456
transform 1 0 77004 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_837
timestamp 1636968456
transform 1 0 78108 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_849
timestamp 1636968456
transform 1 0 79212 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_861
timestamp 1
transform 1 0 80316 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_867
timestamp 1
transform 1 0 80868 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_869
timestamp 1
transform 1 0 81052 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_134_906
timestamp 1
transform 1 0 84456 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_134_914
timestamp 1
transform 1 0 85192 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_134_920
timestamp 1
transform 1 0 85744 0 1 75072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_134_934
timestamp 1636968456
transform 1 0 87032 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_946
timestamp 1636968456
transform 1 0 88136 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_958
timestamp 1636968456
transform 1 0 89240 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_970
timestamp 1
transform 1 0 90344 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_134_976
timestamp 1
transform 1 0 90896 0 1 75072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_134_981
timestamp 1636968456
transform 1 0 91356 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_993
timestamp 1636968456
transform 1 0 92460 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1005
timestamp 1636968456
transform 1 0 93564 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1017
timestamp 1636968456
transform 1 0 94668 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_1029
timestamp 1
transform 1 0 95772 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_1035
timestamp 1
transform 1 0 96324 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1037
timestamp 1636968456
transform 1 0 96508 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1049
timestamp 1636968456
transform 1 0 97612 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1061
timestamp 1636968456
transform 1 0 98716 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1073
timestamp 1636968456
transform 1 0 99820 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_1085
timestamp 1
transform 1 0 100924 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_1091
timestamp 1
transform 1 0 101476 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1093
timestamp 1636968456
transform 1 0 101660 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1105
timestamp 1636968456
transform 1 0 102764 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1117
timestamp 1636968456
transform 1 0 103868 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1129
timestamp 1636968456
transform 1 0 104972 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_1141
timestamp 1
transform 1 0 106076 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_1147
timestamp 1
transform 1 0 106628 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1149
timestamp 1636968456
transform 1 0 106812 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_134_1161
timestamp 1
transform 1 0 107916 0 1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_135_8
timestamp 1636968456
transform 1 0 1840 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_20
timestamp 1636968456
transform 1 0 2944 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_32
timestamp 1636968456
transform 1 0 4048 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_44
timestamp 1636968456
transform 1 0 5152 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_57
timestamp 1636968456
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_69
timestamp 1636968456
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_81
timestamp 1636968456
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_93
timestamp 1636968456
transform 1 0 9660 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_105
timestamp 1
transform 1 0 10764 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_111
timestamp 1
transform 1 0 11316 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_113
timestamp 1636968456
transform 1 0 11500 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_125
timestamp 1636968456
transform 1 0 12604 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_137
timestamp 1636968456
transform 1 0 13708 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_149
timestamp 1636968456
transform 1 0 14812 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_161
timestamp 1
transform 1 0 15916 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_167
timestamp 1
transform 1 0 16468 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_169
timestamp 1636968456
transform 1 0 16652 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_181
timestamp 1636968456
transform 1 0 17756 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_193
timestamp 1636968456
transform 1 0 18860 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_205
timestamp 1636968456
transform 1 0 19964 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_217
timestamp 1
transform 1 0 21068 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_223
timestamp 1
transform 1 0 21620 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_225
timestamp 1636968456
transform 1 0 21804 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_237
timestamp 1636968456
transform 1 0 22908 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_249
timestamp 1636968456
transform 1 0 24012 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_261
timestamp 1636968456
transform 1 0 25116 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_273
timestamp 1
transform 1 0 26220 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_279
timestamp 1
transform 1 0 26772 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_281
timestamp 1636968456
transform 1 0 26956 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_293
timestamp 1636968456
transform 1 0 28060 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_305
timestamp 1636968456
transform 1 0 29164 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_317
timestamp 1636968456
transform 1 0 30268 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_329
timestamp 1
transform 1 0 31372 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_335
timestamp 1
transform 1 0 31924 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_337
timestamp 1636968456
transform 1 0 32108 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_349
timestamp 1636968456
transform 1 0 33212 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_361
timestamp 1636968456
transform 1 0 34316 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_373
timestamp 1636968456
transform 1 0 35420 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_385
timestamp 1
transform 1 0 36524 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_391
timestamp 1
transform 1 0 37076 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_393
timestamp 1636968456
transform 1 0 37260 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_405
timestamp 1636968456
transform 1 0 38364 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_417
timestamp 1636968456
transform 1 0 39468 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_429
timestamp 1636968456
transform 1 0 40572 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_441
timestamp 1
transform 1 0 41676 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_447
timestamp 1
transform 1 0 42228 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_449
timestamp 1636968456
transform 1 0 42412 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_461
timestamp 1636968456
transform 1 0 43516 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_473
timestamp 1636968456
transform 1 0 44620 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_485
timestamp 1636968456
transform 1 0 45724 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_497
timestamp 1
transform 1 0 46828 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_503
timestamp 1
transform 1 0 47380 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_505
timestamp 1636968456
transform 1 0 47564 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_517
timestamp 1636968456
transform 1 0 48668 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_529
timestamp 1636968456
transform 1 0 49772 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_541
timestamp 1636968456
transform 1 0 50876 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_553
timestamp 1
transform 1 0 51980 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_559
timestamp 1
transform 1 0 52532 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_561
timestamp 1636968456
transform 1 0 52716 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_573
timestamp 1636968456
transform 1 0 53820 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_585
timestamp 1636968456
transform 1 0 54924 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_597
timestamp 1636968456
transform 1 0 56028 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_609
timestamp 1
transform 1 0 57132 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_615
timestamp 1
transform 1 0 57684 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_617
timestamp 1636968456
transform 1 0 57868 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_629
timestamp 1636968456
transform 1 0 58972 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_641
timestamp 1636968456
transform 1 0 60076 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_653
timestamp 1636968456
transform 1 0 61180 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_665
timestamp 1
transform 1 0 62284 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_671
timestamp 1
transform 1 0 62836 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_673
timestamp 1636968456
transform 1 0 63020 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_685
timestamp 1636968456
transform 1 0 64124 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_697
timestamp 1636968456
transform 1 0 65228 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_709
timestamp 1636968456
transform 1 0 66332 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_721
timestamp 1
transform 1 0 67436 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_727
timestamp 1
transform 1 0 67988 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_729
timestamp 1636968456
transform 1 0 68172 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_741
timestamp 1636968456
transform 1 0 69276 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_753
timestamp 1636968456
transform 1 0 70380 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_765
timestamp 1636968456
transform 1 0 71484 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_777
timestamp 1
transform 1 0 72588 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_783
timestamp 1
transform 1 0 73140 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_785
timestamp 1636968456
transform 1 0 73324 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_797
timestamp 1636968456
transform 1 0 74428 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_809
timestamp 1636968456
transform 1 0 75532 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_821
timestamp 1636968456
transform 1 0 76636 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_833
timestamp 1
transform 1 0 77740 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_839
timestamp 1
transform 1 0 78292 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_841
timestamp 1636968456
transform 1 0 78476 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_853
timestamp 1636968456
transform 1 0 79580 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_865
timestamp 1636968456
transform 1 0 80684 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_877
timestamp 1
transform 1 0 81788 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_135_885
timestamp 1
transform 1 0 82524 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_135_892
timestamp 1
transform 1 0 83168 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_924
timestamp 1
transform 1 0 86112 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_135_929
timestamp 1
transform 1 0 86572 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_135_955
timestamp 1
transform 1 0 88964 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_135_963
timestamp 1
transform 1 0 89700 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_135_973
timestamp 1
transform 1 0 90620 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_980
timestamp 1636968456
transform 1 0 91264 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_992
timestamp 1636968456
transform 1 0 92368 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_1004
timestamp 1
transform 1 0 93472 0 -1 76160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1009
timestamp 1636968456
transform 1 0 93932 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1021
timestamp 1636968456
transform 1 0 95036 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1033
timestamp 1636968456
transform 1 0 96140 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1045
timestamp 1636968456
transform 1 0 97244 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_1057
timestamp 1
transform 1 0 98348 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_1063
timestamp 1
transform 1 0 98900 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1065
timestamp 1636968456
transform 1 0 99084 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1077
timestamp 1636968456
transform 1 0 100188 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1089
timestamp 1636968456
transform 1 0 101292 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1101
timestamp 1636968456
transform 1 0 102396 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_1113
timestamp 1
transform 1 0 103500 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_1119
timestamp 1
transform 1 0 104052 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1121
timestamp 1636968456
transform 1 0 104236 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1133
timestamp 1636968456
transform 1 0 105340 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1145
timestamp 1636968456
transform 1 0 106444 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_1157
timestamp 1
transform 1 0 107548 0 -1 76160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_136_8
timestamp 1636968456
transform 1 0 1840 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_20
timestamp 1
transform 1 0 2944 0 1 76160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_136_29
timestamp 1636968456
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_41
timestamp 1636968456
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_53
timestamp 1636968456
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_65
timestamp 1636968456
transform 1 0 7084 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1
transform 1 0 8188 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1
transform 1 0 8740 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_85
timestamp 1636968456
transform 1 0 8924 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_97
timestamp 1636968456
transform 1 0 10028 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_109
timestamp 1636968456
transform 1 0 11132 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_121
timestamp 1636968456
transform 1 0 12236 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_133
timestamp 1
transform 1 0 13340 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_139
timestamp 1
transform 1 0 13892 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_141
timestamp 1636968456
transform 1 0 14076 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_153
timestamp 1636968456
transform 1 0 15180 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_165
timestamp 1636968456
transform 1 0 16284 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_177
timestamp 1636968456
transform 1 0 17388 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_189
timestamp 1
transform 1 0 18492 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_195
timestamp 1
transform 1 0 19044 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_197
timestamp 1636968456
transform 1 0 19228 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_209
timestamp 1636968456
transform 1 0 20332 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_221
timestamp 1
transform 1 0 21436 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_136_246
timestamp 1
transform 1 0 23736 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_136_253
timestamp 1
transform 1 0 24380 0 1 76160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_136_260
timestamp 1636968456
transform 1 0 25024 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_272
timestamp 1636968456
transform 1 0 26128 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_284
timestamp 1636968456
transform 1 0 27232 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_296
timestamp 1
transform 1 0 28336 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_307
timestamp 1
transform 1 0 29348 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_309
timestamp 1636968456
transform 1 0 29532 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_136_321
timestamp 1
transform 1 0 30636 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_136_329
timestamp 1
transform 1 0 31372 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_136_335
timestamp 1
transform 1 0 31924 0 1 76160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_136_343
timestamp 1636968456
transform 1 0 32660 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_355
timestamp 1
transform 1 0 33764 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_136_363
timestamp 1
transform 1 0 34500 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_365
timestamp 1636968456
transform 1 0 34684 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_377
timestamp 1636968456
transform 1 0 35788 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_389
timestamp 1636968456
transform 1 0 36892 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_401
timestamp 1636968456
transform 1 0 37996 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_413
timestamp 1
transform 1 0 39100 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_419
timestamp 1
transform 1 0 39652 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_421
timestamp 1636968456
transform 1 0 39836 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_433
timestamp 1636968456
transform 1 0 40940 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_445
timestamp 1636968456
transform 1 0 42044 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_457
timestamp 1636968456
transform 1 0 43148 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_469
timestamp 1
transform 1 0 44252 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_475
timestamp 1
transform 1 0 44804 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_477
timestamp 1636968456
transform 1 0 44988 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_489
timestamp 1636968456
transform 1 0 46092 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_501
timestamp 1636968456
transform 1 0 47196 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_513
timestamp 1636968456
transform 1 0 48300 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_525
timestamp 1
transform 1 0 49404 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_531
timestamp 1
transform 1 0 49956 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_533
timestamp 1636968456
transform 1 0 50140 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_545
timestamp 1636968456
transform 1 0 51244 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_557
timestamp 1636968456
transform 1 0 52348 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_569
timestamp 1636968456
transform 1 0 53452 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_581
timestamp 1
transform 1 0 54556 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_587
timestamp 1
transform 1 0 55108 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_589
timestamp 1636968456
transform 1 0 55292 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_601
timestamp 1636968456
transform 1 0 56396 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_613
timestamp 1636968456
transform 1 0 57500 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_625
timestamp 1636968456
transform 1 0 58604 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_637
timestamp 1
transform 1 0 59708 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_643
timestamp 1
transform 1 0 60260 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_645
timestamp 1636968456
transform 1 0 60444 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_657
timestamp 1636968456
transform 1 0 61548 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_669
timestamp 1636968456
transform 1 0 62652 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_681
timestamp 1636968456
transform 1 0 63756 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_693
timestamp 1
transform 1 0 64860 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_699
timestamp 1
transform 1 0 65412 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_701
timestamp 1636968456
transform 1 0 65596 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_713
timestamp 1636968456
transform 1 0 66700 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_725
timestamp 1636968456
transform 1 0 67804 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_737
timestamp 1636968456
transform 1 0 68908 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_749
timestamp 1
transform 1 0 70012 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_755
timestamp 1
transform 1 0 70564 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_757
timestamp 1636968456
transform 1 0 70748 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_769
timestamp 1636968456
transform 1 0 71852 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_781
timestamp 1636968456
transform 1 0 72956 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_793
timestamp 1636968456
transform 1 0 74060 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_805
timestamp 1
transform 1 0 75164 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_811
timestamp 1
transform 1 0 75716 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_813
timestamp 1636968456
transform 1 0 75900 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_825
timestamp 1636968456
transform 1 0 77004 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_837
timestamp 1636968456
transform 1 0 78108 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_849
timestamp 1636968456
transform 1 0 79212 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_861
timestamp 1
transform 1 0 80316 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_867
timestamp 1
transform 1 0 80868 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_869
timestamp 1636968456
transform 1 0 81052 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_886
timestamp 1
transform 1 0 82616 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_136_914
timestamp 1
transform 1 0 85192 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_918
timestamp 1
transform 1 0 85560 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_136_948
timestamp 1
transform 1 0 88320 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_136_958
timestamp 1
transform 1 0 89240 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_962
timestamp 1
transform 1 0 89608 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_968
timestamp 1636968456
transform 1 0 90160 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_981
timestamp 1636968456
transform 1 0 91356 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_993
timestamp 1636968456
transform 1 0 92460 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1005
timestamp 1636968456
transform 1 0 93564 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1017
timestamp 1636968456
transform 1 0 94668 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_1029
timestamp 1
transform 1 0 95772 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1035
timestamp 1
transform 1 0 96324 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1037
timestamp 1636968456
transform 1 0 96508 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1049
timestamp 1636968456
transform 1 0 97612 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1061
timestamp 1636968456
transform 1 0 98716 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1073
timestamp 1636968456
transform 1 0 99820 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_1085
timestamp 1
transform 1 0 100924 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1091
timestamp 1
transform 1 0 101476 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1093
timestamp 1636968456
transform 1 0 101660 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1105
timestamp 1636968456
transform 1 0 102764 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1117
timestamp 1636968456
transform 1 0 103868 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1129
timestamp 1636968456
transform 1 0 104972 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_1141
timestamp 1
transform 1 0 106076 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1147
timestamp 1
transform 1 0 106628 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1149
timestamp 1636968456
transform 1 0 106812 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_1161
timestamp 1
transform 1 0 107916 0 1 76160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_137_11
timestamp 1636968456
transform 1 0 2116 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_23
timestamp 1636968456
transform 1 0 3220 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_35
timestamp 1636968456
transform 1 0 4324 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_47
timestamp 1
transform 1 0 5428 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_57
timestamp 1636968456
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_69
timestamp 1636968456
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_81
timestamp 1636968456
transform 1 0 8556 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_93
timestamp 1636968456
transform 1 0 9660 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_105
timestamp 1
transform 1 0 10764 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_111
timestamp 1
transform 1 0 11316 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_113
timestamp 1636968456
transform 1 0 11500 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_125
timestamp 1636968456
transform 1 0 12604 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_137
timestamp 1636968456
transform 1 0 13708 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_149
timestamp 1636968456
transform 1 0 14812 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_161
timestamp 1
transform 1 0 15916 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_167
timestamp 1
transform 1 0 16468 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_169
timestamp 1636968456
transform 1 0 16652 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_181
timestamp 1636968456
transform 1 0 17756 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_193
timestamp 1636968456
transform 1 0 18860 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_205
timestamp 1636968456
transform 1 0 19964 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_217
timestamp 1
transform 1 0 21068 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_223
timestamp 1
transform 1 0 21620 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_137_225
timestamp 1
transform 1 0 21804 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_137_233
timestamp 1
transform 1 0 22540 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_137_281
timestamp 1
transform 1 0 26956 0 -1 77248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_137_292
timestamp 1636968456
transform 1 0 27968 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_304
timestamp 1636968456
transform 1 0 29072 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_321
timestamp 1636968456
transform 1 0 30636 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_137_333
timestamp 1
transform 1 0 31740 0 -1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_137_337
timestamp 1636968456
transform 1 0 32108 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_349
timestamp 1636968456
transform 1 0 33212 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_361
timestamp 1636968456
transform 1 0 34316 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_373
timestamp 1636968456
transform 1 0 35420 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_385
timestamp 1
transform 1 0 36524 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_391
timestamp 1
transform 1 0 37076 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_393
timestamp 1636968456
transform 1 0 37260 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_405
timestamp 1636968456
transform 1 0 38364 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_417
timestamp 1636968456
transform 1 0 39468 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_429
timestamp 1636968456
transform 1 0 40572 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_441
timestamp 1
transform 1 0 41676 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_447
timestamp 1
transform 1 0 42228 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_449
timestamp 1636968456
transform 1 0 42412 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_461
timestamp 1636968456
transform 1 0 43516 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_473
timestamp 1636968456
transform 1 0 44620 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_485
timestamp 1636968456
transform 1 0 45724 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_497
timestamp 1
transform 1 0 46828 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_503
timestamp 1
transform 1 0 47380 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_505
timestamp 1636968456
transform 1 0 47564 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_517
timestamp 1636968456
transform 1 0 48668 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_529
timestamp 1636968456
transform 1 0 49772 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_541
timestamp 1636968456
transform 1 0 50876 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_553
timestamp 1
transform 1 0 51980 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_559
timestamp 1
transform 1 0 52532 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_561
timestamp 1636968456
transform 1 0 52716 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_573
timestamp 1636968456
transform 1 0 53820 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_585
timestamp 1636968456
transform 1 0 54924 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_597
timestamp 1636968456
transform 1 0 56028 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_609
timestamp 1
transform 1 0 57132 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_615
timestamp 1
transform 1 0 57684 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_617
timestamp 1636968456
transform 1 0 57868 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_629
timestamp 1636968456
transform 1 0 58972 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_641
timestamp 1636968456
transform 1 0 60076 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_653
timestamp 1636968456
transform 1 0 61180 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_665
timestamp 1
transform 1 0 62284 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_671
timestamp 1
transform 1 0 62836 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_673
timestamp 1636968456
transform 1 0 63020 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_685
timestamp 1636968456
transform 1 0 64124 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_697
timestamp 1636968456
transform 1 0 65228 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_709
timestamp 1636968456
transform 1 0 66332 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_721
timestamp 1
transform 1 0 67436 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_727
timestamp 1
transform 1 0 67988 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_137_729
timestamp 1
transform 1 0 68172 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_137_737
timestamp 1
transform 1 0 68908 0 -1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_137_744
timestamp 1636968456
transform 1 0 69552 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_756
timestamp 1636968456
transform 1 0 70656 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_768
timestamp 1636968456
transform 1 0 71760 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_780
timestamp 1
transform 1 0 72864 0 -1 77248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_137_785
timestamp 1636968456
transform 1 0 73324 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_797
timestamp 1636968456
transform 1 0 74428 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_813
timestamp 1636968456
transform 1 0 75900 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_825
timestamp 1636968456
transform 1 0 77004 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_137_837
timestamp 1
transform 1 0 78108 0 -1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_137_841
timestamp 1636968456
transform 1 0 78476 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_853
timestamp 1636968456
transform 1 0 79580 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_865
timestamp 1
transform 1 0 80684 0 -1 77248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_137_878
timestamp 1636968456
transform 1 0 81880 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_890
timestamp 1
transform 1 0 82984 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_137_897
timestamp 1
transform 1 0 83628 0 -1 77248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_137_905
timestamp 1636968456
transform 1 0 84364 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_137_917
timestamp 1
transform 1 0 85468 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_137_957
timestamp 1
transform 1 0 89148 0 -1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_137_989
timestamp 1636968456
transform 1 0 92092 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_1001
timestamp 1
transform 1 0 93196 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_1007
timestamp 1
transform 1 0 93748 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1009
timestamp 1636968456
transform 1 0 93932 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1021
timestamp 1636968456
transform 1 0 95036 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1033
timestamp 1636968456
transform 1 0 96140 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1045
timestamp 1636968456
transform 1 0 97244 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_1057
timestamp 1
transform 1 0 98348 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_1063
timestamp 1
transform 1 0 98900 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1065
timestamp 1636968456
transform 1 0 99084 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1077
timestamp 1636968456
transform 1 0 100188 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1089
timestamp 1636968456
transform 1 0 101292 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1101
timestamp 1636968456
transform 1 0 102396 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_1113
timestamp 1
transform 1 0 103500 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_1119
timestamp 1
transform 1 0 104052 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1121
timestamp 1636968456
transform 1 0 104236 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1133
timestamp 1636968456
transform 1 0 105340 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1145
timestamp 1636968456
transform 1 0 106444 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_1157
timestamp 1
transform 1 0 107548 0 -1 77248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_138_3
timestamp 1636968456
transform 1 0 1380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_15
timestamp 1636968456
transform 1 0 2484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 1
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_29
timestamp 1636968456
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_41
timestamp 1636968456
transform 1 0 4876 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_53
timestamp 1
transform 1 0 5980 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_57
timestamp 1636968456
transform 1 0 6348 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_69
timestamp 1636968456
transform 1 0 7452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1
transform 1 0 8556 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_85
timestamp 1636968456
transform 1 0 8924 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_97
timestamp 1636968456
transform 1 0 10028 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_109
timestamp 1
transform 1 0 11132 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_113
timestamp 1636968456
transform 1 0 11500 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_125
timestamp 1636968456
transform 1 0 12604 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_137
timestamp 1
transform 1 0 13708 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_141
timestamp 1636968456
transform 1 0 14076 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_153
timestamp 1
transform 1 0 15180 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_138_161
timestamp 1
transform 1 0 15916 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_138_165
timestamp 1
transform 1 0 16284 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_169
timestamp 1636968456
transform 1 0 16652 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_181
timestamp 1636968456
transform 1 0 17756 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_193
timestamp 1
transform 1 0 18860 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_197
timestamp 1
transform 1 0 19228 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_223
timestamp 1
transform 1 0 21620 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_138_227
timestamp 1
transform 1 0 21988 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_138_255
timestamp 1
transform 1 0 24564 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_281
timestamp 1
transform 1 0 26956 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_138_290
timestamp 1
transform 1 0 27784 0 1 77248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_138_296
timestamp 1636968456
transform 1 0 28336 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_311
timestamp 1
transform 1 0 29716 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_138_321
timestamp 1
transform 1 0 30636 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_335
timestamp 1
transform 1 0 31924 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_356
timestamp 1
transform 1 0 33856 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_138_361
timestamp 1
transform 1 0 34316 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_138_382
timestamp 1
transform 1 0 36248 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_138_385
timestamp 1
transform 1 0 36524 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_389
timestamp 1
transform 1 0 36892 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_410
timestamp 1
transform 1 0 38824 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_138_438
timestamp 1
transform 1 0 41400 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_138_466
timestamp 1
transform 1 0 43976 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_138_474
timestamp 1
transform 1 0 44712 0 1 77248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_138_477
timestamp 1636968456
transform 1 0 44988 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_489
timestamp 1636968456
transform 1 0 46092 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_501
timestamp 1
transform 1 0 47196 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_505
timestamp 1636968456
transform 1 0 47564 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_517
timestamp 1636968456
transform 1 0 48668 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_529
timestamp 1
transform 1 0 49772 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_533
timestamp 1636968456
transform 1 0 50140 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_545
timestamp 1636968456
transform 1 0 51244 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_557
timestamp 1
transform 1 0 52348 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_561
timestamp 1636968456
transform 1 0 52716 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_573
timestamp 1636968456
transform 1 0 53820 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_585
timestamp 1
transform 1 0 54924 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_589
timestamp 1636968456
transform 1 0 55292 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_601
timestamp 1636968456
transform 1 0 56396 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_613
timestamp 1
transform 1 0 57500 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_617
timestamp 1636968456
transform 1 0 57868 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_629
timestamp 1636968456
transform 1 0 58972 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_641
timestamp 1
transform 1 0 60076 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_662
timestamp 1
transform 1 0 62008 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_666
timestamp 1
transform 1 0 62376 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_671
timestamp 1
transform 1 0 62836 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_686
timestamp 1
transform 1 0 64216 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_138_694
timestamp 1
transform 1 0 64952 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_699
timestamp 1
transform 1 0 65412 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_714
timestamp 1
transform 1 0 66792 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_138_722
timestamp 1
transform 1 0 67528 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_727
timestamp 1
transform 1 0 67988 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_742
timestamp 1
transform 1 0 69368 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_757
timestamp 1
transform 1 0 70748 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_773
timestamp 1
transform 1 0 72220 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_781
timestamp 1
transform 1 0 72956 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_138_822
timestamp 1
transform 1 0 76728 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_830
timestamp 1
transform 1 0 77464 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_138_839
timestamp 1
transform 1 0 78292 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_138_850
timestamp 1
transform 1 0 79304 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_138_869
timestamp 1
transform 1 0 81052 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_895
timestamp 1
transform 1 0 83444 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_902
timestamp 1
transform 1 0 84088 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_923
timestamp 1
transform 1 0 86020 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_938
timestamp 1636968456
transform 1 0 87400 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_138_950
timestamp 1
transform 1 0 88504 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_138_977
timestamp 1
transform 1 0 90988 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_1003
timestamp 1
transform 1 0 93380 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_1007
timestamp 1
transform 1 0 93748 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_138_1031
timestamp 1
transform 1 0 95956 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_1035
timestamp 1
transform 1 0 96324 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1037
timestamp 1636968456
transform 1 0 96508 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1049
timestamp 1636968456
transform 1 0 97612 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_1061
timestamp 1
transform 1 0 98716 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1065
timestamp 1636968456
transform 1 0 99084 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1077
timestamp 1636968456
transform 1 0 100188 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_1089
timestamp 1
transform 1 0 101292 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1093
timestamp 1636968456
transform 1 0 101660 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1105
timestamp 1636968456
transform 1 0 102764 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_1117
timestamp 1
transform 1 0 103868 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1121
timestamp 1636968456
transform 1 0 104236 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1133
timestamp 1636968456
transform 1 0 105340 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_1145
timestamp 1
transform 1 0 106444 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1149
timestamp 1636968456
transform 1 0 106812 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_1161
timestamp 1
transform 1 0 107916 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_1167
timestamp 1
transform 1 0 108468 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_11
timestamp 1636968456
transform 1 0 2116 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_23
timestamp 1636968456
transform 1 0 3220 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_35
timestamp 1636968456
transform 1 0 4324 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_47
timestamp 1
transform 1 0 5428 0 -1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_139_55
timestamp 1
transform 1 0 6164 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_57
timestamp 1636968456
transform 1 0 6348 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_139_69
timestamp 1
transform 1 0 7452 0 -1 78336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1122
timestamp 1636968456
transform 1 0 104328 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1134
timestamp 1636968456
transform 1 0 105432 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1146
timestamp 1636968456
transform 1 0 106536 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_139_1158
timestamp 1
transform 1 0 107640 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_139_1162
timestamp 1
transform 1 0 108008 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_11
timestamp 1636968456
transform 1 0 2116 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_140_23
timestamp 1
transform 1 0 3220 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_140_27
timestamp 1
transform 1 0 3588 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_29
timestamp 1636968456
transform 1 0 3772 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_41
timestamp 1636968456
transform 1 0 4876 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_53
timestamp 1636968456
transform 1 0 5980 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_65
timestamp 1
transform 1 0 7084 0 1 78336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1122
timestamp 1636968456
transform 1 0 104328 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1134
timestamp 1636968456
transform 1 0 105432 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_140_1146
timestamp 1
transform 1 0 106536 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1148
timestamp 1636968456
transform 1 0 106720 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_140_1160
timestamp 1
transform 1 0 107824 0 1 78336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_141_11
timestamp 1636968456
transform 1 0 2116 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_23
timestamp 1636968456
transform 1 0 3220 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_35
timestamp 1636968456
transform 1 0 4324 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_141_47
timestamp 1
transform 1 0 5428 0 -1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_141_55
timestamp 1
transform 1 0 6164 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_57
timestamp 1636968456
transform 1 0 6348 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_141_69
timestamp 1
transform 1 0 7452 0 -1 79424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1122
timestamp 1636968456
transform 1 0 104328 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1134
timestamp 1636968456
transform 1 0 105432 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1146
timestamp 1636968456
transform 1 0 106536 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_141_1158
timestamp 1
transform 1 0 107640 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_141_1162
timestamp 1
transform 1 0 108008 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_11
timestamp 1636968456
transform 1 0 2116 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_142_23
timestamp 1
transform 1 0 3220 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_142_27
timestamp 1
transform 1 0 3588 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_29
timestamp 1636968456
transform 1 0 3772 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_41
timestamp 1636968456
transform 1 0 4876 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_53
timestamp 1636968456
transform 1 0 5980 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_65
timestamp 1
transform 1 0 7084 0 1 79424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1122
timestamp 1636968456
transform 1 0 104328 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1134
timestamp 1636968456
transform 1 0 105432 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_1146
timestamp 1
transform 1 0 106536 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1148
timestamp 1636968456
transform 1 0 106720 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_142_1160
timestamp 1
transform 1 0 107824 0 1 79424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_143_5
timestamp 1636968456
transform 1 0 1564 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_17
timestamp 1636968456
transform 1 0 2668 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_29
timestamp 1636968456
transform 1 0 3772 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_41
timestamp 1636968456
transform 1 0 4876 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_143_53
timestamp 1
transform 1 0 5980 0 -1 80512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_143_57
timestamp 1636968456
transform 1 0 6348 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_143_69
timestamp 1
transform 1 0 7452 0 -1 80512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1122
timestamp 1636968456
transform 1 0 104328 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1134
timestamp 1636968456
transform 1 0 105432 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1146
timestamp 1636968456
transform 1 0 106536 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_143_1158
timestamp 1
transform 1 0 107640 0 -1 80512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_143_1166
timestamp 1
transform 1 0 108376 0 -1 80512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_144_15
timestamp 1636968456
transform 1 0 2484 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_27
timestamp 1
transform 1 0 3588 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_29
timestamp 1636968456
transform 1 0 3772 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_41
timestamp 1636968456
transform 1 0 4876 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_53
timestamp 1636968456
transform 1 0 5980 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_65
timestamp 1
transform 1 0 7084 0 1 80512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1122
timestamp 1636968456
transform 1 0 104328 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1134
timestamp 1636968456
transform 1 0 105432 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_1146
timestamp 1
transform 1 0 106536 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1148
timestamp 1636968456
transform 1 0 106720 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_144_1160
timestamp 1
transform 1 0 107824 0 1 80512
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_145_11
timestamp 1636968456
transform 1 0 2116 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_23
timestamp 1636968456
transform 1 0 3220 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_35
timestamp 1636968456
transform 1 0 4324 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_145_47
timestamp 1
transform 1 0 5428 0 -1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_145_55
timestamp 1
transform 1 0 6164 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_57
timestamp 1636968456
transform 1 0 6348 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_145_69
timestamp 1
transform 1 0 7452 0 -1 81600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1122
timestamp 1636968456
transform 1 0 104328 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1134
timestamp 1636968456
transform 1 0 105432 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1146
timestamp 1636968456
transform 1 0 106536 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_145_1158
timestamp 1
transform 1 0 107640 0 -1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_145_1166
timestamp 1
transform 1 0 108376 0 -1 81600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_146_11
timestamp 1636968456
transform 1 0 2116 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_146_23
timestamp 1
transform 1 0 3220 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_27
timestamp 1
transform 1 0 3588 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_29
timestamp 1636968456
transform 1 0 3772 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_41
timestamp 1636968456
transform 1 0 4876 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_53
timestamp 1636968456
transform 1 0 5980 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_65
timestamp 1
transform 1 0 7084 0 1 81600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1122
timestamp 1636968456
transform 1 0 104328 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1134
timestamp 1636968456
transform 1 0 105432 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_1146
timestamp 1
transform 1 0 106536 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1148
timestamp 1636968456
transform 1 0 106720 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_1160
timestamp 1
transform 1 0 107824 0 1 81600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_147_11
timestamp 1636968456
transform 1 0 2116 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_23
timestamp 1636968456
transform 1 0 3220 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_35
timestamp 1636968456
transform 1 0 4324 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_47
timestamp 1
transform 1 0 5428 0 -1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_147_55
timestamp 1
transform 1 0 6164 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_57
timestamp 1636968456
transform 1 0 6348 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_147_69
timestamp 1
transform 1 0 7452 0 -1 82688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1122
timestamp 1636968456
transform 1 0 104328 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1134
timestamp 1636968456
transform 1 0 105432 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1146
timestamp 1636968456
transform 1 0 106536 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_1158
timestamp 1
transform 1 0 107640 0 -1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_147_1166
timestamp 1
transform 1 0 108376 0 -1 82688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_148_3
timestamp 1636968456
transform 1 0 1380 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_15
timestamp 1636968456
transform 1 0 2484 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_27
timestamp 1
transform 1 0 3588 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_29
timestamp 1636968456
transform 1 0 3772 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_41
timestamp 1636968456
transform 1 0 4876 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_53
timestamp 1636968456
transform 1 0 5980 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_65
timestamp 1
transform 1 0 7084 0 1 82688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1122
timestamp 1636968456
transform 1 0 104328 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1134
timestamp 1636968456
transform 1 0 105432 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_1146
timestamp 1
transform 1 0 106536 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1148
timestamp 1636968456
transform 1 0 106720 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_148_1160
timestamp 1
transform 1 0 107824 0 1 82688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_149_11
timestamp 1636968456
transform 1 0 2116 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_23
timestamp 1636968456
transform 1 0 3220 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_35
timestamp 1636968456
transform 1 0 4324 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_47
timestamp 1
transform 1 0 5428 0 -1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_149_55
timestamp 1
transform 1 0 6164 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_57
timestamp 1636968456
transform 1 0 6348 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_149_69
timestamp 1
transform 1 0 7452 0 -1 83776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1122
timestamp 1636968456
transform 1 0 104328 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1134
timestamp 1636968456
transform 1 0 105432 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1146
timestamp 1636968456
transform 1 0 106536 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_1158
timestamp 1
transform 1 0 107640 0 -1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_149_1166
timestamp 1
transform 1 0 108376 0 -1 83776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_150_11
timestamp 1636968456
transform 1 0 2116 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_150_23
timestamp 1
transform 1 0 3220 0 1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_150_27
timestamp 1
transform 1 0 3588 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_29
timestamp 1636968456
transform 1 0 3772 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_41
timestamp 1636968456
transform 1 0 4876 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_53
timestamp 1636968456
transform 1 0 5980 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_65
timestamp 1
transform 1 0 7084 0 1 83776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1122
timestamp 1636968456
transform 1 0 104328 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1134
timestamp 1636968456
transform 1 0 105432 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_1146
timestamp 1
transform 1 0 106536 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1148
timestamp 1636968456
transform 1 0 106720 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_1160
timestamp 1
transform 1 0 107824 0 1 83776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_151_11
timestamp 1636968456
transform 1 0 2116 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_23
timestamp 1636968456
transform 1 0 3220 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_35
timestamp 1636968456
transform 1 0 4324 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_47
timestamp 1
transform 1 0 5428 0 -1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_55
timestamp 1
transform 1 0 6164 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_57
timestamp 1636968456
transform 1 0 6348 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_151_69
timestamp 1
transform 1 0 7452 0 -1 84864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1122
timestamp 1636968456
transform 1 0 104328 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1134
timestamp 1636968456
transform 1 0 105432 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1146
timestamp 1636968456
transform 1 0 106536 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_1158
timestamp 1
transform 1 0 107640 0 -1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_1166
timestamp 1
transform 1 0 108376 0 -1 84864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_152_11
timestamp 1636968456
transform 1 0 2116 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_152_23
timestamp 1
transform 1 0 3220 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_152_27
timestamp 1
transform 1 0 3588 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_29
timestamp 1636968456
transform 1 0 3772 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_41
timestamp 1636968456
transform 1 0 4876 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_53
timestamp 1636968456
transform 1 0 5980 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_65
timestamp 1
transform 1 0 7084 0 1 84864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1122
timestamp 1636968456
transform 1 0 104328 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1134
timestamp 1636968456
transform 1 0 105432 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_152_1146
timestamp 1
transform 1 0 106536 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1148
timestamp 1636968456
transform 1 0 106720 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_1160
timestamp 1
transform 1 0 107824 0 1 84864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_153_3
timestamp 1636968456
transform 1 0 1380 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_15
timestamp 1636968456
transform 1 0 2484 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_27
timestamp 1636968456
transform 1 0 3588 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_39
timestamp 1636968456
transform 1 0 4692 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_153_51
timestamp 1
transform 1 0 5796 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_153_55
timestamp 1
transform 1 0 6164 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_57
timestamp 1636968456
transform 1 0 6348 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_153_69
timestamp 1
transform 1 0 7452 0 -1 85952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1122
timestamp 1636968456
transform 1 0 104328 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1134
timestamp 1636968456
transform 1 0 105432 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1146
timestamp 1636968456
transform 1 0 106536 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_153_1158
timestamp 1
transform 1 0 107640 0 -1 85952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_153_1166
timestamp 1
transform 1 0 108376 0 -1 85952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_154_8
timestamp 1636968456
transform 1 0 1840 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_20
timestamp 1
transform 1 0 2944 0 1 85952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_154_29
timestamp 1636968456
transform 1 0 3772 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_41
timestamp 1636968456
transform 1 0 4876 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_53
timestamp 1636968456
transform 1 0 5980 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_65
timestamp 1
transform 1 0 7084 0 1 85952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1122
timestamp 1636968456
transform 1 0 104328 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1134
timestamp 1636968456
transform 1 0 105432 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_1146
timestamp 1
transform 1 0 106536 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1148
timestamp 1636968456
transform 1 0 106720 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_1160
timestamp 1
transform 1 0 107824 0 1 85952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_155_11
timestamp 1636968456
transform 1 0 2116 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_23
timestamp 1636968456
transform 1 0 3220 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_35
timestamp 1636968456
transform 1 0 4324 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_155_47
timestamp 1
transform 1 0 5428 0 -1 87040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_155_55
timestamp 1
transform 1 0 6164 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_57
timestamp 1636968456
transform 1 0 6348 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_155_69
timestamp 1
transform 1 0 7452 0 -1 87040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1122
timestamp 1636968456
transform 1 0 104328 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1134
timestamp 1636968456
transform 1 0 105432 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1146
timestamp 1636968456
transform 1 0 106536 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_155_1158
timestamp 1
transform 1 0 107640 0 -1 87040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_155_1166
timestamp 1
transform 1 0 108376 0 -1 87040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_156_11
timestamp 1636968456
transform 1 0 2116 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_156_23
timestamp 1
transform 1 0 3220 0 1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_156_27
timestamp 1
transform 1 0 3588 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_29
timestamp 1636968456
transform 1 0 3772 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_41
timestamp 1636968456
transform 1 0 4876 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_53
timestamp 1636968456
transform 1 0 5980 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_65
timestamp 1
transform 1 0 7084 0 1 87040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1122
timestamp 1636968456
transform 1 0 104328 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1134
timestamp 1636968456
transform 1 0 105432 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_156_1146
timestamp 1
transform 1 0 106536 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1148
timestamp 1636968456
transform 1 0 106720 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_156_1160
timestamp 1
transform 1 0 107824 0 1 87040
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_157_11
timestamp 1636968456
transform 1 0 2116 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_23
timestamp 1636968456
transform 1 0 3220 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_35
timestamp 1636968456
transform 1 0 4324 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_47
timestamp 1
transform 1 0 5428 0 -1 88128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_157_55
timestamp 1
transform 1 0 6164 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_57
timestamp 1636968456
transform 1 0 6348 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_157_69
timestamp 1
transform 1 0 7452 0 -1 88128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1122
timestamp 1636968456
transform 1 0 104328 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1134
timestamp 1636968456
transform 1 0 105432 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1146
timestamp 1636968456
transform 1 0 106536 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_1158
timestamp 1
transform 1 0 107640 0 -1 88128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_157_1166
timestamp 1
transform 1 0 108376 0 -1 88128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_158_3
timestamp 1636968456
transform 1 0 1380 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_15
timestamp 1636968456
transform 1 0 2484 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_27
timestamp 1
transform 1 0 3588 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_29
timestamp 1636968456
transform 1 0 3772 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_41
timestamp 1636968456
transform 1 0 4876 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_53
timestamp 1636968456
transform 1 0 5980 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_65
timestamp 1
transform 1 0 7084 0 1 88128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1122
timestamp 1636968456
transform 1 0 104328 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1134
timestamp 1636968456
transform 1 0 105432 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_1146
timestamp 1
transform 1 0 106536 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1148
timestamp 1636968456
transform 1 0 106720 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_158_1160
timestamp 1
transform 1 0 107824 0 1 88128
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_159_11
timestamp 1636968456
transform 1 0 2116 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_23
timestamp 1636968456
transform 1 0 3220 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_35
timestamp 1636968456
transform 1 0 4324 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_47
timestamp 1
transform 1 0 5428 0 -1 89216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_159_55
timestamp 1
transform 1 0 6164 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_57
timestamp 1636968456
transform 1 0 6348 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_159_69
timestamp 1
transform 1 0 7452 0 -1 89216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1122
timestamp 1636968456
transform 1 0 104328 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1134
timestamp 1636968456
transform 1 0 105432 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1146
timestamp 1636968456
transform 1 0 106536 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_1158
timestamp 1
transform 1 0 107640 0 -1 89216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_159_1166
timestamp 1
transform 1 0 108376 0 -1 89216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_160_3
timestamp 1636968456
transform 1 0 1380 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_15
timestamp 1636968456
transform 1 0 2484 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_27
timestamp 1
transform 1 0 3588 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_29
timestamp 1636968456
transform 1 0 3772 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_41
timestamp 1636968456
transform 1 0 4876 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_53
timestamp 1636968456
transform 1 0 5980 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_65
timestamp 1
transform 1 0 7084 0 1 89216
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1122
timestamp 1636968456
transform 1 0 104328 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1134
timestamp 1636968456
transform 1 0 105432 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_1146
timestamp 1
transform 1 0 106536 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1148
timestamp 1636968456
transform 1 0 106720 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_160_1160
timestamp 1
transform 1 0 107824 0 1 89216
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_161_3
timestamp 1636968456
transform 1 0 1380 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_15
timestamp 1636968456
transform 1 0 2484 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_27
timestamp 1636968456
transform 1 0 3588 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_39
timestamp 1636968456
transform 1 0 4692 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_161_51
timestamp 1
transform 1 0 5796 0 -1 90304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_161_55
timestamp 1
transform 1 0 6164 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_57
timestamp 1636968456
transform 1 0 6348 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_161_69
timestamp 1
transform 1 0 7452 0 -1 90304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1122
timestamp 1636968456
transform 1 0 104328 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1134
timestamp 1636968456
transform 1 0 105432 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1146
timestamp 1636968456
transform 1 0 106536 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_1158
timestamp 1
transform 1 0 107640 0 -1 90304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_161_1166
timestamp 1
transform 1 0 108376 0 -1 90304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_162_3
timestamp 1636968456
transform 1 0 1380 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_15
timestamp 1636968456
transform 1 0 2484 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_27
timestamp 1
transform 1 0 3588 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_29
timestamp 1636968456
transform 1 0 3772 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_41
timestamp 1636968456
transform 1 0 4876 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_53
timestamp 1636968456
transform 1 0 5980 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_65
timestamp 1
transform 1 0 7084 0 1 90304
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1124
timestamp 1636968456
transform 1 0 104512 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_162_1136
timestamp 1
transform 1 0 105616 0 1 90304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_162_1144
timestamp 1
transform 1 0 106352 0 1 90304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1148
timestamp 1636968456
transform 1 0 106720 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_162_1160
timestamp 1
transform 1 0 107824 0 1 90304
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_163_3
timestamp 1636968456
transform 1 0 1380 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_15
timestamp 1636968456
transform 1 0 2484 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_27
timestamp 1636968456
transform 1 0 3588 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_39
timestamp 1636968456
transform 1 0 4692 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_163_51
timestamp 1
transform 1 0 5796 0 -1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_163_55
timestamp 1
transform 1 0 6164 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_57
timestamp 1636968456
transform 1 0 6348 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_163_69
timestamp 1
transform 1 0 7452 0 -1 91392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1144
timestamp 1636968456
transform 1 0 106352 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1156
timestamp 1636968456
transform 1 0 107456 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_3
timestamp 1636968456
transform 1 0 1380 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_15
timestamp 1636968456
transform 1 0 2484 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_27
timestamp 1
transform 1 0 3588 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_29
timestamp 1636968456
transform 1 0 3772 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_41
timestamp 1636968456
transform 1 0 4876 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_53
timestamp 1636968456
transform 1 0 5980 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_65
timestamp 1
transform 1 0 7084 0 1 91392
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1122
timestamp 1636968456
transform 1 0 104328 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1134
timestamp 1636968456
transform 1 0 105432 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_1146
timestamp 1
transform 1 0 106536 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1148
timestamp 1636968456
transform 1 0 106720 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_164_1160
timestamp 1
transform 1 0 107824 0 1 91392
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_165_3
timestamp 1636968456
transform 1 0 1380 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_15
timestamp 1636968456
transform 1 0 2484 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_27
timestamp 1636968456
transform 1 0 3588 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_39
timestamp 1636968456
transform 1 0 4692 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_165_51
timestamp 1
transform 1 0 5796 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_165_55
timestamp 1
transform 1 0 6164 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_57
timestamp 1636968456
transform 1 0 6348 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_165_69
timestamp 1
transform 1 0 7452 0 -1 92480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1122
timestamp 1636968456
transform 1 0 104328 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1134
timestamp 1636968456
transform 1 0 105432 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1146
timestamp 1636968456
transform 1 0 106536 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_1158
timestamp 1
transform 1 0 107640 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_165_1166
timestamp 1
transform 1 0 108376 0 -1 92480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_166_3
timestamp 1636968456
transform 1 0 1380 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_15
timestamp 1636968456
transform 1 0 2484 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_27
timestamp 1
transform 1 0 3588 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_29
timestamp 1636968456
transform 1 0 3772 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_41
timestamp 1636968456
transform 1 0 4876 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_53
timestamp 1636968456
transform 1 0 5980 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_65
timestamp 1
transform 1 0 7084 0 1 92480
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1124
timestamp 1636968456
transform 1 0 104512 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_1136
timestamp 1
transform 1 0 105616 0 1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_166_1144
timestamp 1
transform 1 0 106352 0 1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1148
timestamp 1636968456
transform 1 0 106720 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_1160
timestamp 1
transform 1 0 107824 0 1 92480
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_167_3
timestamp 1636968456
transform 1 0 1380 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_15
timestamp 1636968456
transform 1 0 2484 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_27
timestamp 1636968456
transform 1 0 3588 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_39
timestamp 1636968456
transform 1 0 4692 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_167_51
timestamp 1
transform 1 0 5796 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_55
timestamp 1
transform 1 0 6164 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_57
timestamp 1636968456
transform 1 0 6348 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_167_69
timestamp 1
transform 1 0 7452 0 -1 93568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1122
timestamp 1636968456
transform 1 0 104328 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1134
timestamp 1636968456
transform 1 0 105432 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1146
timestamp 1636968456
transform 1 0 106536 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_1158
timestamp 1
transform 1 0 107640 0 -1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_167_1166
timestamp 1
transform 1 0 108376 0 -1 93568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_168_3
timestamp 1636968456
transform 1 0 1380 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_15
timestamp 1636968456
transform 1 0 2484 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_27
timestamp 1
transform 1 0 3588 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_29
timestamp 1636968456
transform 1 0 3772 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_41
timestamp 1636968456
transform 1 0 4876 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_53
timestamp 1636968456
transform 1 0 5980 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_65
timestamp 1
transform 1 0 7084 0 1 93568
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1124
timestamp 1636968456
transform 1 0 104512 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_168_1136
timestamp 1
transform 1 0 105616 0 1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_168_1144
timestamp 1
transform 1 0 106352 0 1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1148
timestamp 1636968456
transform 1 0 106720 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_168_1160
timestamp 1
transform 1 0 107824 0 1 93568
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_169_3
timestamp 1636968456
transform 1 0 1380 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_15
timestamp 1636968456
transform 1 0 2484 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_27
timestamp 1636968456
transform 1 0 3588 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_39
timestamp 1636968456
transform 1 0 4692 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_169_51
timestamp 1
transform 1 0 5796 0 -1 94656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_169_55
timestamp 1
transform 1 0 6164 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_57
timestamp 1636968456
transform 1 0 6348 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_169_69
timestamp 1
transform 1 0 7452 0 -1 94656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1122
timestamp 1636968456
transform 1 0 104328 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1134
timestamp 1636968456
transform 1 0 105432 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1146
timestamp 1636968456
transform 1 0 106536 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_169_1158
timestamp 1
transform 1 0 107640 0 -1 94656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_169_1166
timestamp 1
transform 1 0 108376 0 -1 94656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_170_3
timestamp 1636968456
transform 1 0 1380 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_15
timestamp 1636968456
transform 1 0 2484 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_27
timestamp 1
transform 1 0 3588 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_29
timestamp 1636968456
transform 1 0 3772 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_41
timestamp 1636968456
transform 1 0 4876 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_53
timestamp 1636968456
transform 1 0 5980 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_65
timestamp 1
transform 1 0 7084 0 1 94656
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1122
timestamp 1636968456
transform 1 0 104328 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1134
timestamp 1636968456
transform 1 0 105432 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_1146
timestamp 1
transform 1 0 106536 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1148
timestamp 1636968456
transform 1 0 106720 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_170_1160
timestamp 1
transform 1 0 107824 0 1 94656
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_171_3
timestamp 1636968456
transform 1 0 1380 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_15
timestamp 1636968456
transform 1 0 2484 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_27
timestamp 1636968456
transform 1 0 3588 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_39
timestamp 1636968456
transform 1 0 4692 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_171_51
timestamp 1
transform 1 0 5796 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_171_55
timestamp 1
transform 1 0 6164 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_57
timestamp 1636968456
transform 1 0 6348 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_171_69
timestamp 1
transform 1 0 7452 0 -1 95744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1124
timestamp 1636968456
transform 1 0 104512 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1136
timestamp 1636968456
transform 1 0 105616 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1148
timestamp 1636968456
transform 1 0 106720 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_1160
timestamp 1
transform 1 0 107824 0 -1 95744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_172_3
timestamp 1636968456
transform 1 0 1380 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_15
timestamp 1636968456
transform 1 0 2484 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_172_27
timestamp 1
transform 1 0 3588 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_29
timestamp 1636968456
transform 1 0 3772 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_41
timestamp 1636968456
transform 1 0 4876 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_53
timestamp 1636968456
transform 1 0 5980 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_65
timestamp 1
transform 1 0 7084 0 1 95744
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1122
timestamp 1636968456
transform 1 0 104328 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1134
timestamp 1636968456
transform 1 0 105432 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_172_1146
timestamp 1
transform 1 0 106536 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1148
timestamp 1636968456
transform 1 0 106720 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_1160
timestamp 1
transform 1 0 107824 0 1 95744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_173_3
timestamp 1636968456
transform 1 0 1380 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_15
timestamp 1636968456
transform 1 0 2484 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_27
timestamp 1636968456
transform 1 0 3588 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_39
timestamp 1636968456
transform 1 0 4692 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_173_51
timestamp 1
transform 1 0 5796 0 -1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_173_55
timestamp 1
transform 1 0 6164 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_57
timestamp 1636968456
transform 1 0 6348 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_173_69
timestamp 1
transform 1 0 7452 0 -1 96832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1122
timestamp 1636968456
transform 1 0 104328 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1134
timestamp 1636968456
transform 1 0 105432 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1146
timestamp 1636968456
transform 1 0 106536 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_1158
timestamp 1
transform 1 0 107640 0 -1 96832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_173_1166
timestamp 1
transform 1 0 108376 0 -1 96832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_174_3
timestamp 1636968456
transform 1 0 1380 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_15
timestamp 1636968456
transform 1 0 2484 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_174_27
timestamp 1
transform 1 0 3588 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_29
timestamp 1636968456
transform 1 0 3772 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_41
timestamp 1636968456
transform 1 0 4876 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_53
timestamp 1636968456
transform 1 0 5980 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_65
timestamp 1
transform 1 0 7084 0 1 96832
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1122
timestamp 1636968456
transform 1 0 104328 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1134
timestamp 1636968456
transform 1 0 105432 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_174_1146
timestamp 1
transform 1 0 106536 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1148
timestamp 1636968456
transform 1 0 106720 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_174_1160
timestamp 1
transform 1 0 107824 0 1 96832
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_175_3
timestamp 1636968456
transform 1 0 1380 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_15
timestamp 1636968456
transform 1 0 2484 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_27
timestamp 1636968456
transform 1 0 3588 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_39
timestamp 1636968456
transform 1 0 4692 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_175_51
timestamp 1
transform 1 0 5796 0 -1 97920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_175_55
timestamp 1
transform 1 0 6164 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_57
timestamp 1636968456
transform 1 0 6348 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_175_69
timestamp 1
transform 1 0 7452 0 -1 97920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1122
timestamp 1636968456
transform 1 0 104328 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1134
timestamp 1636968456
transform 1 0 105432 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1146
timestamp 1636968456
transform 1 0 106536 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_175_1158
timestamp 1
transform 1 0 107640 0 -1 97920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_175_1166
timestamp 1
transform 1 0 108376 0 -1 97920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_176_3
timestamp 1636968456
transform 1 0 1380 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_15
timestamp 1636968456
transform 1 0 2484 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_176_27
timestamp 1
transform 1 0 3588 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_29
timestamp 1636968456
transform 1 0 3772 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_41
timestamp 1636968456
transform 1 0 4876 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_53
timestamp 1636968456
transform 1 0 5980 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_65
timestamp 1
transform 1 0 7084 0 1 97920
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1122
timestamp 1636968456
transform 1 0 104328 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1134
timestamp 1636968456
transform 1 0 105432 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_176_1146
timestamp 1
transform 1 0 106536 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1148
timestamp 1636968456
transform 1 0 106720 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_176_1160
timestamp 1
transform 1 0 107824 0 1 97920
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_177_3
timestamp 1636968456
transform 1 0 1380 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_15
timestamp 1636968456
transform 1 0 2484 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_27
timestamp 1636968456
transform 1 0 3588 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_39
timestamp 1636968456
transform 1 0 4692 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_177_51
timestamp 1
transform 1 0 5796 0 -1 99008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_177_55
timestamp 1
transform 1 0 6164 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_57
timestamp 1636968456
transform 1 0 6348 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_177_69
timestamp 1
transform 1 0 7452 0 -1 99008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1122
timestamp 1636968456
transform 1 0 104328 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1134
timestamp 1636968456
transform 1 0 105432 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1146
timestamp 1636968456
transform 1 0 106536 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_177_1158
timestamp 1
transform 1 0 107640 0 -1 99008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_177_1166
timestamp 1
transform 1 0 108376 0 -1 99008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_178_3
timestamp 1636968456
transform 1 0 1380 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_15
timestamp 1636968456
transform 1 0 2484 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_178_27
timestamp 1
transform 1 0 3588 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_29
timestamp 1636968456
transform 1 0 3772 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_41
timestamp 1636968456
transform 1 0 4876 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_53
timestamp 1636968456
transform 1 0 5980 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_65
timestamp 1
transform 1 0 7084 0 1 99008
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1122
timestamp 1636968456
transform 1 0 104328 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1134
timestamp 1636968456
transform 1 0 105432 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_178_1146
timestamp 1
transform 1 0 106536 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1148
timestamp 1636968456
transform 1 0 106720 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_178_1160
timestamp 1
transform 1 0 107824 0 1 99008
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_179_3
timestamp 1636968456
transform 1 0 1380 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_15
timestamp 1636968456
transform 1 0 2484 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_27
timestamp 1636968456
transform 1 0 3588 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_39
timestamp 1636968456
transform 1 0 4692 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_179_51
timestamp 1
transform 1 0 5796 0 -1 100096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_179_55
timestamp 1
transform 1 0 6164 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_57
timestamp 1636968456
transform 1 0 6348 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_179_69
timestamp 1
transform 1 0 7452 0 -1 100096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1122
timestamp 1636968456
transform 1 0 104328 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1134
timestamp 1636968456
transform 1 0 105432 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1146
timestamp 1636968456
transform 1 0 106536 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_1158
timestamp 1
transform 1 0 107640 0 -1 100096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_179_1166
timestamp 1
transform 1 0 108376 0 -1 100096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_180_3
timestamp 1636968456
transform 1 0 1380 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_15
timestamp 1636968456
transform 1 0 2484 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_180_27
timestamp 1
transform 1 0 3588 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_29
timestamp 1636968456
transform 1 0 3772 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_41
timestamp 1636968456
transform 1 0 4876 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_53
timestamp 1636968456
transform 1 0 5980 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_65
timestamp 1
transform 1 0 7084 0 1 100096
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1122
timestamp 1636968456
transform 1 0 104328 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1134
timestamp 1636968456
transform 1 0 105432 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_180_1146
timestamp 1
transform 1 0 106536 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1148
timestamp 1636968456
transform 1 0 106720 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_180_1160
timestamp 1
transform 1 0 107824 0 1 100096
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_181_3
timestamp 1636968456
transform 1 0 1380 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_15
timestamp 1636968456
transform 1 0 2484 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_27
timestamp 1636968456
transform 1 0 3588 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_39
timestamp 1636968456
transform 1 0 4692 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_181_51
timestamp 1
transform 1 0 5796 0 -1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_181_55
timestamp 1
transform 1 0 6164 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_57
timestamp 1636968456
transform 1 0 6348 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_181_69
timestamp 1
transform 1 0 7452 0 -1 101184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1122
timestamp 1636968456
transform 1 0 104328 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1134
timestamp 1636968456
transform 1 0 105432 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1146
timestamp 1636968456
transform 1 0 106536 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_181_1158
timestamp 1
transform 1 0 107640 0 -1 101184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_181_1166
timestamp 1
transform 1 0 108376 0 -1 101184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_182_3
timestamp 1636968456
transform 1 0 1380 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_15
timestamp 1636968456
transform 1 0 2484 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_182_27
timestamp 1
transform 1 0 3588 0 1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_182_29
timestamp 1636968456
transform 1 0 3772 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_41
timestamp 1636968456
transform 1 0 4876 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_53
timestamp 1636968456
transform 1 0 5980 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_65
timestamp 1
transform 1 0 7084 0 1 101184
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1122
timestamp 1636968456
transform 1 0 104328 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1134
timestamp 1636968456
transform 1 0 105432 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_182_1146
timestamp 1
transform 1 0 106536 0 1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1148
timestamp 1636968456
transform 1 0 106720 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_182_1160
timestamp 1
transform 1 0 107824 0 1 101184
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_183_3
timestamp 1636968456
transform 1 0 1380 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_15
timestamp 1636968456
transform 1 0 2484 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_27
timestamp 1636968456
transform 1 0 3588 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_39
timestamp 1636968456
transform 1 0 4692 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_183_51
timestamp 1
transform 1 0 5796 0 -1 102272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_183_55
timestamp 1
transform 1 0 6164 0 -1 102272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_183_57
timestamp 1636968456
transform 1 0 6348 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_183_69
timestamp 1
transform 1 0 7452 0 -1 102272
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_183_1122
timestamp 1636968456
transform 1 0 104328 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_1134
timestamp 1636968456
transform 1 0 105432 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_1146
timestamp 1636968456
transform 1 0 106536 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_183_1158
timestamp 1
transform 1 0 107640 0 -1 102272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_183_1166
timestamp 1
transform 1 0 108376 0 -1 102272
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_184_3
timestamp 1636968456
transform 1 0 1380 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_15
timestamp 1636968456
transform 1 0 2484 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_184_27
timestamp 1
transform 1 0 3588 0 1 102272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_184_29
timestamp 1636968456
transform 1 0 3772 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_41
timestamp 1636968456
transform 1 0 4876 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_53
timestamp 1636968456
transform 1 0 5980 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_65
timestamp 1
transform 1 0 7084 0 1 102272
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_184_1122
timestamp 1636968456
transform 1 0 104328 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_1134
timestamp 1636968456
transform 1 0 105432 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_184_1146
timestamp 1
transform 1 0 106536 0 1 102272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_184_1148
timestamp 1636968456
transform 1 0 106720 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_184_1160
timestamp 1
transform 1 0 107824 0 1 102272
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_185_3
timestamp 1636968456
transform 1 0 1380 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_15
timestamp 1636968456
transform 1 0 2484 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_27
timestamp 1636968456
transform 1 0 3588 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_39
timestamp 1636968456
transform 1 0 4692 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_185_51
timestamp 1
transform 1 0 5796 0 -1 103360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_185_55
timestamp 1
transform 1 0 6164 0 -1 103360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_185_57
timestamp 1636968456
transform 1 0 6348 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_185_69
timestamp 1
transform 1 0 7452 0 -1 103360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_185_1122
timestamp 1636968456
transform 1 0 104328 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_1134
timestamp 1636968456
transform 1 0 105432 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_1146
timestamp 1636968456
transform 1 0 106536 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_185_1158
timestamp 1
transform 1 0 107640 0 -1 103360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_185_1166
timestamp 1
transform 1 0 108376 0 -1 103360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_186_3
timestamp 1636968456
transform 1 0 1380 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_15
timestamp 1636968456
transform 1 0 2484 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_186_27
timestamp 1
transform 1 0 3588 0 1 103360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_186_29
timestamp 1636968456
transform 1 0 3772 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_41
timestamp 1636968456
transform 1 0 4876 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_53
timestamp 1636968456
transform 1 0 5980 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_65
timestamp 1
transform 1 0 7084 0 1 103360
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_186_1122
timestamp 1636968456
transform 1 0 104328 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_1134
timestamp 1636968456
transform 1 0 105432 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_186_1146
timestamp 1
transform 1 0 106536 0 1 103360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_186_1148
timestamp 1636968456
transform 1 0 106720 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_1160
timestamp 1
transform 1 0 107824 0 1 103360
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_187_8
timestamp 1636968456
transform 1 0 1840 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_20
timestamp 1636968456
transform 1 0 2944 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_32
timestamp 1636968456
transform 1 0 4048 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_44
timestamp 1636968456
transform 1 0 5152 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_57
timestamp 1636968456
transform 1 0 6348 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_187_69
timestamp 1
transform 1 0 7452 0 -1 104448
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_187_1122
timestamp 1636968456
transform 1 0 104328 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_1134
timestamp 1636968456
transform 1 0 105432 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_1146
timestamp 1636968456
transform 1 0 106536 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_187_1158
timestamp 1
transform 1 0 107640 0 -1 104448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_187_1166
timestamp 1
transform 1 0 108376 0 -1 104448
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_188_3
timestamp 1636968456
transform 1 0 1380 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_15
timestamp 1636968456
transform 1 0 2484 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_188_27
timestamp 1
transform 1 0 3588 0 1 104448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_188_29
timestamp 1636968456
transform 1 0 3772 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_41
timestamp 1636968456
transform 1 0 4876 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_53
timestamp 1636968456
transform 1 0 5980 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_65
timestamp 1
transform 1 0 7084 0 1 104448
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_188_1122
timestamp 1636968456
transform 1 0 104328 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_1134
timestamp 1636968456
transform 1 0 105432 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_188_1146
timestamp 1
transform 1 0 106536 0 1 104448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_188_1148
timestamp 1636968456
transform 1 0 106720 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_188_1160
timestamp 1
transform 1 0 107824 0 1 104448
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_189_3
timestamp 1636968456
transform 1 0 1380 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_15
timestamp 1636968456
transform 1 0 2484 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_27
timestamp 1636968456
transform 1 0 3588 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_39
timestamp 1636968456
transform 1 0 4692 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_189_51
timestamp 1
transform 1 0 5796 0 -1 105536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_189_55
timestamp 1
transform 1 0 6164 0 -1 105536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_189_57
timestamp 1636968456
transform 1 0 6348 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_189_69
timestamp 1
transform 1 0 7452 0 -1 105536
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_189_1122
timestamp 1636968456
transform 1 0 104328 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_1134
timestamp 1636968456
transform 1 0 105432 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_1146
timestamp 1636968456
transform 1 0 106536 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_189_1158
timestamp 1
transform 1 0 107640 0 -1 105536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_189_1166
timestamp 1
transform 1 0 108376 0 -1 105536
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_190_8
timestamp 1636968456
transform 1 0 1840 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_190_20
timestamp 1
transform 1 0 2944 0 1 105536
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_190_29
timestamp 1636968456
transform 1 0 3772 0 1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_190_41
timestamp 1636968456
transform 1 0 4876 0 1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_190_53
timestamp 1636968456
transform 1 0 5980 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_65
timestamp 1
transform 1 0 7084 0 1 105536
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_190_1122
timestamp 1636968456
transform 1 0 104328 0 1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_190_1134
timestamp 1636968456
transform 1 0 105432 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_190_1146
timestamp 1
transform 1 0 106536 0 1 105536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_190_1148
timestamp 1636968456
transform 1 0 106720 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_190_1160
timestamp 1
transform 1 0 107824 0 1 105536
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_191_3
timestamp 1636968456
transform 1 0 1380 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_15
timestamp 1636968456
transform 1 0 2484 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_27
timestamp 1636968456
transform 1 0 3588 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_39
timestamp 1636968456
transform 1 0 4692 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_191_51
timestamp 1
transform 1 0 5796 0 -1 106624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_191_55
timestamp 1
transform 1 0 6164 0 -1 106624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_191_57
timestamp 1636968456
transform 1 0 6348 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_191_69
timestamp 1
transform 1 0 7452 0 -1 106624
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_191_1122
timestamp 1636968456
transform 1 0 104328 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_1134
timestamp 1636968456
transform 1 0 105432 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_1146
timestamp 1636968456
transform 1 0 106536 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_191_1158
timestamp 1
transform 1 0 107640 0 -1 106624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_191_1166
timestamp 1
transform 1 0 108376 0 -1 106624
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_192_8
timestamp 1636968456
transform 1 0 1840 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_20
timestamp 1
transform 1 0 2944 0 1 106624
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_192_29
timestamp 1636968456
transform 1 0 3772 0 1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_192_41
timestamp 1636968456
transform 1 0 4876 0 1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_192_53
timestamp 1636968456
transform 1 0 5980 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_65
timestamp 1
transform 1 0 7084 0 1 106624
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_192_1122
timestamp 1636968456
transform 1 0 104328 0 1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_192_1134
timestamp 1636968456
transform 1 0 105432 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_192_1146
timestamp 1
transform 1 0 106536 0 1 106624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_192_1148
timestamp 1636968456
transform 1 0 106720 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_1160
timestamp 1
transform 1 0 107824 0 1 106624
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_193_3
timestamp 1636968456
transform 1 0 1380 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_15
timestamp 1636968456
transform 1 0 2484 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_27
timestamp 1636968456
transform 1 0 3588 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_39
timestamp 1636968456
transform 1 0 4692 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_193_51
timestamp 1
transform 1 0 5796 0 -1 107712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_193_55
timestamp 1
transform 1 0 6164 0 -1 107712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_193_57
timestamp 1636968456
transform 1 0 6348 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_193_69
timestamp 1
transform 1 0 7452 0 -1 107712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_193_1122
timestamp 1636968456
transform 1 0 104328 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_1134
timestamp 1636968456
transform 1 0 105432 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_1146
timestamp 1636968456
transform 1 0 106536 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_193_1158
timestamp 1
transform 1 0 107640 0 -1 107712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_193_1166
timestamp 1
transform 1 0 108376 0 -1 107712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_194_3
timestamp 1636968456
transform 1 0 1380 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_15
timestamp 1636968456
transform 1 0 2484 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_194_27
timestamp 1
transform 1 0 3588 0 1 107712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_194_29
timestamp 1636968456
transform 1 0 3772 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_41
timestamp 1636968456
transform 1 0 4876 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_53
timestamp 1636968456
transform 1 0 5980 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_65
timestamp 1
transform 1 0 7084 0 1 107712
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_194_1122
timestamp 1636968456
transform 1 0 104328 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_1134
timestamp 1636968456
transform 1 0 105432 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_194_1146
timestamp 1
transform 1 0 106536 0 1 107712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_194_1148
timestamp 1636968456
transform 1 0 106720 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_194_1160
timestamp 1
transform 1 0 107824 0 1 107712
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_195_8
timestamp 1636968456
transform 1 0 1840 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_20
timestamp 1636968456
transform 1 0 2944 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_32
timestamp 1636968456
transform 1 0 4048 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_44
timestamp 1636968456
transform 1 0 5152 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_57
timestamp 1636968456
transform 1 0 6348 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_195_69
timestamp 1
transform 1 0 7452 0 -1 108800
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_195_1122
timestamp 1636968456
transform 1 0 104328 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_1134
timestamp 1636968456
transform 1 0 105432 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_1146
timestamp 1636968456
transform 1 0 106536 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_195_1158
timestamp 1
transform 1 0 107640 0 -1 108800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_195_1166
timestamp 1
transform 1 0 108376 0 -1 108800
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_196_3
timestamp 1636968456
transform 1 0 1380 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_15
timestamp 1636968456
transform 1 0 2484 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_196_27
timestamp 1
transform 1 0 3588 0 1 108800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_196_29
timestamp 1636968456
transform 1 0 3772 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_41
timestamp 1636968456
transform 1 0 4876 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_53
timestamp 1636968456
transform 1 0 5980 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_65
timestamp 1
transform 1 0 7084 0 1 108800
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_196_1122
timestamp 1636968456
transform 1 0 104328 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_1134
timestamp 1636968456
transform 1 0 105432 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_196_1146
timestamp 1
transform 1 0 106536 0 1 108800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_196_1148
timestamp 1636968456
transform 1 0 106720 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_196_1160
timestamp 1
transform 1 0 107824 0 1 108800
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_197_8
timestamp 1636968456
transform 1 0 1840 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_20
timestamp 1636968456
transform 1 0 2944 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_32
timestamp 1636968456
transform 1 0 4048 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_44
timestamp 1636968456
transform 1 0 5152 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_57
timestamp 1636968456
transform 1 0 6348 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_197_69
timestamp 1
transform 1 0 7452 0 -1 109888
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_197_1122
timestamp 1636968456
transform 1 0 104328 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_1134
timestamp 1636968456
transform 1 0 105432 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_1146
timestamp 1636968456
transform 1 0 106536 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_197_1158
timestamp 1
transform 1 0 107640 0 -1 109888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_197_1166
timestamp 1
transform 1 0 108376 0 -1 109888
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_198_3
timestamp 1636968456
transform 1 0 1380 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_15
timestamp 1636968456
transform 1 0 2484 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_198_27
timestamp 1
transform 1 0 3588 0 1 109888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_198_29
timestamp 1636968456
transform 1 0 3772 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_41
timestamp 1636968456
transform 1 0 4876 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_53
timestamp 1636968456
transform 1 0 5980 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_65
timestamp 1
transform 1 0 7084 0 1 109888
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_198_1122
timestamp 1636968456
transform 1 0 104328 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_1134
timestamp 1636968456
transform 1 0 105432 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_198_1146
timestamp 1
transform 1 0 106536 0 1 109888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_198_1148
timestamp 1636968456
transform 1 0 106720 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_198_1160
timestamp 1
transform 1 0 107824 0 1 109888
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_199_3
timestamp 1636968456
transform 1 0 1380 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_15
timestamp 1636968456
transform 1 0 2484 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_27
timestamp 1636968456
transform 1 0 3588 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_39
timestamp 1636968456
transform 1 0 4692 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_199_51
timestamp 1
transform 1 0 5796 0 -1 110976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_199_55
timestamp 1
transform 1 0 6164 0 -1 110976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_199_57
timestamp 1636968456
transform 1 0 6348 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_199_69
timestamp 1
transform 1 0 7452 0 -1 110976
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_199_1122
timestamp 1636968456
transform 1 0 104328 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_1134
timestamp 1636968456
transform 1 0 105432 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_1146
timestamp 1636968456
transform 1 0 106536 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_1158
timestamp 1
transform 1 0 107640 0 -1 110976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_199_1166
timestamp 1
transform 1 0 108376 0 -1 110976
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_200_8
timestamp 1636968456
transform 1 0 1840 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_200_20
timestamp 1
transform 1 0 2944 0 1 110976
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_200_29
timestamp 1636968456
transform 1 0 3772 0 1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_200_41
timestamp 1636968456
transform 1 0 4876 0 1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_200_53
timestamp 1636968456
transform 1 0 5980 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_65
timestamp 1
transform 1 0 7084 0 1 110976
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_200_1122
timestamp 1636968456
transform 1 0 104328 0 1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_200_1134
timestamp 1636968456
transform 1 0 105432 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_200_1146
timestamp 1
transform 1 0 106536 0 1 110976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_200_1148
timestamp 1636968456
transform 1 0 106720 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_200_1160
timestamp 1
transform 1 0 107824 0 1 110976
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_201_3
timestamp 1636968456
transform 1 0 1380 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_15
timestamp 1636968456
transform 1 0 2484 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_27
timestamp 1636968456
transform 1 0 3588 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_39
timestamp 1636968456
transform 1 0 4692 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_201_51
timestamp 1
transform 1 0 5796 0 -1 112064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_201_55
timestamp 1
transform 1 0 6164 0 -1 112064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_201_57
timestamp 1636968456
transform 1 0 6348 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_201_69
timestamp 1
transform 1 0 7452 0 -1 112064
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_201_1122
timestamp 1636968456
transform 1 0 104328 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_1134
timestamp 1636968456
transform 1 0 105432 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_1146
timestamp 1636968456
transform 1 0 106536 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_201_1158
timestamp 1
transform 1 0 107640 0 -1 112064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_201_1166
timestamp 1
transform 1 0 108376 0 -1 112064
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_202_3
timestamp 1636968456
transform 1 0 1380 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_15
timestamp 1636968456
transform 1 0 2484 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_202_27
timestamp 1
transform 1 0 3588 0 1 112064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_202_29
timestamp 1636968456
transform 1 0 3772 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_41
timestamp 1636968456
transform 1 0 4876 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_53
timestamp 1636968456
transform 1 0 5980 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_65
timestamp 1
transform 1 0 7084 0 1 112064
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_202_1122
timestamp 1636968456
transform 1 0 104328 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_1134
timestamp 1636968456
transform 1 0 105432 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_202_1146
timestamp 1
transform 1 0 106536 0 1 112064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_202_1148
timestamp 1636968456
transform 1 0 106720 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_202_1160
timestamp 1
transform 1 0 107824 0 1 112064
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_203_3
timestamp 1636968456
transform 1 0 1380 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_15
timestamp 1636968456
transform 1 0 2484 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_27
timestamp 1636968456
transform 1 0 3588 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_39
timestamp 1636968456
transform 1 0 4692 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_203_51
timestamp 1
transform 1 0 5796 0 -1 113152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_203_55
timestamp 1
transform 1 0 6164 0 -1 113152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_203_57
timestamp 1636968456
transform 1 0 6348 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_203_69
timestamp 1
transform 1 0 7452 0 -1 113152
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_203_1122
timestamp 1636968456
transform 1 0 104328 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_1134
timestamp 1636968456
transform 1 0 105432 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_1146
timestamp 1636968456
transform 1 0 106536 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_203_1158
timestamp 1
transform 1 0 107640 0 -1 113152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_203_1166
timestamp 1
transform 1 0 108376 0 -1 113152
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_204_3
timestamp 1636968456
transform 1 0 1380 0 1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_204_15
timestamp 1636968456
transform 1 0 2484 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_204_27
timestamp 1
transform 1 0 3588 0 1 113152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_204_29
timestamp 1636968456
transform 1 0 3772 0 1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_204_41
timestamp 1636968456
transform 1 0 4876 0 1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_204_53
timestamp 1636968456
transform 1 0 5980 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_65
timestamp 1
transform 1 0 7084 0 1 113152
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_204_1122
timestamp 1636968456
transform 1 0 104328 0 1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_204_1134
timestamp 1636968456
transform 1 0 105432 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_204_1146
timestamp 1
transform 1 0 106536 0 1 113152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_204_1148
timestamp 1636968456
transform 1 0 106720 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_204_1160
timestamp 1
transform 1 0 107824 0 1 113152
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_205_3
timestamp 1636968456
transform 1 0 1380 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_15
timestamp 1636968456
transform 1 0 2484 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_27
timestamp 1636968456
transform 1 0 3588 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_39
timestamp 1636968456
transform 1 0 4692 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_205_51
timestamp 1
transform 1 0 5796 0 -1 114240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_205_55
timestamp 1
transform 1 0 6164 0 -1 114240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_205_57
timestamp 1636968456
transform 1 0 6348 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_205_69
timestamp 1
transform 1 0 7452 0 -1 114240
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_205_1122
timestamp 1636968456
transform 1 0 104328 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_1134
timestamp 1636968456
transform 1 0 105432 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_1146
timestamp 1636968456
transform 1 0 106536 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_205_1158
timestamp 1
transform 1 0 107640 0 -1 114240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_205_1166
timestamp 1
transform 1 0 108376 0 -1 114240
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_206_3
timestamp 1636968456
transform 1 0 1380 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_15
timestamp 1636968456
transform 1 0 2484 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_206_27
timestamp 1
transform 1 0 3588 0 1 114240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_206_29
timestamp 1636968456
transform 1 0 3772 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_41
timestamp 1636968456
transform 1 0 4876 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_53
timestamp 1636968456
transform 1 0 5980 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_65
timestamp 1
transform 1 0 7084 0 1 114240
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_206_1122
timestamp 1636968456
transform 1 0 104328 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_1134
timestamp 1636968456
transform 1 0 105432 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_206_1146
timestamp 1
transform 1 0 106536 0 1 114240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_206_1148
timestamp 1636968456
transform 1 0 106720 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_206_1160
timestamp 1
transform 1 0 107824 0 1 114240
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_207_3
timestamp 1636968456
transform 1 0 1380 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_15
timestamp 1636968456
transform 1 0 2484 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_27
timestamp 1636968456
transform 1 0 3588 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_39
timestamp 1636968456
transform 1 0 4692 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_207_51
timestamp 1
transform 1 0 5796 0 -1 115328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_55
timestamp 1
transform 1 0 6164 0 -1 115328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_207_57
timestamp 1636968456
transform 1 0 6348 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_207_69
timestamp 1
transform 1 0 7452 0 -1 115328
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_207_1122
timestamp 1636968456
transform 1 0 104328 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_1134
timestamp 1636968456
transform 1 0 105432 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_1146
timestamp 1636968456
transform 1 0 106536 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_207_1158
timestamp 1
transform 1 0 107640 0 -1 115328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_207_1166
timestamp 1
transform 1 0 108376 0 -1 115328
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_208_3
timestamp 1636968456
transform 1 0 1380 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_15
timestamp 1636968456
transform 1 0 2484 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_208_27
timestamp 1
transform 1 0 3588 0 1 115328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_208_29
timestamp 1636968456
transform 1 0 3772 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_41
timestamp 1636968456
transform 1 0 4876 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_53
timestamp 1636968456
transform 1 0 5980 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_65
timestamp 1
transform 1 0 7084 0 1 115328
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_208_1122
timestamp 1636968456
transform 1 0 104328 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_1134
timestamp 1636968456
transform 1 0 105432 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_208_1146
timestamp 1
transform 1 0 106536 0 1 115328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_208_1148
timestamp 1636968456
transform 1 0 106720 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_208_1160
timestamp 1
transform 1 0 107824 0 1 115328
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_209_3
timestamp 1636968456
transform 1 0 1380 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_15
timestamp 1636968456
transform 1 0 2484 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_27
timestamp 1636968456
transform 1 0 3588 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_39
timestamp 1636968456
transform 1 0 4692 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_209_51
timestamp 1
transform 1 0 5796 0 -1 116416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_55
timestamp 1
transform 1 0 6164 0 -1 116416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_209_57
timestamp 1636968456
transform 1 0 6348 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_209_69
timestamp 1
transform 1 0 7452 0 -1 116416
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_209_1122
timestamp 1636968456
transform 1 0 104328 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_1134
timestamp 1636968456
transform 1 0 105432 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_1146
timestamp 1636968456
transform 1 0 106536 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_209_1158
timestamp 1
transform 1 0 107640 0 -1 116416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_209_1166
timestamp 1
transform 1 0 108376 0 -1 116416
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_210_3
timestamp 1636968456
transform 1 0 1380 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_15
timestamp 1636968456
transform 1 0 2484 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_210_27
timestamp 1
transform 1 0 3588 0 1 116416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_210_29
timestamp 1636968456
transform 1 0 3772 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_41
timestamp 1636968456
transform 1 0 4876 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_53
timestamp 1636968456
transform 1 0 5980 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_65
timestamp 1
transform 1 0 7084 0 1 116416
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_210_1122
timestamp 1636968456
transform 1 0 104328 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_1134
timestamp 1636968456
transform 1 0 105432 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_210_1146
timestamp 1
transform 1 0 106536 0 1 116416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_210_1148
timestamp 1636968456
transform 1 0 106720 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_210_1160
timestamp 1
transform 1 0 107824 0 1 116416
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_211_3
timestamp 1636968456
transform 1 0 1380 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_15
timestamp 1636968456
transform 1 0 2484 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_27
timestamp 1636968456
transform 1 0 3588 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_39
timestamp 1636968456
transform 1 0 4692 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_211_51
timestamp 1
transform 1 0 5796 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_211_55
timestamp 1
transform 1 0 6164 0 -1 117504
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_211_57
timestamp 1636968456
transform 1 0 6348 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_211_69
timestamp 1
transform 1 0 7452 0 -1 117504
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_211_1122
timestamp 1636968456
transform 1 0 104328 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_1134
timestamp 1636968456
transform 1 0 105432 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_1146
timestamp 1636968456
transform 1 0 106536 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_211_1158
timestamp 1
transform 1 0 107640 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_211_1166
timestamp 1
transform 1 0 108376 0 -1 117504
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_212_3
timestamp 1636968456
transform 1 0 1380 0 1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_212_15
timestamp 1636968456
transform 1 0 2484 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_212_27
timestamp 1
transform 1 0 3588 0 1 117504
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_212_29
timestamp 1636968456
transform 1 0 3772 0 1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_212_41
timestamp 1636968456
transform 1 0 4876 0 1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_212_53
timestamp 1636968456
transform 1 0 5980 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_212_65
timestamp 1
transform 1 0 7084 0 1 117504
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_212_1122
timestamp 1636968456
transform 1 0 104328 0 1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_212_1134
timestamp 1636968456
transform 1 0 105432 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_212_1146
timestamp 1
transform 1 0 106536 0 1 117504
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_212_1148
timestamp 1636968456
transform 1 0 106720 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_212_1160
timestamp 1
transform 1 0 107824 0 1 117504
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_213_3
timestamp 1636968456
transform 1 0 1380 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_15
timestamp 1636968456
transform 1 0 2484 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_27
timestamp 1636968456
transform 1 0 3588 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_39
timestamp 1636968456
transform 1 0 4692 0 -1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_213_51
timestamp 1
transform 1 0 5796 0 -1 118592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_213_55
timestamp 1
transform 1 0 6164 0 -1 118592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_213_57
timestamp 1636968456
transform 1 0 6348 0 -1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_213_69
timestamp 1
transform 1 0 7452 0 -1 118592
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_213_1122
timestamp 1636968456
transform 1 0 104328 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_1134
timestamp 1636968456
transform 1 0 105432 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_1146
timestamp 1636968456
transform 1 0 106536 0 -1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_213_1158
timestamp 1
transform 1 0 107640 0 -1 118592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_213_1166
timestamp 1
transform 1 0 108376 0 -1 118592
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_214_3
timestamp 1636968456
transform 1 0 1380 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_15
timestamp 1636968456
transform 1 0 2484 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_214_27
timestamp 1
transform 1 0 3588 0 1 118592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_214_29
timestamp 1636968456
transform 1 0 3772 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_41
timestamp 1636968456
transform 1 0 4876 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_53
timestamp 1636968456
transform 1 0 5980 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_214_65
timestamp 1
transform 1 0 7084 0 1 118592
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_214_1122
timestamp 1636968456
transform 1 0 104328 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_1134
timestamp 1636968456
transform 1 0 105432 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_214_1146
timestamp 1
transform 1 0 106536 0 1 118592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_214_1148
timestamp 1636968456
transform 1 0 106720 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_214_1160
timestamp 1
transform 1 0 107824 0 1 118592
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_215_3
timestamp 1636968456
transform 1 0 1380 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_15
timestamp 1636968456
transform 1 0 2484 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_27
timestamp 1636968456
transform 1 0 3588 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_39
timestamp 1636968456
transform 1 0 4692 0 -1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_215_51
timestamp 1
transform 1 0 5796 0 -1 119680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_215_55
timestamp 1
transform 1 0 6164 0 -1 119680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_215_57
timestamp 1636968456
transform 1 0 6348 0 -1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_215_69
timestamp 1
transform 1 0 7452 0 -1 119680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_215_1122
timestamp 1636968456
transform 1 0 104328 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_1134
timestamp 1636968456
transform 1 0 105432 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_1146
timestamp 1636968456
transform 1 0 106536 0 -1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_215_1158
timestamp 1
transform 1 0 107640 0 -1 119680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_215_1166
timestamp 1
transform 1 0 108376 0 -1 119680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_216_3
timestamp 1636968456
transform 1 0 1380 0 1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_216_15
timestamp 1636968456
transform 1 0 2484 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_216_27
timestamp 1
transform 1 0 3588 0 1 119680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_216_29
timestamp 1636968456
transform 1 0 3772 0 1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_216_41
timestamp 1636968456
transform 1 0 4876 0 1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_216_53
timestamp 1636968456
transform 1 0 5980 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_216_65
timestamp 1
transform 1 0 7084 0 1 119680
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_216_1122
timestamp 1636968456
transform 1 0 104328 0 1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_216_1134
timestamp 1636968456
transform 1 0 105432 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_216_1146
timestamp 1
transform 1 0 106536 0 1 119680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_216_1148
timestamp 1636968456
transform 1 0 106720 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_216_1160
timestamp 1
transform 1 0 107824 0 1 119680
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_217_3
timestamp 1636968456
transform 1 0 1380 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_15
timestamp 1636968456
transform 1 0 2484 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_27
timestamp 1636968456
transform 1 0 3588 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_39
timestamp 1636968456
transform 1 0 4692 0 -1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_217_51
timestamp 1
transform 1 0 5796 0 -1 120768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_217_55
timestamp 1
transform 1 0 6164 0 -1 120768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_217_57
timestamp 1636968456
transform 1 0 6348 0 -1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_217_69
timestamp 1
transform 1 0 7452 0 -1 120768
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_217_1122
timestamp 1636968456
transform 1 0 104328 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_1134
timestamp 1636968456
transform 1 0 105432 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_1146
timestamp 1636968456
transform 1 0 106536 0 -1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_217_1158
timestamp 1
transform 1 0 107640 0 -1 120768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_217_1166
timestamp 1
transform 1 0 108376 0 -1 120768
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_218_3
timestamp 1636968456
transform 1 0 1380 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_15
timestamp 1636968456
transform 1 0 2484 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_218_27
timestamp 1
transform 1 0 3588 0 1 120768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_218_29
timestamp 1636968456
transform 1 0 3772 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_41
timestamp 1636968456
transform 1 0 4876 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_53
timestamp 1636968456
transform 1 0 5980 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_218_65
timestamp 1
transform 1 0 7084 0 1 120768
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_218_1122
timestamp 1636968456
transform 1 0 104328 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_1134
timestamp 1636968456
transform 1 0 105432 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_218_1146
timestamp 1
transform 1 0 106536 0 1 120768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_218_1148
timestamp 1636968456
transform 1 0 106720 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_218_1160
timestamp 1
transform 1 0 107824 0 1 120768
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_219_3
timestamp 1636968456
transform 1 0 1380 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_15
timestamp 1636968456
transform 1 0 2484 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_27
timestamp 1636968456
transform 1 0 3588 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_39
timestamp 1636968456
transform 1 0 4692 0 -1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_219_51
timestamp 1
transform 1 0 5796 0 -1 121856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_219_55
timestamp 1
transform 1 0 6164 0 -1 121856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_219_57
timestamp 1636968456
transform 1 0 6348 0 -1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_219_69
timestamp 1
transform 1 0 7452 0 -1 121856
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_219_1122
timestamp 1636968456
transform 1 0 104328 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_1134
timestamp 1636968456
transform 1 0 105432 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_1146
timestamp 1636968456
transform 1 0 106536 0 -1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_219_1158
timestamp 1
transform 1 0 107640 0 -1 121856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_219_1166
timestamp 1
transform 1 0 108376 0 -1 121856
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_220_3
timestamp 1636968456
transform 1 0 1380 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_15
timestamp 1636968456
transform 1 0 2484 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_220_27
timestamp 1
transform 1 0 3588 0 1 121856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_220_29
timestamp 1636968456
transform 1 0 3772 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_41
timestamp 1636968456
transform 1 0 4876 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_53
timestamp 1636968456
transform 1 0 5980 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_220_65
timestamp 1
transform 1 0 7084 0 1 121856
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_220_1122
timestamp 1636968456
transform 1 0 104328 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_1134
timestamp 1636968456
transform 1 0 105432 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_220_1146
timestamp 1
transform 1 0 106536 0 1 121856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_220_1148
timestamp 1636968456
transform 1 0 106720 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_220_1160
timestamp 1
transform 1 0 107824 0 1 121856
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_221_3
timestamp 1636968456
transform 1 0 1380 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_15
timestamp 1636968456
transform 1 0 2484 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_27
timestamp 1636968456
transform 1 0 3588 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_39
timestamp 1636968456
transform 1 0 4692 0 -1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_221_51
timestamp 1
transform 1 0 5796 0 -1 122944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_221_55
timestamp 1
transform 1 0 6164 0 -1 122944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_221_57
timestamp 1636968456
transform 1 0 6348 0 -1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_221_69
timestamp 1
transform 1 0 7452 0 -1 122944
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_221_1122
timestamp 1636968456
transform 1 0 104328 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_1134
timestamp 1636968456
transform 1 0 105432 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_1146
timestamp 1636968456
transform 1 0 106536 0 -1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_221_1158
timestamp 1
transform 1 0 107640 0 -1 122944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_221_1166
timestamp 1
transform 1 0 108376 0 -1 122944
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_222_3
timestamp 1636968456
transform 1 0 1380 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_15
timestamp 1636968456
transform 1 0 2484 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_222_27
timestamp 1
transform 1 0 3588 0 1 122944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_222_29
timestamp 1636968456
transform 1 0 3772 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_41
timestamp 1636968456
transform 1 0 4876 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_53
timestamp 1636968456
transform 1 0 5980 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_222_65
timestamp 1
transform 1 0 7084 0 1 122944
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_222_1122
timestamp 1636968456
transform 1 0 104328 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_1134
timestamp 1636968456
transform 1 0 105432 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_222_1146
timestamp 1
transform 1 0 106536 0 1 122944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_222_1148
timestamp 1636968456
transform 1 0 106720 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_222_1160
timestamp 1
transform 1 0 107824 0 1 122944
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_223_3
timestamp 1636968456
transform 1 0 1380 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_15
timestamp 1636968456
transform 1 0 2484 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_27
timestamp 1636968456
transform 1 0 3588 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_39
timestamp 1636968456
transform 1 0 4692 0 -1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_223_51
timestamp 1
transform 1 0 5796 0 -1 124032
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_223_55
timestamp 1
transform 1 0 6164 0 -1 124032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_223_57
timestamp 1636968456
transform 1 0 6348 0 -1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_223_69
timestamp 1
transform 1 0 7452 0 -1 124032
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_223_1122
timestamp 1636968456
transform 1 0 104328 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_1134
timestamp 1636968456
transform 1 0 105432 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_1146
timestamp 1636968456
transform 1 0 106536 0 -1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_223_1158
timestamp 1
transform 1 0 107640 0 -1 124032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_223_1166
timestamp 1
transform 1 0 108376 0 -1 124032
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_224_3
timestamp 1636968456
transform 1 0 1380 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_15
timestamp 1636968456
transform 1 0 2484 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_224_27
timestamp 1
transform 1 0 3588 0 1 124032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_224_29
timestamp 1636968456
transform 1 0 3772 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_41
timestamp 1636968456
transform 1 0 4876 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_53
timestamp 1636968456
transform 1 0 5980 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_224_65
timestamp 1
transform 1 0 7084 0 1 124032
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_224_1122
timestamp 1636968456
transform 1 0 104328 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_1134
timestamp 1636968456
transform 1 0 105432 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_224_1146
timestamp 1
transform 1 0 106536 0 1 124032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_224_1148
timestamp 1636968456
transform 1 0 106720 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_224_1160
timestamp 1
transform 1 0 107824 0 1 124032
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_225_3
timestamp 1636968456
transform 1 0 1380 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_15
timestamp 1636968456
transform 1 0 2484 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_27
timestamp 1636968456
transform 1 0 3588 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_39
timestamp 1636968456
transform 1 0 4692 0 -1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_225_51
timestamp 1
transform 1 0 5796 0 -1 125120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_225_55
timestamp 1
transform 1 0 6164 0 -1 125120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_225_57
timestamp 1636968456
transform 1 0 6348 0 -1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_225_69
timestamp 1
transform 1 0 7452 0 -1 125120
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_225_1122
timestamp 1636968456
transform 1 0 104328 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_1134
timestamp 1636968456
transform 1 0 105432 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_1146
timestamp 1636968456
transform 1 0 106536 0 -1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_225_1158
timestamp 1
transform 1 0 107640 0 -1 125120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_225_1166
timestamp 1
transform 1 0 108376 0 -1 125120
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_226_3
timestamp 1636968456
transform 1 0 1380 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_15
timestamp 1636968456
transform 1 0 2484 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_226_27
timestamp 1
transform 1 0 3588 0 1 125120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_226_29
timestamp 1636968456
transform 1 0 3772 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_41
timestamp 1636968456
transform 1 0 4876 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_53
timestamp 1636968456
transform 1 0 5980 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_226_65
timestamp 1
transform 1 0 7084 0 1 125120
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_226_1122
timestamp 1636968456
transform 1 0 104328 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_1134
timestamp 1636968456
transform 1 0 105432 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_226_1146
timestamp 1
transform 1 0 106536 0 1 125120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_226_1148
timestamp 1636968456
transform 1 0 106720 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_226_1160
timestamp 1
transform 1 0 107824 0 1 125120
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_227_3
timestamp 1636968456
transform 1 0 1380 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_15
timestamp 1636968456
transform 1 0 2484 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_27
timestamp 1636968456
transform 1 0 3588 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_39
timestamp 1636968456
transform 1 0 4692 0 -1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_227_51
timestamp 1
transform 1 0 5796 0 -1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_227_55
timestamp 1
transform 1 0 6164 0 -1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_227_57
timestamp 1636968456
transform 1 0 6348 0 -1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_227_69
timestamp 1
transform 1 0 7452 0 -1 126208
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_227_1122
timestamp 1636968456
transform 1 0 104328 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_1134
timestamp 1636968456
transform 1 0 105432 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_1146
timestamp 1636968456
transform 1 0 106536 0 -1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_227_1158
timestamp 1
transform 1 0 107640 0 -1 126208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_227_1166
timestamp 1
transform 1 0 108376 0 -1 126208
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_228_3
timestamp 1636968456
transform 1 0 1380 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_15
timestamp 1636968456
transform 1 0 2484 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_228_27
timestamp 1
transform 1 0 3588 0 1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_228_29
timestamp 1636968456
transform 1 0 3772 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_41
timestamp 1636968456
transform 1 0 4876 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_53
timestamp 1636968456
transform 1 0 5980 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_228_65
timestamp 1
transform 1 0 7084 0 1 126208
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1122
timestamp 1636968456
transform 1 0 104328 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1134
timestamp 1636968456
transform 1 0 105432 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_228_1146
timestamp 1
transform 1 0 106536 0 1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1148
timestamp 1636968456
transform 1 0 106720 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_228_1160
timestamp 1
transform 1 0 107824 0 1 126208
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_229_3
timestamp 1636968456
transform 1 0 1380 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_15
timestamp 1636968456
transform 1 0 2484 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_27
timestamp 1636968456
transform 1 0 3588 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_39
timestamp 1636968456
transform 1 0 4692 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_229_51
timestamp 1
transform 1 0 5796 0 -1 127296
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_229_55
timestamp 1
transform 1 0 6164 0 -1 127296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_229_57
timestamp 1636968456
transform 1 0 6348 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_229_69
timestamp 1
transform 1 0 7452 0 -1 127296
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1122
timestamp 1636968456
transform 1 0 104328 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1134
timestamp 1636968456
transform 1 0 105432 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1146
timestamp 1636968456
transform 1 0 106536 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_229_1158
timestamp 1
transform 1 0 107640 0 -1 127296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_229_1166
timestamp 1
transform 1 0 108376 0 -1 127296
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_230_3
timestamp 1636968456
transform 1 0 1380 0 1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_230_15
timestamp 1636968456
transform 1 0 2484 0 1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_230_27
timestamp 1
transform 1 0 3588 0 1 127296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_230_29
timestamp 1636968456
transform 1 0 3772 0 1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_230_41
timestamp 1636968456
transform 1 0 4876 0 1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_230_53
timestamp 1636968456
transform 1 0 5980 0 1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_230_65
timestamp 1
transform 1 0 7084 0 1 127296
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_230_1122
timestamp 1636968456
transform 1 0 104328 0 1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_230_1134
timestamp 1636968456
transform 1 0 105432 0 1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_230_1146
timestamp 1
transform 1 0 106536 0 1 127296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_230_1148
timestamp 1636968456
transform 1 0 106720 0 1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_230_1160
timestamp 1
transform 1 0 107824 0 1 127296
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_231_3
timestamp 1636968456
transform 1 0 1380 0 -1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_231_15
timestamp 1636968456
transform 1 0 2484 0 -1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_231_27
timestamp 1636968456
transform 1 0 3588 0 -1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_231_39
timestamp 1636968456
transform 1 0 4692 0 -1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_231_51
timestamp 1
transform 1 0 5796 0 -1 128384
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_231_55
timestamp 1
transform 1 0 6164 0 -1 128384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_231_57
timestamp 1636968456
transform 1 0 6348 0 -1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_231_69
timestamp 1
transform 1 0 7452 0 -1 128384
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_231_1122
timestamp 1636968456
transform 1 0 104328 0 -1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_231_1134
timestamp 1636968456
transform 1 0 105432 0 -1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_231_1146
timestamp 1636968456
transform 1 0 106536 0 -1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_231_1158
timestamp 1
transform 1 0 107640 0 -1 128384
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_231_1166
timestamp 1
transform 1 0 108376 0 -1 128384
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_232_3
timestamp 1636968456
transform 1 0 1380 0 1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_232_15
timestamp 1636968456
transform 1 0 2484 0 1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_232_27
timestamp 1
transform 1 0 3588 0 1 128384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_232_29
timestamp 1636968456
transform 1 0 3772 0 1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_232_41
timestamp 1636968456
transform 1 0 4876 0 1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_232_53
timestamp 1636968456
transform 1 0 5980 0 1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_232_65
timestamp 1
transform 1 0 7084 0 1 128384
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_232_1122
timestamp 1636968456
transform 1 0 104328 0 1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_232_1134
timestamp 1636968456
transform 1 0 105432 0 1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_232_1146
timestamp 1
transform 1 0 106536 0 1 128384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_232_1148
timestamp 1636968456
transform 1 0 106720 0 1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_232_1160
timestamp 1
transform 1 0 107824 0 1 128384
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_233_3
timestamp 1636968456
transform 1 0 1380 0 -1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_233_15
timestamp 1636968456
transform 1 0 2484 0 -1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_233_27
timestamp 1636968456
transform 1 0 3588 0 -1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_233_39
timestamp 1636968456
transform 1 0 4692 0 -1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_233_51
timestamp 1
transform 1 0 5796 0 -1 129472
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_233_55
timestamp 1
transform 1 0 6164 0 -1 129472
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_233_57
timestamp 1636968456
transform 1 0 6348 0 -1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_233_69
timestamp 1
transform 1 0 7452 0 -1 129472
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_233_1122
timestamp 1636968456
transform 1 0 104328 0 -1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_233_1134
timestamp 1636968456
transform 1 0 105432 0 -1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_233_1146
timestamp 1636968456
transform 1 0 106536 0 -1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_233_1158
timestamp 1
transform 1 0 107640 0 -1 129472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_233_1166
timestamp 1
transform 1 0 108376 0 -1 129472
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_234_3
timestamp 1636968456
transform 1 0 1380 0 1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_234_15
timestamp 1636968456
transform 1 0 2484 0 1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_234_27
timestamp 1
transform 1 0 3588 0 1 129472
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_234_29
timestamp 1636968456
transform 1 0 3772 0 1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_234_41
timestamp 1636968456
transform 1 0 4876 0 1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_234_53
timestamp 1636968456
transform 1 0 5980 0 1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_234_65
timestamp 1
transform 1 0 7084 0 1 129472
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_234_1125
timestamp 1636968456
transform 1 0 104604 0 1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_234_1137
timestamp 1
transform 1 0 105708 0 1 129472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_234_1145
timestamp 1
transform 1 0 106444 0 1 129472
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_234_1148
timestamp 1636968456
transform 1 0 106720 0 1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_234_1160
timestamp 1
transform 1 0 107824 0 1 129472
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_235_3
timestamp 1636968456
transform 1 0 1380 0 -1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_235_15
timestamp 1636968456
transform 1 0 2484 0 -1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_235_27
timestamp 1636968456
transform 1 0 3588 0 -1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_235_39
timestamp 1636968456
transform 1 0 4692 0 -1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_235_51
timestamp 1
transform 1 0 5796 0 -1 130560
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_235_55
timestamp 1
transform 1 0 6164 0 -1 130560
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_235_57
timestamp 1636968456
transform 1 0 6348 0 -1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_235_69
timestamp 1
transform 1 0 7452 0 -1 130560
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_235_1122
timestamp 1636968456
transform 1 0 104328 0 -1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_235_1134
timestamp 1636968456
transform 1 0 105432 0 -1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_235_1146
timestamp 1636968456
transform 1 0 106536 0 -1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_235_1158
timestamp 1
transform 1 0 107640 0 -1 130560
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_235_1166
timestamp 1
transform 1 0 108376 0 -1 130560
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_236_3
timestamp 1636968456
transform 1 0 1380 0 1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_236_15
timestamp 1636968456
transform 1 0 2484 0 1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_236_27
timestamp 1
transform 1 0 3588 0 1 130560
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_236_29
timestamp 1636968456
transform 1 0 3772 0 1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_236_41
timestamp 1636968456
transform 1 0 4876 0 1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_236_53
timestamp 1636968456
transform 1 0 5980 0 1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_236_65
timestamp 1
transform 1 0 7084 0 1 130560
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_236_1122
timestamp 1636968456
transform 1 0 104328 0 1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_236_1134
timestamp 1636968456
transform 1 0 105432 0 1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_236_1146
timestamp 1
transform 1 0 106536 0 1 130560
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_236_1148
timestamp 1636968456
transform 1 0 106720 0 1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_236_1160
timestamp 1
transform 1 0 107824 0 1 130560
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_237_3
timestamp 1636968456
transform 1 0 1380 0 -1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_237_15
timestamp 1636968456
transform 1 0 2484 0 -1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_237_27
timestamp 1636968456
transform 1 0 3588 0 -1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_237_39
timestamp 1636968456
transform 1 0 4692 0 -1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_237_51
timestamp 1
transform 1 0 5796 0 -1 131648
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_237_55
timestamp 1
transform 1 0 6164 0 -1 131648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_237_57
timestamp 1636968456
transform 1 0 6348 0 -1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_237_69
timestamp 1
transform 1 0 7452 0 -1 131648
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_237_1122
timestamp 1636968456
transform 1 0 104328 0 -1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_237_1134
timestamp 1636968456
transform 1 0 105432 0 -1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_237_1146
timestamp 1636968456
transform 1 0 106536 0 -1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_237_1158
timestamp 1
transform 1 0 107640 0 -1 131648
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_237_1166
timestamp 1
transform 1 0 108376 0 -1 131648
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_238_3
timestamp 1636968456
transform 1 0 1380 0 1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_238_15
timestamp 1636968456
transform 1 0 2484 0 1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_238_27
timestamp 1
transform 1 0 3588 0 1 131648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_238_29
timestamp 1636968456
transform 1 0 3772 0 1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_238_41
timestamp 1636968456
transform 1 0 4876 0 1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_238_53
timestamp 1636968456
transform 1 0 5980 0 1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_238_65
timestamp 1
transform 1 0 7084 0 1 131648
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_238_1122
timestamp 1636968456
transform 1 0 104328 0 1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_238_1134
timestamp 1636968456
transform 1 0 105432 0 1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_238_1146
timestamp 1
transform 1 0 106536 0 1 131648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_238_1148
timestamp 1636968456
transform 1 0 106720 0 1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_238_1160
timestamp 1
transform 1 0 107824 0 1 131648
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_239_3
timestamp 1636968456
transform 1 0 1380 0 -1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_239_15
timestamp 1636968456
transform 1 0 2484 0 -1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_239_27
timestamp 1636968456
transform 1 0 3588 0 -1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_239_39
timestamp 1636968456
transform 1 0 4692 0 -1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_239_51
timestamp 1
transform 1 0 5796 0 -1 132736
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_239_55
timestamp 1
transform 1 0 6164 0 -1 132736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_239_57
timestamp 1636968456
transform 1 0 6348 0 -1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_239_69
timestamp 1
transform 1 0 7452 0 -1 132736
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_239_1122
timestamp 1636968456
transform 1 0 104328 0 -1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_239_1134
timestamp 1636968456
transform 1 0 105432 0 -1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_239_1146
timestamp 1636968456
transform 1 0 106536 0 -1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_239_1158
timestamp 1
transform 1 0 107640 0 -1 132736
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_239_1166
timestamp 1
transform 1 0 108376 0 -1 132736
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_240_3
timestamp 1636968456
transform 1 0 1380 0 1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_240_15
timestamp 1636968456
transform 1 0 2484 0 1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_240_27
timestamp 1
transform 1 0 3588 0 1 132736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_240_29
timestamp 1636968456
transform 1 0 3772 0 1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_240_41
timestamp 1636968456
transform 1 0 4876 0 1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_240_53
timestamp 1636968456
transform 1 0 5980 0 1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_240_65
timestamp 1
transform 1 0 7084 0 1 132736
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_240_1122
timestamp 1636968456
transform 1 0 104328 0 1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_240_1134
timestamp 1636968456
transform 1 0 105432 0 1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_240_1146
timestamp 1
transform 1 0 106536 0 1 132736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_240_1148
timestamp 1636968456
transform 1 0 106720 0 1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_240_1160
timestamp 1
transform 1 0 107824 0 1 132736
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_241_3
timestamp 1636968456
transform 1 0 1380 0 -1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_241_15
timestamp 1636968456
transform 1 0 2484 0 -1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_241_27
timestamp 1636968456
transform 1 0 3588 0 -1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_241_39
timestamp 1636968456
transform 1 0 4692 0 -1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_241_51
timestamp 1
transform 1 0 5796 0 -1 133824
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_241_55
timestamp 1
transform 1 0 6164 0 -1 133824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_241_57
timestamp 1636968456
transform 1 0 6348 0 -1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_241_69
timestamp 1
transform 1 0 7452 0 -1 133824
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_241_1122
timestamp 1636968456
transform 1 0 104328 0 -1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_241_1134
timestamp 1636968456
transform 1 0 105432 0 -1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_241_1146
timestamp 1636968456
transform 1 0 106536 0 -1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_241_1158
timestamp 1
transform 1 0 107640 0 -1 133824
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_241_1166
timestamp 1
transform 1 0 108376 0 -1 133824
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_242_3
timestamp 1636968456
transform 1 0 1380 0 1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_242_15
timestamp 1636968456
transform 1 0 2484 0 1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_242_27
timestamp 1
transform 1 0 3588 0 1 133824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_242_29
timestamp 1636968456
transform 1 0 3772 0 1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_242_41
timestamp 1636968456
transform 1 0 4876 0 1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_242_53
timestamp 1636968456
transform 1 0 5980 0 1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_242_65
timestamp 1
transform 1 0 7084 0 1 133824
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_242_1122
timestamp 1636968456
transform 1 0 104328 0 1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_242_1134
timestamp 1636968456
transform 1 0 105432 0 1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_242_1146
timestamp 1
transform 1 0 106536 0 1 133824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_242_1148
timestamp 1636968456
transform 1 0 106720 0 1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_242_1160
timestamp 1
transform 1 0 107824 0 1 133824
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_243_3
timestamp 1636968456
transform 1 0 1380 0 -1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_243_15
timestamp 1636968456
transform 1 0 2484 0 -1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_243_27
timestamp 1636968456
transform 1 0 3588 0 -1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_243_39
timestamp 1636968456
transform 1 0 4692 0 -1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_243_51
timestamp 1
transform 1 0 5796 0 -1 134912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_243_55
timestamp 1
transform 1 0 6164 0 -1 134912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_243_57
timestamp 1636968456
transform 1 0 6348 0 -1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_243_69
timestamp 1
transform 1 0 7452 0 -1 134912
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_243_1122
timestamp 1636968456
transform 1 0 104328 0 -1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_243_1134
timestamp 1636968456
transform 1 0 105432 0 -1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_243_1146
timestamp 1636968456
transform 1 0 106536 0 -1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_243_1158
timestamp 1
transform 1 0 107640 0 -1 134912
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_243_1166
timestamp 1
transform 1 0 108376 0 -1 134912
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_244_3
timestamp 1636968456
transform 1 0 1380 0 1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_244_15
timestamp 1636968456
transform 1 0 2484 0 1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_244_27
timestamp 1
transform 1 0 3588 0 1 134912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_244_29
timestamp 1636968456
transform 1 0 3772 0 1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_244_41
timestamp 1636968456
transform 1 0 4876 0 1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_244_53
timestamp 1636968456
transform 1 0 5980 0 1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_244_65
timestamp 1
transform 1 0 7084 0 1 134912
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_244_1122
timestamp 1636968456
transform 1 0 104328 0 1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_244_1134
timestamp 1636968456
transform 1 0 105432 0 1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_244_1146
timestamp 1
transform 1 0 106536 0 1 134912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_244_1148
timestamp 1636968456
transform 1 0 106720 0 1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_244_1160
timestamp 1
transform 1 0 107824 0 1 134912
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_245_3
timestamp 1636968456
transform 1 0 1380 0 -1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_245_15
timestamp 1636968456
transform 1 0 2484 0 -1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_245_27
timestamp 1636968456
transform 1 0 3588 0 -1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_245_39
timestamp 1636968456
transform 1 0 4692 0 -1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_245_51
timestamp 1
transform 1 0 5796 0 -1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_245_55
timestamp 1
transform 1 0 6164 0 -1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_245_57
timestamp 1636968456
transform 1 0 6348 0 -1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_245_69
timestamp 1
transform 1 0 7452 0 -1 136000
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_245_1122
timestamp 1636968456
transform 1 0 104328 0 -1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_245_1134
timestamp 1636968456
transform 1 0 105432 0 -1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_245_1146
timestamp 1636968456
transform 1 0 106536 0 -1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_245_1158
timestamp 1
transform 1 0 107640 0 -1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_245_1166
timestamp 1
transform 1 0 108376 0 -1 136000
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_246_3
timestamp 1636968456
transform 1 0 1380 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_15
timestamp 1636968456
transform 1 0 2484 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_246_27
timestamp 1
transform 1 0 3588 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_29
timestamp 1636968456
transform 1 0 3772 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_41
timestamp 1636968456
transform 1 0 4876 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_53
timestamp 1
transform 1 0 5980 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_57
timestamp 1636968456
transform 1 0 6348 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_69
timestamp 1636968456
transform 1 0 7452 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_81
timestamp 1
transform 1 0 8556 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_85
timestamp 1636968456
transform 1 0 8924 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_97
timestamp 1636968456
transform 1 0 10028 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_109
timestamp 1
transform 1 0 11132 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_113
timestamp 1636968456
transform 1 0 11500 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_125
timestamp 1636968456
transform 1 0 12604 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_137
timestamp 1
transform 1 0 13708 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_141
timestamp 1636968456
transform 1 0 14076 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_153
timestamp 1636968456
transform 1 0 15180 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_165
timestamp 1
transform 1 0 16284 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_169
timestamp 1636968456
transform 1 0 16652 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_181
timestamp 1636968456
transform 1 0 17756 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_193
timestamp 1
transform 1 0 18860 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_197
timestamp 1636968456
transform 1 0 19228 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_209
timestamp 1636968456
transform 1 0 20332 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_221
timestamp 1
transform 1 0 21436 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_225
timestamp 1636968456
transform 1 0 21804 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_237
timestamp 1636968456
transform 1 0 22908 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_249
timestamp 1
transform 1 0 24012 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_253
timestamp 1636968456
transform 1 0 24380 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_265
timestamp 1636968456
transform 1 0 25484 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_277
timestamp 1
transform 1 0 26588 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_281
timestamp 1636968456
transform 1 0 26956 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_293
timestamp 1636968456
transform 1 0 28060 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_305
timestamp 1
transform 1 0 29164 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_309
timestamp 1636968456
transform 1 0 29532 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_321
timestamp 1636968456
transform 1 0 30636 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_333
timestamp 1
transform 1 0 31740 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_337
timestamp 1636968456
transform 1 0 32108 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_349
timestamp 1636968456
transform 1 0 33212 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_361
timestamp 1
transform 1 0 34316 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_365
timestamp 1636968456
transform 1 0 34684 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_377
timestamp 1
transform 1 0 35788 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_246_382
timestamp 1
transform 1 0 36248 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_246_390
timestamp 1
transform 1 0 36984 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_246_393
timestamp 1
transform 1 0 37260 0 1 136000
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_246_407
timestamp 1636968456
transform 1 0 38548 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_246_419
timestamp 1
transform 1 0 39652 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_246_421
timestamp 1
transform 1 0 39836 0 1 136000
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_246_427
timestamp 1
transform 1 0 40388 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_434
timestamp 1636968456
transform 1 0 41032 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_246_446
timestamp 1
transform 1 0 42136 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_246_449
timestamp 1
transform 1 0 42412 0 1 136000
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_246_459
timestamp 1636968456
transform 1 0 43332 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_246_471
timestamp 1
transform 1 0 44436 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_246_475
timestamp 1
transform 1 0 44804 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_246_477
timestamp 1
transform 1 0 44988 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_484
timestamp 1636968456
transform 1 0 45632 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_496
timestamp 1
transform 1 0 46736 0 1 136000
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_246_511
timestamp 1636968456
transform 1 0 48116 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_523
timestamp 1
transform 1 0 49220 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_246_531
timestamp 1
transform 1 0 49956 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_533
timestamp 1636968456
transform 1 0 50140 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_545
timestamp 1636968456
transform 1 0 51244 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_557
timestamp 1
transform 1 0 52348 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_246_561
timestamp 1
transform 1 0 52716 0 1 136000
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_246_575
timestamp 1636968456
transform 1 0 54004 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_246_587
timestamp 1
transform 1 0 55108 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_246_589
timestamp 1
transform 1 0 55292 0 1 136000
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_246_599
timestamp 1636968456
transform 1 0 56212 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_246_611
timestamp 1
transform 1 0 57316 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_246_615
timestamp 1
transform 1 0 57684 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_246_617
timestamp 1
transform 1 0 57868 0 1 136000
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_246_625
timestamp 1636968456
transform 1 0 58604 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_246_637
timestamp 1
transform 1 0 59708 0 1 136000
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_246_643
timestamp 1
transform 1 0 60260 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_246_645
timestamp 1
transform 1 0 60444 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_652
timestamp 1636968456
transform 1 0 61088 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_664
timestamp 1
transform 1 0 62192 0 1 136000
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_246_679
timestamp 1636968456
transform 1 0 63572 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_246_691
timestamp 1
transform 1 0 64676 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_246_699
timestamp 1
transform 1 0 65412 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_701
timestamp 1636968456
transform 1 0 65596 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_713
timestamp 1
transform 1 0 66700 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_246_727
timestamp 1
transform 1 0 67988 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_729
timestamp 1636968456
transform 1 0 68172 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_246_741
timestamp 1
transform 1 0 69276 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_246_751
timestamp 1
transform 1 0 70196 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_246_755
timestamp 1
transform 1 0 70564 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_757
timestamp 1636968456
transform 1 0 70748 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_246_769
timestamp 1
transform 1 0 71852 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_246_777
timestamp 1
transform 1 0 72588 0 1 136000
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_246_783
timestamp 1
transform 1 0 73140 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_246_785
timestamp 1
transform 1 0 73324 0 1 136000
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_246_799
timestamp 1636968456
transform 1 0 74612 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_246_811
timestamp 1
transform 1 0 75716 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_813
timestamp 1636968456
transform 1 0 75900 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_825
timestamp 1636968456
transform 1 0 77004 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_837
timestamp 1
transform 1 0 78108 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_841
timestamp 1636968456
transform 1 0 78476 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_853
timestamp 1636968456
transform 1 0 79580 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_865
timestamp 1
transform 1 0 80684 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_869
timestamp 1636968456
transform 1 0 81052 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_881
timestamp 1636968456
transform 1 0 82156 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_893
timestamp 1
transform 1 0 83260 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_897
timestamp 1636968456
transform 1 0 83628 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_909
timestamp 1636968456
transform 1 0 84732 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_921
timestamp 1
transform 1 0 85836 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_246_927
timestamp 1
transform 1 0 86388 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_246_935
timestamp 1
transform 1 0 87124 0 1 136000
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_246_939
timestamp 1636968456
transform 1 0 87492 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_246_951
timestamp 1
transform 1 0 88596 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_953
timestamp 1636968456
transform 1 0 88780 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_965
timestamp 1636968456
transform 1 0 89884 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_977
timestamp 1
transform 1 0 90988 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_981
timestamp 1636968456
transform 1 0 91356 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_993
timestamp 1636968456
transform 1 0 92460 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_1005
timestamp 1
transform 1 0 93564 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1009
timestamp 1636968456
transform 1 0 93932 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_1021
timestamp 1
transform 1 0 95036 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_246_1029
timestamp 1
transform 1 0 95772 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_246_1032
timestamp 1
transform 1 0 96048 0 1 136000
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1037
timestamp 1636968456
transform 1 0 96508 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1049
timestamp 1636968456
transform 1 0 97612 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_1061
timestamp 1
transform 1 0 98716 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1065
timestamp 1636968456
transform 1 0 99084 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1077
timestamp 1636968456
transform 1 0 100188 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_1089
timestamp 1
transform 1 0 101292 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1093
timestamp 1636968456
transform 1 0 101660 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1105
timestamp 1636968456
transform 1 0 102764 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_1117
timestamp 1
transform 1 0 103868 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1121
timestamp 1636968456
transform 1 0 104236 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1133
timestamp 1636968456
transform 1 0 105340 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_1145
timestamp 1
transform 1 0 106444 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1149
timestamp 1636968456
transform 1 0 106812 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_246_1161
timestamp 1
transform 1 0 107916 0 1 136000
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_246_1167
timestamp 1
transform 1 0 108468 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_3
timestamp 1636968456
transform 1 0 1380 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_15
timestamp 1636968456
transform 1 0 2484 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_27
timestamp 1636968456
transform 1 0 3588 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_39
timestamp 1636968456
transform 1 0 4692 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_247_51
timestamp 1
transform 1 0 5796 0 -1 137088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_247_55
timestamp 1
transform 1 0 6164 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_57
timestamp 1636968456
transform 1 0 6348 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_69
timestamp 1636968456
transform 1 0 7452 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_81
timestamp 1636968456
transform 1 0 8556 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_93
timestamp 1636968456
transform 1 0 9660 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_105
timestamp 1
transform 1 0 10764 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_111
timestamp 1
transform 1 0 11316 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_113
timestamp 1636968456
transform 1 0 11500 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_125
timestamp 1636968456
transform 1 0 12604 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_137
timestamp 1636968456
transform 1 0 13708 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_149
timestamp 1636968456
transform 1 0 14812 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_161
timestamp 1
transform 1 0 15916 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_167
timestamp 1
transform 1 0 16468 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_169
timestamp 1636968456
transform 1 0 16652 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_181
timestamp 1636968456
transform 1 0 17756 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_193
timestamp 1636968456
transform 1 0 18860 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_205
timestamp 1636968456
transform 1 0 19964 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_217
timestamp 1
transform 1 0 21068 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_223
timestamp 1
transform 1 0 21620 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_225
timestamp 1636968456
transform 1 0 21804 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_237
timestamp 1636968456
transform 1 0 22908 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_249
timestamp 1636968456
transform 1 0 24012 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_261
timestamp 1636968456
transform 1 0 25116 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_273
timestamp 1
transform 1 0 26220 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_279
timestamp 1
transform 1 0 26772 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_281
timestamp 1636968456
transform 1 0 26956 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_293
timestamp 1636968456
transform 1 0 28060 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_305
timestamp 1636968456
transform 1 0 29164 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_317
timestamp 1636968456
transform 1 0 30268 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_329
timestamp 1
transform 1 0 31372 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_335
timestamp 1
transform 1 0 31924 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_337
timestamp 1636968456
transform 1 0 32108 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_349
timestamp 1636968456
transform 1 0 33212 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_361
timestamp 1636968456
transform 1 0 34316 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_373
timestamp 1636968456
transform 1 0 35420 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_385
timestamp 1
transform 1 0 36524 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_391
timestamp 1
transform 1 0 37076 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_393
timestamp 1636968456
transform 1 0 37260 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_405
timestamp 1636968456
transform 1 0 38364 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_417
timestamp 1636968456
transform 1 0 39468 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_429
timestamp 1636968456
transform 1 0 40572 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_441
timestamp 1
transform 1 0 41676 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_447
timestamp 1
transform 1 0 42228 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_449
timestamp 1636968456
transform 1 0 42412 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_461
timestamp 1636968456
transform 1 0 43516 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_473
timestamp 1636968456
transform 1 0 44620 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_485
timestamp 1636968456
transform 1 0 45724 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_497
timestamp 1
transform 1 0 46828 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_503
timestamp 1
transform 1 0 47380 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_505
timestamp 1636968456
transform 1 0 47564 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_517
timestamp 1636968456
transform 1 0 48668 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_529
timestamp 1636968456
transform 1 0 49772 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_541
timestamp 1636968456
transform 1 0 50876 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_553
timestamp 1
transform 1 0 51980 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_559
timestamp 1
transform 1 0 52532 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_561
timestamp 1636968456
transform 1 0 52716 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_573
timestamp 1636968456
transform 1 0 53820 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_585
timestamp 1636968456
transform 1 0 54924 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_597
timestamp 1636968456
transform 1 0 56028 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_609
timestamp 1
transform 1 0 57132 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_615
timestamp 1
transform 1 0 57684 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_617
timestamp 1636968456
transform 1 0 57868 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_629
timestamp 1636968456
transform 1 0 58972 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_641
timestamp 1636968456
transform 1 0 60076 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_653
timestamp 1636968456
transform 1 0 61180 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_665
timestamp 1
transform 1 0 62284 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_671
timestamp 1
transform 1 0 62836 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_673
timestamp 1636968456
transform 1 0 63020 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_685
timestamp 1636968456
transform 1 0 64124 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_697
timestamp 1636968456
transform 1 0 65228 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_709
timestamp 1636968456
transform 1 0 66332 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_721
timestamp 1
transform 1 0 67436 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_727
timestamp 1
transform 1 0 67988 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_729
timestamp 1636968456
transform 1 0 68172 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_741
timestamp 1636968456
transform 1 0 69276 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_753
timestamp 1636968456
transform 1 0 70380 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_765
timestamp 1636968456
transform 1 0 71484 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_777
timestamp 1
transform 1 0 72588 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_783
timestamp 1
transform 1 0 73140 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_785
timestamp 1636968456
transform 1 0 73324 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_797
timestamp 1636968456
transform 1 0 74428 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_809
timestamp 1636968456
transform 1 0 75532 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_821
timestamp 1636968456
transform 1 0 76636 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_833
timestamp 1
transform 1 0 77740 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_839
timestamp 1
transform 1 0 78292 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_841
timestamp 1636968456
transform 1 0 78476 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_853
timestamp 1636968456
transform 1 0 79580 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_865
timestamp 1636968456
transform 1 0 80684 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_877
timestamp 1636968456
transform 1 0 81788 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_889
timestamp 1
transform 1 0 82892 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_895
timestamp 1
transform 1 0 83444 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_897
timestamp 1636968456
transform 1 0 83628 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_909
timestamp 1636968456
transform 1 0 84732 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_921
timestamp 1636968456
transform 1 0 85836 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_933
timestamp 1636968456
transform 1 0 86940 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_945
timestamp 1
transform 1 0 88044 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_951
timestamp 1
transform 1 0 88596 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_953
timestamp 1636968456
transform 1 0 88780 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_965
timestamp 1636968456
transform 1 0 89884 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_977
timestamp 1636968456
transform 1 0 90988 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_989
timestamp 1636968456
transform 1 0 92092 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_1001
timestamp 1
transform 1 0 93196 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_1007
timestamp 1
transform 1 0 93748 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1009
timestamp 1636968456
transform 1 0 93932 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1021
timestamp 1636968456
transform 1 0 95036 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1033
timestamp 1636968456
transform 1 0 96140 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1045
timestamp 1636968456
transform 1 0 97244 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_1057
timestamp 1
transform 1 0 98348 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_1063
timestamp 1
transform 1 0 98900 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1065
timestamp 1636968456
transform 1 0 99084 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1077
timestamp 1636968456
transform 1 0 100188 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1089
timestamp 1636968456
transform 1 0 101292 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1101
timestamp 1636968456
transform 1 0 102396 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_1113
timestamp 1
transform 1 0 103500 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_1119
timestamp 1
transform 1 0 104052 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1121
timestamp 1636968456
transform 1 0 104236 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1133
timestamp 1636968456
transform 1 0 105340 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1145
timestamp 1636968456
transform 1 0 106444 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_247_1157
timestamp 1
transform 1 0 107548 0 -1 137088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_247_1165
timestamp 1
transform 1 0 108284 0 -1 137088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_248_3
timestamp 1636968456
transform 1 0 1380 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_15
timestamp 1636968456
transform 1 0 2484 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_248_27
timestamp 1
transform 1 0 3588 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_29
timestamp 1636968456
transform 1 0 3772 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_41
timestamp 1636968456
transform 1 0 4876 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_53
timestamp 1636968456
transform 1 0 5980 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_65
timestamp 1636968456
transform 1 0 7084 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_77
timestamp 1
transform 1 0 8188 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_83
timestamp 1
transform 1 0 8740 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_85
timestamp 1636968456
transform 1 0 8924 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_97
timestamp 1636968456
transform 1 0 10028 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_109
timestamp 1636968456
transform 1 0 11132 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_121
timestamp 1636968456
transform 1 0 12236 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_133
timestamp 1
transform 1 0 13340 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_139
timestamp 1
transform 1 0 13892 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_141
timestamp 1636968456
transform 1 0 14076 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_153
timestamp 1636968456
transform 1 0 15180 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_165
timestamp 1636968456
transform 1 0 16284 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_177
timestamp 1636968456
transform 1 0 17388 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_189
timestamp 1
transform 1 0 18492 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_195
timestamp 1
transform 1 0 19044 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_197
timestamp 1636968456
transform 1 0 19228 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_209
timestamp 1636968456
transform 1 0 20332 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_221
timestamp 1636968456
transform 1 0 21436 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_233
timestamp 1636968456
transform 1 0 22540 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_245
timestamp 1
transform 1 0 23644 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_251
timestamp 1
transform 1 0 24196 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_253
timestamp 1636968456
transform 1 0 24380 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_265
timestamp 1636968456
transform 1 0 25484 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_277
timestamp 1636968456
transform 1 0 26588 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_289
timestamp 1636968456
transform 1 0 27692 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_301
timestamp 1
transform 1 0 28796 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_307
timestamp 1
transform 1 0 29348 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_309
timestamp 1636968456
transform 1 0 29532 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_321
timestamp 1636968456
transform 1 0 30636 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_333
timestamp 1636968456
transform 1 0 31740 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_345
timestamp 1636968456
transform 1 0 32844 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_357
timestamp 1
transform 1 0 33948 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_363
timestamp 1
transform 1 0 34500 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_365
timestamp 1636968456
transform 1 0 34684 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_377
timestamp 1636968456
transform 1 0 35788 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_389
timestamp 1636968456
transform 1 0 36892 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_401
timestamp 1636968456
transform 1 0 37996 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_413
timestamp 1
transform 1 0 39100 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_419
timestamp 1
transform 1 0 39652 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_421
timestamp 1636968456
transform 1 0 39836 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_433
timestamp 1636968456
transform 1 0 40940 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_445
timestamp 1636968456
transform 1 0 42044 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_457
timestamp 1636968456
transform 1 0 43148 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_469
timestamp 1
transform 1 0 44252 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_475
timestamp 1
transform 1 0 44804 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_477
timestamp 1636968456
transform 1 0 44988 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_489
timestamp 1636968456
transform 1 0 46092 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_501
timestamp 1636968456
transform 1 0 47196 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_513
timestamp 1636968456
transform 1 0 48300 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_525
timestamp 1
transform 1 0 49404 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_531
timestamp 1
transform 1 0 49956 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_533
timestamp 1636968456
transform 1 0 50140 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_545
timestamp 1636968456
transform 1 0 51244 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_557
timestamp 1636968456
transform 1 0 52348 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_569
timestamp 1636968456
transform 1 0 53452 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_581
timestamp 1
transform 1 0 54556 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_587
timestamp 1
transform 1 0 55108 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_589
timestamp 1636968456
transform 1 0 55292 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_601
timestamp 1636968456
transform 1 0 56396 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_613
timestamp 1636968456
transform 1 0 57500 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_625
timestamp 1636968456
transform 1 0 58604 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_637
timestamp 1
transform 1 0 59708 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_643
timestamp 1
transform 1 0 60260 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_645
timestamp 1636968456
transform 1 0 60444 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_657
timestamp 1636968456
transform 1 0 61548 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_669
timestamp 1636968456
transform 1 0 62652 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_681
timestamp 1636968456
transform 1 0 63756 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_693
timestamp 1
transform 1 0 64860 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_699
timestamp 1
transform 1 0 65412 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_701
timestamp 1636968456
transform 1 0 65596 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_713
timestamp 1636968456
transform 1 0 66700 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_725
timestamp 1636968456
transform 1 0 67804 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_737
timestamp 1636968456
transform 1 0 68908 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_749
timestamp 1
transform 1 0 70012 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_755
timestamp 1
transform 1 0 70564 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_757
timestamp 1636968456
transform 1 0 70748 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_769
timestamp 1636968456
transform 1 0 71852 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_781
timestamp 1636968456
transform 1 0 72956 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_793
timestamp 1636968456
transform 1 0 74060 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_805
timestamp 1
transform 1 0 75164 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_811
timestamp 1
transform 1 0 75716 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_813
timestamp 1636968456
transform 1 0 75900 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_825
timestamp 1636968456
transform 1 0 77004 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_837
timestamp 1636968456
transform 1 0 78108 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_849
timestamp 1636968456
transform 1 0 79212 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_861
timestamp 1
transform 1 0 80316 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_867
timestamp 1
transform 1 0 80868 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_869
timestamp 1636968456
transform 1 0 81052 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_881
timestamp 1636968456
transform 1 0 82156 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_893
timestamp 1636968456
transform 1 0 83260 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_905
timestamp 1636968456
transform 1 0 84364 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_917
timestamp 1
transform 1 0 85468 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_923
timestamp 1
transform 1 0 86020 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_925
timestamp 1636968456
transform 1 0 86204 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_937
timestamp 1636968456
transform 1 0 87308 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_949
timestamp 1636968456
transform 1 0 88412 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_961
timestamp 1636968456
transform 1 0 89516 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_973
timestamp 1
transform 1 0 90620 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_979
timestamp 1
transform 1 0 91172 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_981
timestamp 1636968456
transform 1 0 91356 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_993
timestamp 1636968456
transform 1 0 92460 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1005
timestamp 1636968456
transform 1 0 93564 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1017
timestamp 1636968456
transform 1 0 94668 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_1029
timestamp 1
transform 1 0 95772 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_1035
timestamp 1
transform 1 0 96324 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1037
timestamp 1636968456
transform 1 0 96508 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1049
timestamp 1636968456
transform 1 0 97612 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1061
timestamp 1636968456
transform 1 0 98716 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1073
timestamp 1636968456
transform 1 0 99820 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_1085
timestamp 1
transform 1 0 100924 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_1091
timestamp 1
transform 1 0 101476 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1093
timestamp 1636968456
transform 1 0 101660 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1105
timestamp 1636968456
transform 1 0 102764 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1117
timestamp 1636968456
transform 1 0 103868 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1129
timestamp 1636968456
transform 1 0 104972 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_1141
timestamp 1
transform 1 0 106076 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_1147
timestamp 1
transform 1 0 106628 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1149
timestamp 1636968456
transform 1 0 106812 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_1161
timestamp 1
transform 1 0 107916 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_1167
timestamp 1
transform 1 0 108468 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_3
timestamp 1636968456
transform 1 0 1380 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_15
timestamp 1636968456
transform 1 0 2484 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_27
timestamp 1636968456
transform 1 0 3588 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_39
timestamp 1636968456
transform 1 0 4692 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_249_51
timestamp 1
transform 1 0 5796 0 -1 138176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_249_55
timestamp 1
transform 1 0 6164 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_57
timestamp 1636968456
transform 1 0 6348 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_69
timestamp 1636968456
transform 1 0 7452 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_81
timestamp 1636968456
transform 1 0 8556 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_93
timestamp 1636968456
transform 1 0 9660 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_105
timestamp 1
transform 1 0 10764 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_111
timestamp 1
transform 1 0 11316 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_113
timestamp 1636968456
transform 1 0 11500 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_125
timestamp 1636968456
transform 1 0 12604 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_137
timestamp 1636968456
transform 1 0 13708 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_149
timestamp 1636968456
transform 1 0 14812 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_161
timestamp 1
transform 1 0 15916 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_167
timestamp 1
transform 1 0 16468 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_169
timestamp 1636968456
transform 1 0 16652 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_181
timestamp 1636968456
transform 1 0 17756 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_193
timestamp 1636968456
transform 1 0 18860 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_205
timestamp 1636968456
transform 1 0 19964 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_217
timestamp 1
transform 1 0 21068 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_223
timestamp 1
transform 1 0 21620 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_225
timestamp 1636968456
transform 1 0 21804 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_237
timestamp 1636968456
transform 1 0 22908 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_249
timestamp 1636968456
transform 1 0 24012 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_261
timestamp 1636968456
transform 1 0 25116 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_273
timestamp 1
transform 1 0 26220 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_279
timestamp 1
transform 1 0 26772 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_281
timestamp 1636968456
transform 1 0 26956 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_293
timestamp 1636968456
transform 1 0 28060 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_305
timestamp 1636968456
transform 1 0 29164 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_317
timestamp 1636968456
transform 1 0 30268 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_329
timestamp 1
transform 1 0 31372 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_335
timestamp 1
transform 1 0 31924 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_337
timestamp 1636968456
transform 1 0 32108 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_349
timestamp 1636968456
transform 1 0 33212 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_361
timestamp 1636968456
transform 1 0 34316 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_373
timestamp 1636968456
transform 1 0 35420 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_385
timestamp 1
transform 1 0 36524 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_391
timestamp 1
transform 1 0 37076 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_393
timestamp 1636968456
transform 1 0 37260 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_405
timestamp 1636968456
transform 1 0 38364 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_417
timestamp 1636968456
transform 1 0 39468 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_429
timestamp 1636968456
transform 1 0 40572 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_441
timestamp 1
transform 1 0 41676 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_447
timestamp 1
transform 1 0 42228 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_449
timestamp 1636968456
transform 1 0 42412 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_461
timestamp 1636968456
transform 1 0 43516 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_473
timestamp 1636968456
transform 1 0 44620 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_485
timestamp 1636968456
transform 1 0 45724 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_497
timestamp 1
transform 1 0 46828 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_503
timestamp 1
transform 1 0 47380 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_505
timestamp 1636968456
transform 1 0 47564 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_517
timestamp 1636968456
transform 1 0 48668 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_529
timestamp 1636968456
transform 1 0 49772 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_541
timestamp 1636968456
transform 1 0 50876 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_553
timestamp 1
transform 1 0 51980 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_559
timestamp 1
transform 1 0 52532 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_561
timestamp 1636968456
transform 1 0 52716 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_573
timestamp 1636968456
transform 1 0 53820 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_585
timestamp 1636968456
transform 1 0 54924 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_597
timestamp 1636968456
transform 1 0 56028 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_609
timestamp 1
transform 1 0 57132 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_615
timestamp 1
transform 1 0 57684 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_617
timestamp 1636968456
transform 1 0 57868 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_629
timestamp 1636968456
transform 1 0 58972 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_641
timestamp 1636968456
transform 1 0 60076 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_653
timestamp 1636968456
transform 1 0 61180 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_665
timestamp 1
transform 1 0 62284 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_671
timestamp 1
transform 1 0 62836 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_673
timestamp 1636968456
transform 1 0 63020 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_685
timestamp 1636968456
transform 1 0 64124 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_697
timestamp 1636968456
transform 1 0 65228 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_709
timestamp 1636968456
transform 1 0 66332 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_721
timestamp 1
transform 1 0 67436 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_727
timestamp 1
transform 1 0 67988 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_729
timestamp 1636968456
transform 1 0 68172 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_741
timestamp 1636968456
transform 1 0 69276 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_753
timestamp 1636968456
transform 1 0 70380 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_765
timestamp 1636968456
transform 1 0 71484 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_777
timestamp 1
transform 1 0 72588 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_783
timestamp 1
transform 1 0 73140 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_785
timestamp 1636968456
transform 1 0 73324 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_797
timestamp 1636968456
transform 1 0 74428 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_809
timestamp 1636968456
transform 1 0 75532 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_821
timestamp 1636968456
transform 1 0 76636 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_833
timestamp 1
transform 1 0 77740 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_839
timestamp 1
transform 1 0 78292 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_841
timestamp 1636968456
transform 1 0 78476 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_853
timestamp 1636968456
transform 1 0 79580 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_865
timestamp 1636968456
transform 1 0 80684 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_877
timestamp 1636968456
transform 1 0 81788 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_889
timestamp 1
transform 1 0 82892 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_895
timestamp 1
transform 1 0 83444 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_897
timestamp 1636968456
transform 1 0 83628 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_909
timestamp 1636968456
transform 1 0 84732 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_921
timestamp 1636968456
transform 1 0 85836 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_933
timestamp 1636968456
transform 1 0 86940 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_945
timestamp 1
transform 1 0 88044 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_951
timestamp 1
transform 1 0 88596 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_953
timestamp 1636968456
transform 1 0 88780 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_965
timestamp 1636968456
transform 1 0 89884 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_977
timestamp 1636968456
transform 1 0 90988 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_989
timestamp 1636968456
transform 1 0 92092 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_1001
timestamp 1
transform 1 0 93196 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_1007
timestamp 1
transform 1 0 93748 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1009
timestamp 1636968456
transform 1 0 93932 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1021
timestamp 1636968456
transform 1 0 95036 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1033
timestamp 1636968456
transform 1 0 96140 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1045
timestamp 1636968456
transform 1 0 97244 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_1057
timestamp 1
transform 1 0 98348 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_1063
timestamp 1
transform 1 0 98900 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1065
timestamp 1636968456
transform 1 0 99084 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1077
timestamp 1636968456
transform 1 0 100188 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1089
timestamp 1636968456
transform 1 0 101292 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1101
timestamp 1636968456
transform 1 0 102396 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_1113
timestamp 1
transform 1 0 103500 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_1119
timestamp 1
transform 1 0 104052 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1121
timestamp 1636968456
transform 1 0 104236 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1133
timestamp 1636968456
transform 1 0 105340 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1145
timestamp 1636968456
transform 1 0 106444 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_249_1157
timestamp 1
transform 1 0 107548 0 -1 138176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_249_1165
timestamp 1
transform 1 0 108284 0 -1 138176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_250_3
timestamp 1636968456
transform 1 0 1380 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_15
timestamp 1636968456
transform 1 0 2484 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_250_27
timestamp 1
transform 1 0 3588 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_29
timestamp 1636968456
transform 1 0 3772 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_41
timestamp 1636968456
transform 1 0 4876 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_53
timestamp 1636968456
transform 1 0 5980 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_65
timestamp 1636968456
transform 1 0 7084 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_77
timestamp 1
transform 1 0 8188 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_83
timestamp 1
transform 1 0 8740 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_85
timestamp 1636968456
transform 1 0 8924 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_97
timestamp 1636968456
transform 1 0 10028 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_109
timestamp 1636968456
transform 1 0 11132 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_121
timestamp 1636968456
transform 1 0 12236 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_133
timestamp 1
transform 1 0 13340 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_139
timestamp 1
transform 1 0 13892 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_141
timestamp 1636968456
transform 1 0 14076 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_153
timestamp 1636968456
transform 1 0 15180 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_165
timestamp 1636968456
transform 1 0 16284 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_177
timestamp 1636968456
transform 1 0 17388 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_189
timestamp 1
transform 1 0 18492 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_195
timestamp 1
transform 1 0 19044 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_197
timestamp 1636968456
transform 1 0 19228 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_209
timestamp 1636968456
transform 1 0 20332 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_221
timestamp 1636968456
transform 1 0 21436 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_233
timestamp 1636968456
transform 1 0 22540 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_245
timestamp 1
transform 1 0 23644 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_251
timestamp 1
transform 1 0 24196 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_253
timestamp 1636968456
transform 1 0 24380 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_265
timestamp 1636968456
transform 1 0 25484 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_277
timestamp 1636968456
transform 1 0 26588 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_289
timestamp 1636968456
transform 1 0 27692 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_301
timestamp 1
transform 1 0 28796 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_307
timestamp 1
transform 1 0 29348 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_309
timestamp 1636968456
transform 1 0 29532 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_321
timestamp 1636968456
transform 1 0 30636 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_333
timestamp 1636968456
transform 1 0 31740 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_345
timestamp 1636968456
transform 1 0 32844 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_357
timestamp 1
transform 1 0 33948 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_363
timestamp 1
transform 1 0 34500 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_365
timestamp 1636968456
transform 1 0 34684 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_377
timestamp 1636968456
transform 1 0 35788 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_389
timestamp 1636968456
transform 1 0 36892 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_401
timestamp 1636968456
transform 1 0 37996 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_413
timestamp 1
transform 1 0 39100 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_419
timestamp 1
transform 1 0 39652 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_421
timestamp 1636968456
transform 1 0 39836 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_433
timestamp 1636968456
transform 1 0 40940 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_445
timestamp 1636968456
transform 1 0 42044 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_457
timestamp 1636968456
transform 1 0 43148 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_469
timestamp 1
transform 1 0 44252 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_475
timestamp 1
transform 1 0 44804 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_477
timestamp 1636968456
transform 1 0 44988 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_489
timestamp 1636968456
transform 1 0 46092 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_501
timestamp 1636968456
transform 1 0 47196 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_513
timestamp 1636968456
transform 1 0 48300 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_525
timestamp 1
transform 1 0 49404 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_531
timestamp 1
transform 1 0 49956 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_533
timestamp 1636968456
transform 1 0 50140 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_545
timestamp 1636968456
transform 1 0 51244 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_557
timestamp 1636968456
transform 1 0 52348 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_569
timestamp 1636968456
transform 1 0 53452 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_581
timestamp 1
transform 1 0 54556 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_587
timestamp 1
transform 1 0 55108 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_589
timestamp 1636968456
transform 1 0 55292 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_601
timestamp 1636968456
transform 1 0 56396 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_613
timestamp 1636968456
transform 1 0 57500 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_625
timestamp 1636968456
transform 1 0 58604 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_637
timestamp 1
transform 1 0 59708 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_643
timestamp 1
transform 1 0 60260 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_645
timestamp 1636968456
transform 1 0 60444 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_657
timestamp 1636968456
transform 1 0 61548 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_669
timestamp 1636968456
transform 1 0 62652 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_681
timestamp 1636968456
transform 1 0 63756 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_693
timestamp 1
transform 1 0 64860 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_699
timestamp 1
transform 1 0 65412 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_701
timestamp 1636968456
transform 1 0 65596 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_713
timestamp 1636968456
transform 1 0 66700 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_725
timestamp 1636968456
transform 1 0 67804 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_737
timestamp 1636968456
transform 1 0 68908 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_749
timestamp 1
transform 1 0 70012 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_755
timestamp 1
transform 1 0 70564 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_757
timestamp 1636968456
transform 1 0 70748 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_769
timestamp 1636968456
transform 1 0 71852 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_781
timestamp 1636968456
transform 1 0 72956 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_793
timestamp 1636968456
transform 1 0 74060 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_805
timestamp 1
transform 1 0 75164 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_811
timestamp 1
transform 1 0 75716 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_813
timestamp 1636968456
transform 1 0 75900 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_825
timestamp 1636968456
transform 1 0 77004 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_837
timestamp 1636968456
transform 1 0 78108 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_849
timestamp 1636968456
transform 1 0 79212 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_861
timestamp 1
transform 1 0 80316 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_867
timestamp 1
transform 1 0 80868 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_869
timestamp 1636968456
transform 1 0 81052 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_881
timestamp 1636968456
transform 1 0 82156 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_893
timestamp 1636968456
transform 1 0 83260 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_905
timestamp 1636968456
transform 1 0 84364 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_917
timestamp 1
transform 1 0 85468 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_923
timestamp 1
transform 1 0 86020 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_925
timestamp 1636968456
transform 1 0 86204 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_937
timestamp 1636968456
transform 1 0 87308 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_949
timestamp 1636968456
transform 1 0 88412 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_961
timestamp 1636968456
transform 1 0 89516 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_973
timestamp 1
transform 1 0 90620 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_979
timestamp 1
transform 1 0 91172 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_981
timestamp 1636968456
transform 1 0 91356 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_993
timestamp 1636968456
transform 1 0 92460 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1005
timestamp 1636968456
transform 1 0 93564 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1017
timestamp 1636968456
transform 1 0 94668 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_1029
timestamp 1
transform 1 0 95772 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_1035
timestamp 1
transform 1 0 96324 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1037
timestamp 1636968456
transform 1 0 96508 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1049
timestamp 1636968456
transform 1 0 97612 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1061
timestamp 1636968456
transform 1 0 98716 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1073
timestamp 1636968456
transform 1 0 99820 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_1085
timestamp 1
transform 1 0 100924 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_1091
timestamp 1
transform 1 0 101476 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1093
timestamp 1636968456
transform 1 0 101660 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1105
timestamp 1636968456
transform 1 0 102764 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1117
timestamp 1636968456
transform 1 0 103868 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1129
timestamp 1636968456
transform 1 0 104972 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_1141
timestamp 1
transform 1 0 106076 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_1147
timestamp 1
transform 1 0 106628 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1149
timestamp 1636968456
transform 1 0 106812 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_1161
timestamp 1
transform 1 0 107916 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_1167
timestamp 1
transform 1 0 108468 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_3
timestamp 1636968456
transform 1 0 1380 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_15
timestamp 1636968456
transform 1 0 2484 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_27
timestamp 1636968456
transform 1 0 3588 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_39
timestamp 1636968456
transform 1 0 4692 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_251_51
timestamp 1
transform 1 0 5796 0 -1 139264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_251_55
timestamp 1
transform 1 0 6164 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_57
timestamp 1636968456
transform 1 0 6348 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_69
timestamp 1636968456
transform 1 0 7452 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_81
timestamp 1636968456
transform 1 0 8556 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_93
timestamp 1636968456
transform 1 0 9660 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_105
timestamp 1
transform 1 0 10764 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_111
timestamp 1
transform 1 0 11316 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_113
timestamp 1636968456
transform 1 0 11500 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_125
timestamp 1636968456
transform 1 0 12604 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_137
timestamp 1636968456
transform 1 0 13708 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_149
timestamp 1636968456
transform 1 0 14812 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_161
timestamp 1
transform 1 0 15916 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_167
timestamp 1
transform 1 0 16468 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_169
timestamp 1636968456
transform 1 0 16652 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_181
timestamp 1636968456
transform 1 0 17756 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_193
timestamp 1636968456
transform 1 0 18860 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_205
timestamp 1636968456
transform 1 0 19964 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_217
timestamp 1
transform 1 0 21068 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_223
timestamp 1
transform 1 0 21620 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_225
timestamp 1636968456
transform 1 0 21804 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_237
timestamp 1636968456
transform 1 0 22908 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_249
timestamp 1636968456
transform 1 0 24012 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_261
timestamp 1636968456
transform 1 0 25116 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_273
timestamp 1
transform 1 0 26220 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_279
timestamp 1
transform 1 0 26772 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_281
timestamp 1636968456
transform 1 0 26956 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_293
timestamp 1636968456
transform 1 0 28060 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_305
timestamp 1636968456
transform 1 0 29164 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_317
timestamp 1636968456
transform 1 0 30268 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_329
timestamp 1
transform 1 0 31372 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_335
timestamp 1
transform 1 0 31924 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_337
timestamp 1636968456
transform 1 0 32108 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_349
timestamp 1636968456
transform 1 0 33212 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_361
timestamp 1636968456
transform 1 0 34316 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_373
timestamp 1636968456
transform 1 0 35420 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_385
timestamp 1
transform 1 0 36524 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_391
timestamp 1
transform 1 0 37076 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_393
timestamp 1636968456
transform 1 0 37260 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_405
timestamp 1636968456
transform 1 0 38364 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_417
timestamp 1636968456
transform 1 0 39468 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_429
timestamp 1636968456
transform 1 0 40572 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_441
timestamp 1
transform 1 0 41676 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_447
timestamp 1
transform 1 0 42228 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_449
timestamp 1636968456
transform 1 0 42412 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_461
timestamp 1636968456
transform 1 0 43516 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_473
timestamp 1636968456
transform 1 0 44620 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_485
timestamp 1636968456
transform 1 0 45724 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_497
timestamp 1
transform 1 0 46828 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_503
timestamp 1
transform 1 0 47380 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_505
timestamp 1636968456
transform 1 0 47564 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_517
timestamp 1636968456
transform 1 0 48668 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_529
timestamp 1636968456
transform 1 0 49772 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_541
timestamp 1636968456
transform 1 0 50876 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_553
timestamp 1
transform 1 0 51980 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_559
timestamp 1
transform 1 0 52532 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_561
timestamp 1636968456
transform 1 0 52716 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_573
timestamp 1636968456
transform 1 0 53820 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_585
timestamp 1636968456
transform 1 0 54924 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_597
timestamp 1636968456
transform 1 0 56028 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_609
timestamp 1
transform 1 0 57132 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_615
timestamp 1
transform 1 0 57684 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_617
timestamp 1636968456
transform 1 0 57868 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_629
timestamp 1636968456
transform 1 0 58972 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_641
timestamp 1636968456
transform 1 0 60076 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_653
timestamp 1636968456
transform 1 0 61180 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_665
timestamp 1
transform 1 0 62284 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_671
timestamp 1
transform 1 0 62836 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_673
timestamp 1636968456
transform 1 0 63020 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_685
timestamp 1636968456
transform 1 0 64124 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_697
timestamp 1636968456
transform 1 0 65228 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_709
timestamp 1636968456
transform 1 0 66332 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_721
timestamp 1
transform 1 0 67436 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_727
timestamp 1
transform 1 0 67988 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_729
timestamp 1636968456
transform 1 0 68172 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_741
timestamp 1636968456
transform 1 0 69276 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_753
timestamp 1636968456
transform 1 0 70380 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_765
timestamp 1636968456
transform 1 0 71484 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_777
timestamp 1
transform 1 0 72588 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_783
timestamp 1
transform 1 0 73140 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_785
timestamp 1636968456
transform 1 0 73324 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_797
timestamp 1636968456
transform 1 0 74428 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_809
timestamp 1636968456
transform 1 0 75532 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_821
timestamp 1636968456
transform 1 0 76636 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_833
timestamp 1
transform 1 0 77740 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_839
timestamp 1
transform 1 0 78292 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_841
timestamp 1636968456
transform 1 0 78476 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_853
timestamp 1636968456
transform 1 0 79580 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_865
timestamp 1636968456
transform 1 0 80684 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_877
timestamp 1636968456
transform 1 0 81788 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_889
timestamp 1
transform 1 0 82892 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_895
timestamp 1
transform 1 0 83444 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_897
timestamp 1636968456
transform 1 0 83628 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_909
timestamp 1636968456
transform 1 0 84732 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_921
timestamp 1636968456
transform 1 0 85836 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_933
timestamp 1636968456
transform 1 0 86940 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_945
timestamp 1
transform 1 0 88044 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_951
timestamp 1
transform 1 0 88596 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_953
timestamp 1636968456
transform 1 0 88780 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_965
timestamp 1636968456
transform 1 0 89884 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_977
timestamp 1636968456
transform 1 0 90988 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_989
timestamp 1636968456
transform 1 0 92092 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_1001
timestamp 1
transform 1 0 93196 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_1007
timestamp 1
transform 1 0 93748 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1009
timestamp 1636968456
transform 1 0 93932 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1021
timestamp 1636968456
transform 1 0 95036 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1033
timestamp 1636968456
transform 1 0 96140 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1045
timestamp 1636968456
transform 1 0 97244 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_1057
timestamp 1
transform 1 0 98348 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_1063
timestamp 1
transform 1 0 98900 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1065
timestamp 1636968456
transform 1 0 99084 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1077
timestamp 1636968456
transform 1 0 100188 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1089
timestamp 1636968456
transform 1 0 101292 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1101
timestamp 1636968456
transform 1 0 102396 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_1113
timestamp 1
transform 1 0 103500 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_1119
timestamp 1
transform 1 0 104052 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1121
timestamp 1636968456
transform 1 0 104236 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1133
timestamp 1636968456
transform 1 0 105340 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1145
timestamp 1636968456
transform 1 0 106444 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_251_1157
timestamp 1
transform 1 0 107548 0 -1 139264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_251_1165
timestamp 1
transform 1 0 108284 0 -1 139264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_252_3
timestamp 1636968456
transform 1 0 1380 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_15
timestamp 1636968456
transform 1 0 2484 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_252_27
timestamp 1
transform 1 0 3588 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_29
timestamp 1636968456
transform 1 0 3772 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_41
timestamp 1636968456
transform 1 0 4876 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_53
timestamp 1636968456
transform 1 0 5980 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_65
timestamp 1636968456
transform 1 0 7084 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_77
timestamp 1
transform 1 0 8188 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_83
timestamp 1
transform 1 0 8740 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_85
timestamp 1636968456
transform 1 0 8924 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_97
timestamp 1636968456
transform 1 0 10028 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_109
timestamp 1636968456
transform 1 0 11132 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_121
timestamp 1636968456
transform 1 0 12236 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_133
timestamp 1
transform 1 0 13340 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_139
timestamp 1
transform 1 0 13892 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_141
timestamp 1636968456
transform 1 0 14076 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_153
timestamp 1636968456
transform 1 0 15180 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_165
timestamp 1636968456
transform 1 0 16284 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_177
timestamp 1636968456
transform 1 0 17388 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_189
timestamp 1
transform 1 0 18492 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_195
timestamp 1
transform 1 0 19044 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_197
timestamp 1636968456
transform 1 0 19228 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_209
timestamp 1636968456
transform 1 0 20332 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_221
timestamp 1636968456
transform 1 0 21436 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_233
timestamp 1636968456
transform 1 0 22540 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_245
timestamp 1
transform 1 0 23644 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_251
timestamp 1
transform 1 0 24196 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_253
timestamp 1636968456
transform 1 0 24380 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_265
timestamp 1636968456
transform 1 0 25484 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_277
timestamp 1636968456
transform 1 0 26588 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_289
timestamp 1636968456
transform 1 0 27692 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_301
timestamp 1
transform 1 0 28796 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_307
timestamp 1
transform 1 0 29348 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_309
timestamp 1636968456
transform 1 0 29532 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_321
timestamp 1636968456
transform 1 0 30636 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_333
timestamp 1636968456
transform 1 0 31740 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_345
timestamp 1636968456
transform 1 0 32844 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_357
timestamp 1
transform 1 0 33948 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_363
timestamp 1
transform 1 0 34500 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_365
timestamp 1636968456
transform 1 0 34684 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_377
timestamp 1636968456
transform 1 0 35788 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_389
timestamp 1636968456
transform 1 0 36892 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_401
timestamp 1636968456
transform 1 0 37996 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_413
timestamp 1
transform 1 0 39100 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_419
timestamp 1
transform 1 0 39652 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_421
timestamp 1636968456
transform 1 0 39836 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_433
timestamp 1636968456
transform 1 0 40940 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_445
timestamp 1636968456
transform 1 0 42044 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_457
timestamp 1636968456
transform 1 0 43148 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_469
timestamp 1
transform 1 0 44252 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_475
timestamp 1
transform 1 0 44804 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_477
timestamp 1636968456
transform 1 0 44988 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_489
timestamp 1636968456
transform 1 0 46092 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_501
timestamp 1636968456
transform 1 0 47196 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_513
timestamp 1636968456
transform 1 0 48300 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_525
timestamp 1
transform 1 0 49404 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_531
timestamp 1
transform 1 0 49956 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_533
timestamp 1636968456
transform 1 0 50140 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_545
timestamp 1636968456
transform 1 0 51244 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_557
timestamp 1636968456
transform 1 0 52348 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_569
timestamp 1636968456
transform 1 0 53452 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_581
timestamp 1
transform 1 0 54556 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_587
timestamp 1
transform 1 0 55108 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_589
timestamp 1636968456
transform 1 0 55292 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_601
timestamp 1636968456
transform 1 0 56396 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_613
timestamp 1636968456
transform 1 0 57500 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_625
timestamp 1636968456
transform 1 0 58604 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_637
timestamp 1
transform 1 0 59708 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_643
timestamp 1
transform 1 0 60260 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_645
timestamp 1636968456
transform 1 0 60444 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_657
timestamp 1636968456
transform 1 0 61548 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_669
timestamp 1636968456
transform 1 0 62652 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_681
timestamp 1636968456
transform 1 0 63756 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_693
timestamp 1
transform 1 0 64860 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_699
timestamp 1
transform 1 0 65412 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_701
timestamp 1636968456
transform 1 0 65596 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_713
timestamp 1636968456
transform 1 0 66700 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_725
timestamp 1636968456
transform 1 0 67804 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_737
timestamp 1636968456
transform 1 0 68908 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_749
timestamp 1
transform 1 0 70012 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_755
timestamp 1
transform 1 0 70564 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_757
timestamp 1636968456
transform 1 0 70748 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_769
timestamp 1636968456
transform 1 0 71852 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_781
timestamp 1636968456
transform 1 0 72956 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_793
timestamp 1636968456
transform 1 0 74060 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_805
timestamp 1
transform 1 0 75164 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_811
timestamp 1
transform 1 0 75716 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_813
timestamp 1636968456
transform 1 0 75900 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_825
timestamp 1636968456
transform 1 0 77004 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_837
timestamp 1636968456
transform 1 0 78108 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_849
timestamp 1636968456
transform 1 0 79212 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_861
timestamp 1
transform 1 0 80316 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_867
timestamp 1
transform 1 0 80868 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_869
timestamp 1636968456
transform 1 0 81052 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_881
timestamp 1636968456
transform 1 0 82156 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_893
timestamp 1636968456
transform 1 0 83260 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_905
timestamp 1636968456
transform 1 0 84364 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_917
timestamp 1
transform 1 0 85468 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_923
timestamp 1
transform 1 0 86020 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_925
timestamp 1636968456
transform 1 0 86204 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_937
timestamp 1636968456
transform 1 0 87308 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_949
timestamp 1636968456
transform 1 0 88412 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_961
timestamp 1636968456
transform 1 0 89516 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_973
timestamp 1
transform 1 0 90620 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_979
timestamp 1
transform 1 0 91172 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_981
timestamp 1636968456
transform 1 0 91356 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_993
timestamp 1636968456
transform 1 0 92460 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1005
timestamp 1636968456
transform 1 0 93564 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1017
timestamp 1636968456
transform 1 0 94668 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_1029
timestamp 1
transform 1 0 95772 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_1035
timestamp 1
transform 1 0 96324 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1037
timestamp 1636968456
transform 1 0 96508 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1049
timestamp 1636968456
transform 1 0 97612 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1061
timestamp 1636968456
transform 1 0 98716 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1073
timestamp 1636968456
transform 1 0 99820 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_1085
timestamp 1
transform 1 0 100924 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_1091
timestamp 1
transform 1 0 101476 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1093
timestamp 1636968456
transform 1 0 101660 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1105
timestamp 1636968456
transform 1 0 102764 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1117
timestamp 1636968456
transform 1 0 103868 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1129
timestamp 1636968456
transform 1 0 104972 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_1141
timestamp 1
transform 1 0 106076 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_1147
timestamp 1
transform 1 0 106628 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1149
timestamp 1636968456
transform 1 0 106812 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_1161
timestamp 1
transform 1 0 107916 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_1167
timestamp 1
transform 1 0 108468 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_3
timestamp 1636968456
transform 1 0 1380 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_15
timestamp 1636968456
transform 1 0 2484 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_27
timestamp 1636968456
transform 1 0 3588 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_39
timestamp 1636968456
transform 1 0 4692 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_253_51
timestamp 1
transform 1 0 5796 0 -1 140352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_253_55
timestamp 1
transform 1 0 6164 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_57
timestamp 1636968456
transform 1 0 6348 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_69
timestamp 1636968456
transform 1 0 7452 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_81
timestamp 1636968456
transform 1 0 8556 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_93
timestamp 1636968456
transform 1 0 9660 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_105
timestamp 1
transform 1 0 10764 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_111
timestamp 1
transform 1 0 11316 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_113
timestamp 1636968456
transform 1 0 11500 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_125
timestamp 1636968456
transform 1 0 12604 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_137
timestamp 1636968456
transform 1 0 13708 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_149
timestamp 1636968456
transform 1 0 14812 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_161
timestamp 1
transform 1 0 15916 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_167
timestamp 1
transform 1 0 16468 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_169
timestamp 1636968456
transform 1 0 16652 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_181
timestamp 1636968456
transform 1 0 17756 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_193
timestamp 1636968456
transform 1 0 18860 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_205
timestamp 1636968456
transform 1 0 19964 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_217
timestamp 1
transform 1 0 21068 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_223
timestamp 1
transform 1 0 21620 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_225
timestamp 1636968456
transform 1 0 21804 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_237
timestamp 1636968456
transform 1 0 22908 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_249
timestamp 1636968456
transform 1 0 24012 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_261
timestamp 1636968456
transform 1 0 25116 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_273
timestamp 1
transform 1 0 26220 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_279
timestamp 1
transform 1 0 26772 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_281
timestamp 1636968456
transform 1 0 26956 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_293
timestamp 1636968456
transform 1 0 28060 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_305
timestamp 1636968456
transform 1 0 29164 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_317
timestamp 1636968456
transform 1 0 30268 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_329
timestamp 1
transform 1 0 31372 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_335
timestamp 1
transform 1 0 31924 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_337
timestamp 1636968456
transform 1 0 32108 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_349
timestamp 1636968456
transform 1 0 33212 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_361
timestamp 1636968456
transform 1 0 34316 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_373
timestamp 1636968456
transform 1 0 35420 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_385
timestamp 1
transform 1 0 36524 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_391
timestamp 1
transform 1 0 37076 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_393
timestamp 1636968456
transform 1 0 37260 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_405
timestamp 1636968456
transform 1 0 38364 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_417
timestamp 1636968456
transform 1 0 39468 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_429
timestamp 1636968456
transform 1 0 40572 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_441
timestamp 1
transform 1 0 41676 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_447
timestamp 1
transform 1 0 42228 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_449
timestamp 1636968456
transform 1 0 42412 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_461
timestamp 1636968456
transform 1 0 43516 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_473
timestamp 1636968456
transform 1 0 44620 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_485
timestamp 1636968456
transform 1 0 45724 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_497
timestamp 1
transform 1 0 46828 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_503
timestamp 1
transform 1 0 47380 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_505
timestamp 1636968456
transform 1 0 47564 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_517
timestamp 1636968456
transform 1 0 48668 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_529
timestamp 1636968456
transform 1 0 49772 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_541
timestamp 1636968456
transform 1 0 50876 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_553
timestamp 1
transform 1 0 51980 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_559
timestamp 1
transform 1 0 52532 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_561
timestamp 1636968456
transform 1 0 52716 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_573
timestamp 1636968456
transform 1 0 53820 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_585
timestamp 1636968456
transform 1 0 54924 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_597
timestamp 1636968456
transform 1 0 56028 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_609
timestamp 1
transform 1 0 57132 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_615
timestamp 1
transform 1 0 57684 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_617
timestamp 1636968456
transform 1 0 57868 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_629
timestamp 1636968456
transform 1 0 58972 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_641
timestamp 1636968456
transform 1 0 60076 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_653
timestamp 1636968456
transform 1 0 61180 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_665
timestamp 1
transform 1 0 62284 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_671
timestamp 1
transform 1 0 62836 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_673
timestamp 1636968456
transform 1 0 63020 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_685
timestamp 1636968456
transform 1 0 64124 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_697
timestamp 1636968456
transform 1 0 65228 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_709
timestamp 1636968456
transform 1 0 66332 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_721
timestamp 1
transform 1 0 67436 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_727
timestamp 1
transform 1 0 67988 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_729
timestamp 1636968456
transform 1 0 68172 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_741
timestamp 1636968456
transform 1 0 69276 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_753
timestamp 1636968456
transform 1 0 70380 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_765
timestamp 1636968456
transform 1 0 71484 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_777
timestamp 1
transform 1 0 72588 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_783
timestamp 1
transform 1 0 73140 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_785
timestamp 1636968456
transform 1 0 73324 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_797
timestamp 1636968456
transform 1 0 74428 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_809
timestamp 1636968456
transform 1 0 75532 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_821
timestamp 1636968456
transform 1 0 76636 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_833
timestamp 1
transform 1 0 77740 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_839
timestamp 1
transform 1 0 78292 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_841
timestamp 1636968456
transform 1 0 78476 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_853
timestamp 1636968456
transform 1 0 79580 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_865
timestamp 1636968456
transform 1 0 80684 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_877
timestamp 1636968456
transform 1 0 81788 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_889
timestamp 1
transform 1 0 82892 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_895
timestamp 1
transform 1 0 83444 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_897
timestamp 1636968456
transform 1 0 83628 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_909
timestamp 1636968456
transform 1 0 84732 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_921
timestamp 1636968456
transform 1 0 85836 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_933
timestamp 1636968456
transform 1 0 86940 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_945
timestamp 1
transform 1 0 88044 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_951
timestamp 1
transform 1 0 88596 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_953
timestamp 1636968456
transform 1 0 88780 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_965
timestamp 1636968456
transform 1 0 89884 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_977
timestamp 1636968456
transform 1 0 90988 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_989
timestamp 1636968456
transform 1 0 92092 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_1001
timestamp 1
transform 1 0 93196 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_1007
timestamp 1
transform 1 0 93748 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1009
timestamp 1636968456
transform 1 0 93932 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1021
timestamp 1636968456
transform 1 0 95036 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1033
timestamp 1636968456
transform 1 0 96140 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1045
timestamp 1636968456
transform 1 0 97244 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_1057
timestamp 1
transform 1 0 98348 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_1063
timestamp 1
transform 1 0 98900 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1065
timestamp 1636968456
transform 1 0 99084 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1077
timestamp 1636968456
transform 1 0 100188 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1089
timestamp 1636968456
transform 1 0 101292 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1101
timestamp 1636968456
transform 1 0 102396 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_1113
timestamp 1
transform 1 0 103500 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_1119
timestamp 1
transform 1 0 104052 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1121
timestamp 1636968456
transform 1 0 104236 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1133
timestamp 1636968456
transform 1 0 105340 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1145
timestamp 1636968456
transform 1 0 106444 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_253_1157
timestamp 1
transform 1 0 107548 0 -1 140352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_253_1165
timestamp 1
transform 1 0 108284 0 -1 140352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_254_3
timestamp 1636968456
transform 1 0 1380 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_15
timestamp 1636968456
transform 1 0 2484 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_254_27
timestamp 1
transform 1 0 3588 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_29
timestamp 1636968456
transform 1 0 3772 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_41
timestamp 1636968456
transform 1 0 4876 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_53
timestamp 1636968456
transform 1 0 5980 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_65
timestamp 1636968456
transform 1 0 7084 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_77
timestamp 1
transform 1 0 8188 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_83
timestamp 1
transform 1 0 8740 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_85
timestamp 1636968456
transform 1 0 8924 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_97
timestamp 1636968456
transform 1 0 10028 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_109
timestamp 1636968456
transform 1 0 11132 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_121
timestamp 1636968456
transform 1 0 12236 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_133
timestamp 1
transform 1 0 13340 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_139
timestamp 1
transform 1 0 13892 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_141
timestamp 1636968456
transform 1 0 14076 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_153
timestamp 1636968456
transform 1 0 15180 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_165
timestamp 1636968456
transform 1 0 16284 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_177
timestamp 1636968456
transform 1 0 17388 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_189
timestamp 1
transform 1 0 18492 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_195
timestamp 1
transform 1 0 19044 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_197
timestamp 1636968456
transform 1 0 19228 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_209
timestamp 1636968456
transform 1 0 20332 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_221
timestamp 1636968456
transform 1 0 21436 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_233
timestamp 1636968456
transform 1 0 22540 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_245
timestamp 1
transform 1 0 23644 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_251
timestamp 1
transform 1 0 24196 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_253
timestamp 1636968456
transform 1 0 24380 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_265
timestamp 1636968456
transform 1 0 25484 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_277
timestamp 1636968456
transform 1 0 26588 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_289
timestamp 1636968456
transform 1 0 27692 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_301
timestamp 1
transform 1 0 28796 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_307
timestamp 1
transform 1 0 29348 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_309
timestamp 1636968456
transform 1 0 29532 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_321
timestamp 1636968456
transform 1 0 30636 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_333
timestamp 1636968456
transform 1 0 31740 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_345
timestamp 1636968456
transform 1 0 32844 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_357
timestamp 1
transform 1 0 33948 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_363
timestamp 1
transform 1 0 34500 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_365
timestamp 1636968456
transform 1 0 34684 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_377
timestamp 1636968456
transform 1 0 35788 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_389
timestamp 1636968456
transform 1 0 36892 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_401
timestamp 1636968456
transform 1 0 37996 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_413
timestamp 1
transform 1 0 39100 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_419
timestamp 1
transform 1 0 39652 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_421
timestamp 1636968456
transform 1 0 39836 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_433
timestamp 1636968456
transform 1 0 40940 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_445
timestamp 1636968456
transform 1 0 42044 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_457
timestamp 1636968456
transform 1 0 43148 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_469
timestamp 1
transform 1 0 44252 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_475
timestamp 1
transform 1 0 44804 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_477
timestamp 1636968456
transform 1 0 44988 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_489
timestamp 1636968456
transform 1 0 46092 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_501
timestamp 1636968456
transform 1 0 47196 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_513
timestamp 1636968456
transform 1 0 48300 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_525
timestamp 1
transform 1 0 49404 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_531
timestamp 1
transform 1 0 49956 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_533
timestamp 1636968456
transform 1 0 50140 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_545
timestamp 1636968456
transform 1 0 51244 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_557
timestamp 1636968456
transform 1 0 52348 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_569
timestamp 1636968456
transform 1 0 53452 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_581
timestamp 1
transform 1 0 54556 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_587
timestamp 1
transform 1 0 55108 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_589
timestamp 1636968456
transform 1 0 55292 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_601
timestamp 1636968456
transform 1 0 56396 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_613
timestamp 1636968456
transform 1 0 57500 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_625
timestamp 1636968456
transform 1 0 58604 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_637
timestamp 1
transform 1 0 59708 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_643
timestamp 1
transform 1 0 60260 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_645
timestamp 1636968456
transform 1 0 60444 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_657
timestamp 1636968456
transform 1 0 61548 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_669
timestamp 1636968456
transform 1 0 62652 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_681
timestamp 1636968456
transform 1 0 63756 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_693
timestamp 1
transform 1 0 64860 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_699
timestamp 1
transform 1 0 65412 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_701
timestamp 1636968456
transform 1 0 65596 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_713
timestamp 1636968456
transform 1 0 66700 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_725
timestamp 1636968456
transform 1 0 67804 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_737
timestamp 1636968456
transform 1 0 68908 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_749
timestamp 1
transform 1 0 70012 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_755
timestamp 1
transform 1 0 70564 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_757
timestamp 1636968456
transform 1 0 70748 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_769
timestamp 1636968456
transform 1 0 71852 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_781
timestamp 1636968456
transform 1 0 72956 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_793
timestamp 1636968456
transform 1 0 74060 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_805
timestamp 1
transform 1 0 75164 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_811
timestamp 1
transform 1 0 75716 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_813
timestamp 1636968456
transform 1 0 75900 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_825
timestamp 1636968456
transform 1 0 77004 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_837
timestamp 1636968456
transform 1 0 78108 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_849
timestamp 1636968456
transform 1 0 79212 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_861
timestamp 1
transform 1 0 80316 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_867
timestamp 1
transform 1 0 80868 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_869
timestamp 1636968456
transform 1 0 81052 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_881
timestamp 1636968456
transform 1 0 82156 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_893
timestamp 1636968456
transform 1 0 83260 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_905
timestamp 1636968456
transform 1 0 84364 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_917
timestamp 1
transform 1 0 85468 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_923
timestamp 1
transform 1 0 86020 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_925
timestamp 1636968456
transform 1 0 86204 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_937
timestamp 1636968456
transform 1 0 87308 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_949
timestamp 1636968456
transform 1 0 88412 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_961
timestamp 1636968456
transform 1 0 89516 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_973
timestamp 1
transform 1 0 90620 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_979
timestamp 1
transform 1 0 91172 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_981
timestamp 1636968456
transform 1 0 91356 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_993
timestamp 1636968456
transform 1 0 92460 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1005
timestamp 1636968456
transform 1 0 93564 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1017
timestamp 1636968456
transform 1 0 94668 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_1029
timestamp 1
transform 1 0 95772 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_1035
timestamp 1
transform 1 0 96324 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1037
timestamp 1636968456
transform 1 0 96508 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1049
timestamp 1636968456
transform 1 0 97612 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1061
timestamp 1636968456
transform 1 0 98716 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1073
timestamp 1636968456
transform 1 0 99820 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_1085
timestamp 1
transform 1 0 100924 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_1091
timestamp 1
transform 1 0 101476 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1093
timestamp 1636968456
transform 1 0 101660 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1105
timestamp 1636968456
transform 1 0 102764 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1117
timestamp 1636968456
transform 1 0 103868 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1129
timestamp 1636968456
transform 1 0 104972 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_1141
timestamp 1
transform 1 0 106076 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_1147
timestamp 1
transform 1 0 106628 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1149
timestamp 1636968456
transform 1 0 106812 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_1161
timestamp 1
transform 1 0 107916 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_1167
timestamp 1
transform 1 0 108468 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_3
timestamp 1636968456
transform 1 0 1380 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_15
timestamp 1636968456
transform 1 0 2484 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_27
timestamp 1636968456
transform 1 0 3588 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_39
timestamp 1636968456
transform 1 0 4692 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_255_51
timestamp 1
transform 1 0 5796 0 -1 141440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_255_55
timestamp 1
transform 1 0 6164 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_57
timestamp 1636968456
transform 1 0 6348 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_69
timestamp 1636968456
transform 1 0 7452 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_81
timestamp 1636968456
transform 1 0 8556 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_93
timestamp 1636968456
transform 1 0 9660 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_105
timestamp 1
transform 1 0 10764 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_111
timestamp 1
transform 1 0 11316 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_113
timestamp 1636968456
transform 1 0 11500 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_125
timestamp 1636968456
transform 1 0 12604 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_137
timestamp 1636968456
transform 1 0 13708 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_149
timestamp 1636968456
transform 1 0 14812 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_161
timestamp 1
transform 1 0 15916 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_167
timestamp 1
transform 1 0 16468 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_169
timestamp 1636968456
transform 1 0 16652 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_181
timestamp 1636968456
transform 1 0 17756 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_193
timestamp 1636968456
transform 1 0 18860 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_205
timestamp 1636968456
transform 1 0 19964 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_217
timestamp 1
transform 1 0 21068 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_223
timestamp 1
transform 1 0 21620 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_225
timestamp 1636968456
transform 1 0 21804 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_237
timestamp 1636968456
transform 1 0 22908 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_249
timestamp 1636968456
transform 1 0 24012 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_261
timestamp 1636968456
transform 1 0 25116 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_273
timestamp 1
transform 1 0 26220 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_279
timestamp 1
transform 1 0 26772 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_281
timestamp 1636968456
transform 1 0 26956 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_293
timestamp 1636968456
transform 1 0 28060 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_305
timestamp 1636968456
transform 1 0 29164 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_317
timestamp 1636968456
transform 1 0 30268 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_329
timestamp 1
transform 1 0 31372 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_335
timestamp 1
transform 1 0 31924 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_337
timestamp 1636968456
transform 1 0 32108 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_349
timestamp 1636968456
transform 1 0 33212 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_361
timestamp 1636968456
transform 1 0 34316 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_373
timestamp 1636968456
transform 1 0 35420 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_385
timestamp 1
transform 1 0 36524 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_391
timestamp 1
transform 1 0 37076 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_393
timestamp 1636968456
transform 1 0 37260 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_405
timestamp 1636968456
transform 1 0 38364 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_417
timestamp 1636968456
transform 1 0 39468 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_429
timestamp 1636968456
transform 1 0 40572 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_441
timestamp 1
transform 1 0 41676 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_447
timestamp 1
transform 1 0 42228 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_449
timestamp 1636968456
transform 1 0 42412 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_461
timestamp 1636968456
transform 1 0 43516 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_473
timestamp 1636968456
transform 1 0 44620 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_485
timestamp 1636968456
transform 1 0 45724 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_497
timestamp 1
transform 1 0 46828 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_503
timestamp 1
transform 1 0 47380 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_505
timestamp 1636968456
transform 1 0 47564 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_517
timestamp 1636968456
transform 1 0 48668 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_529
timestamp 1636968456
transform 1 0 49772 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_541
timestamp 1636968456
transform 1 0 50876 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_553
timestamp 1
transform 1 0 51980 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_559
timestamp 1
transform 1 0 52532 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_561
timestamp 1636968456
transform 1 0 52716 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_573
timestamp 1636968456
transform 1 0 53820 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_585
timestamp 1636968456
transform 1 0 54924 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_597
timestamp 1636968456
transform 1 0 56028 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_609
timestamp 1
transform 1 0 57132 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_615
timestamp 1
transform 1 0 57684 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_617
timestamp 1636968456
transform 1 0 57868 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_629
timestamp 1636968456
transform 1 0 58972 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_641
timestamp 1636968456
transform 1 0 60076 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_653
timestamp 1636968456
transform 1 0 61180 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_665
timestamp 1
transform 1 0 62284 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_671
timestamp 1
transform 1 0 62836 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_673
timestamp 1636968456
transform 1 0 63020 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_685
timestamp 1636968456
transform 1 0 64124 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_697
timestamp 1636968456
transform 1 0 65228 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_709
timestamp 1636968456
transform 1 0 66332 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_721
timestamp 1
transform 1 0 67436 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_727
timestamp 1
transform 1 0 67988 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_729
timestamp 1636968456
transform 1 0 68172 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_741
timestamp 1636968456
transform 1 0 69276 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_753
timestamp 1636968456
transform 1 0 70380 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_765
timestamp 1636968456
transform 1 0 71484 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_777
timestamp 1
transform 1 0 72588 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_783
timestamp 1
transform 1 0 73140 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_785
timestamp 1636968456
transform 1 0 73324 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_797
timestamp 1636968456
transform 1 0 74428 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_809
timestamp 1636968456
transform 1 0 75532 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_821
timestamp 1636968456
transform 1 0 76636 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_833
timestamp 1
transform 1 0 77740 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_839
timestamp 1
transform 1 0 78292 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_841
timestamp 1636968456
transform 1 0 78476 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_853
timestamp 1636968456
transform 1 0 79580 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_865
timestamp 1636968456
transform 1 0 80684 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_877
timestamp 1636968456
transform 1 0 81788 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_889
timestamp 1
transform 1 0 82892 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_895
timestamp 1
transform 1 0 83444 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_897
timestamp 1636968456
transform 1 0 83628 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_909
timestamp 1636968456
transform 1 0 84732 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_921
timestamp 1636968456
transform 1 0 85836 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_933
timestamp 1636968456
transform 1 0 86940 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_945
timestamp 1
transform 1 0 88044 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_951
timestamp 1
transform 1 0 88596 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_953
timestamp 1636968456
transform 1 0 88780 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_965
timestamp 1636968456
transform 1 0 89884 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_977
timestamp 1636968456
transform 1 0 90988 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_989
timestamp 1636968456
transform 1 0 92092 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_1001
timestamp 1
transform 1 0 93196 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_1007
timestamp 1
transform 1 0 93748 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1009
timestamp 1636968456
transform 1 0 93932 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1021
timestamp 1636968456
transform 1 0 95036 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1033
timestamp 1636968456
transform 1 0 96140 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1045
timestamp 1636968456
transform 1 0 97244 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_1057
timestamp 1
transform 1 0 98348 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_1063
timestamp 1
transform 1 0 98900 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1065
timestamp 1636968456
transform 1 0 99084 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1077
timestamp 1636968456
transform 1 0 100188 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1089
timestamp 1636968456
transform 1 0 101292 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1101
timestamp 1636968456
transform 1 0 102396 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_1113
timestamp 1
transform 1 0 103500 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_1119
timestamp 1
transform 1 0 104052 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1121
timestamp 1636968456
transform 1 0 104236 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1133
timestamp 1636968456
transform 1 0 105340 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1145
timestamp 1636968456
transform 1 0 106444 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_255_1157
timestamp 1
transform 1 0 107548 0 -1 141440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_255_1165
timestamp 1
transform 1 0 108284 0 -1 141440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_256_3
timestamp 1636968456
transform 1 0 1380 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_15
timestamp 1636968456
transform 1 0 2484 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_256_27
timestamp 1
transform 1 0 3588 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_29
timestamp 1636968456
transform 1 0 3772 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_41
timestamp 1636968456
transform 1 0 4876 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_53
timestamp 1636968456
transform 1 0 5980 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_65
timestamp 1636968456
transform 1 0 7084 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_77
timestamp 1
transform 1 0 8188 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_83
timestamp 1
transform 1 0 8740 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_85
timestamp 1636968456
transform 1 0 8924 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_97
timestamp 1636968456
transform 1 0 10028 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_109
timestamp 1636968456
transform 1 0 11132 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_121
timestamp 1636968456
transform 1 0 12236 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_133
timestamp 1
transform 1 0 13340 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_139
timestamp 1
transform 1 0 13892 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_141
timestamp 1636968456
transform 1 0 14076 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_153
timestamp 1636968456
transform 1 0 15180 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_165
timestamp 1636968456
transform 1 0 16284 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_177
timestamp 1636968456
transform 1 0 17388 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_189
timestamp 1
transform 1 0 18492 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_195
timestamp 1
transform 1 0 19044 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_197
timestamp 1636968456
transform 1 0 19228 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_209
timestamp 1636968456
transform 1 0 20332 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_221
timestamp 1636968456
transform 1 0 21436 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_233
timestamp 1636968456
transform 1 0 22540 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_245
timestamp 1
transform 1 0 23644 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_251
timestamp 1
transform 1 0 24196 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_253
timestamp 1636968456
transform 1 0 24380 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_265
timestamp 1636968456
transform 1 0 25484 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_277
timestamp 1636968456
transform 1 0 26588 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_289
timestamp 1636968456
transform 1 0 27692 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_301
timestamp 1
transform 1 0 28796 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_307
timestamp 1
transform 1 0 29348 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_309
timestamp 1636968456
transform 1 0 29532 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_321
timestamp 1636968456
transform 1 0 30636 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_333
timestamp 1636968456
transform 1 0 31740 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_345
timestamp 1636968456
transform 1 0 32844 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_357
timestamp 1
transform 1 0 33948 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_363
timestamp 1
transform 1 0 34500 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_365
timestamp 1636968456
transform 1 0 34684 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_377
timestamp 1636968456
transform 1 0 35788 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_389
timestamp 1636968456
transform 1 0 36892 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_401
timestamp 1636968456
transform 1 0 37996 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_413
timestamp 1
transform 1 0 39100 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_419
timestamp 1
transform 1 0 39652 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_421
timestamp 1636968456
transform 1 0 39836 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_433
timestamp 1636968456
transform 1 0 40940 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_445
timestamp 1636968456
transform 1 0 42044 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_457
timestamp 1636968456
transform 1 0 43148 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_469
timestamp 1
transform 1 0 44252 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_475
timestamp 1
transform 1 0 44804 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_477
timestamp 1636968456
transform 1 0 44988 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_489
timestamp 1636968456
transform 1 0 46092 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_501
timestamp 1636968456
transform 1 0 47196 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_513
timestamp 1636968456
transform 1 0 48300 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_525
timestamp 1
transform 1 0 49404 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_531
timestamp 1
transform 1 0 49956 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_533
timestamp 1636968456
transform 1 0 50140 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_545
timestamp 1636968456
transform 1 0 51244 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_557
timestamp 1636968456
transform 1 0 52348 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_569
timestamp 1636968456
transform 1 0 53452 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_581
timestamp 1
transform 1 0 54556 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_587
timestamp 1
transform 1 0 55108 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_589
timestamp 1636968456
transform 1 0 55292 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_601
timestamp 1636968456
transform 1 0 56396 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_613
timestamp 1636968456
transform 1 0 57500 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_625
timestamp 1636968456
transform 1 0 58604 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_637
timestamp 1
transform 1 0 59708 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_643
timestamp 1
transform 1 0 60260 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_645
timestamp 1636968456
transform 1 0 60444 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_657
timestamp 1636968456
transform 1 0 61548 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_669
timestamp 1636968456
transform 1 0 62652 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_681
timestamp 1636968456
transform 1 0 63756 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_693
timestamp 1
transform 1 0 64860 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_699
timestamp 1
transform 1 0 65412 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_701
timestamp 1636968456
transform 1 0 65596 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_713
timestamp 1636968456
transform 1 0 66700 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_725
timestamp 1636968456
transform 1 0 67804 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_737
timestamp 1636968456
transform 1 0 68908 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_749
timestamp 1
transform 1 0 70012 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_755
timestamp 1
transform 1 0 70564 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_757
timestamp 1636968456
transform 1 0 70748 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_769
timestamp 1636968456
transform 1 0 71852 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_781
timestamp 1636968456
transform 1 0 72956 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_793
timestamp 1636968456
transform 1 0 74060 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_805
timestamp 1
transform 1 0 75164 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_811
timestamp 1
transform 1 0 75716 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_813
timestamp 1636968456
transform 1 0 75900 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_825
timestamp 1636968456
transform 1 0 77004 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_837
timestamp 1636968456
transform 1 0 78108 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_849
timestamp 1636968456
transform 1 0 79212 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_861
timestamp 1
transform 1 0 80316 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_867
timestamp 1
transform 1 0 80868 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_869
timestamp 1636968456
transform 1 0 81052 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_881
timestamp 1636968456
transform 1 0 82156 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_893
timestamp 1636968456
transform 1 0 83260 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_905
timestamp 1636968456
transform 1 0 84364 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_917
timestamp 1
transform 1 0 85468 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_923
timestamp 1
transform 1 0 86020 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_925
timestamp 1636968456
transform 1 0 86204 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_937
timestamp 1636968456
transform 1 0 87308 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_949
timestamp 1636968456
transform 1 0 88412 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_961
timestamp 1636968456
transform 1 0 89516 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_973
timestamp 1
transform 1 0 90620 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_979
timestamp 1
transform 1 0 91172 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_981
timestamp 1636968456
transform 1 0 91356 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_993
timestamp 1636968456
transform 1 0 92460 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1005
timestamp 1636968456
transform 1 0 93564 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1017
timestamp 1636968456
transform 1 0 94668 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_1029
timestamp 1
transform 1 0 95772 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_1035
timestamp 1
transform 1 0 96324 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1037
timestamp 1636968456
transform 1 0 96508 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1049
timestamp 1636968456
transform 1 0 97612 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1061
timestamp 1636968456
transform 1 0 98716 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1073
timestamp 1636968456
transform 1 0 99820 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_1085
timestamp 1
transform 1 0 100924 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_1091
timestamp 1
transform 1 0 101476 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1093
timestamp 1636968456
transform 1 0 101660 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1105
timestamp 1636968456
transform 1 0 102764 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1117
timestamp 1636968456
transform 1 0 103868 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1129
timestamp 1636968456
transform 1 0 104972 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_1141
timestamp 1
transform 1 0 106076 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_1147
timestamp 1
transform 1 0 106628 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1149
timestamp 1636968456
transform 1 0 106812 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_1161
timestamp 1
transform 1 0 107916 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_1167
timestamp 1
transform 1 0 108468 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_3
timestamp 1636968456
transform 1 0 1380 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_15
timestamp 1636968456
transform 1 0 2484 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_27
timestamp 1636968456
transform 1 0 3588 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_39
timestamp 1636968456
transform 1 0 4692 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_257_51
timestamp 1
transform 1 0 5796 0 -1 142528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_257_55
timestamp 1
transform 1 0 6164 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_57
timestamp 1636968456
transform 1 0 6348 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_69
timestamp 1636968456
transform 1 0 7452 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_81
timestamp 1636968456
transform 1 0 8556 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_93
timestamp 1636968456
transform 1 0 9660 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_105
timestamp 1
transform 1 0 10764 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_111
timestamp 1
transform 1 0 11316 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_113
timestamp 1636968456
transform 1 0 11500 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_125
timestamp 1636968456
transform 1 0 12604 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_137
timestamp 1636968456
transform 1 0 13708 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_149
timestamp 1636968456
transform 1 0 14812 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_161
timestamp 1
transform 1 0 15916 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_167
timestamp 1
transform 1 0 16468 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_169
timestamp 1636968456
transform 1 0 16652 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_181
timestamp 1636968456
transform 1 0 17756 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_193
timestamp 1636968456
transform 1 0 18860 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_205
timestamp 1636968456
transform 1 0 19964 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_217
timestamp 1
transform 1 0 21068 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_223
timestamp 1
transform 1 0 21620 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_225
timestamp 1636968456
transform 1 0 21804 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_237
timestamp 1636968456
transform 1 0 22908 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_249
timestamp 1636968456
transform 1 0 24012 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_261
timestamp 1636968456
transform 1 0 25116 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_273
timestamp 1
transform 1 0 26220 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_279
timestamp 1
transform 1 0 26772 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_281
timestamp 1636968456
transform 1 0 26956 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_293
timestamp 1636968456
transform 1 0 28060 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_305
timestamp 1636968456
transform 1 0 29164 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_317
timestamp 1636968456
transform 1 0 30268 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_329
timestamp 1
transform 1 0 31372 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_335
timestamp 1
transform 1 0 31924 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_337
timestamp 1636968456
transform 1 0 32108 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_349
timestamp 1636968456
transform 1 0 33212 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_361
timestamp 1636968456
transform 1 0 34316 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_373
timestamp 1636968456
transform 1 0 35420 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_385
timestamp 1
transform 1 0 36524 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_391
timestamp 1
transform 1 0 37076 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_393
timestamp 1636968456
transform 1 0 37260 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_405
timestamp 1636968456
transform 1 0 38364 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_417
timestamp 1636968456
transform 1 0 39468 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_429
timestamp 1636968456
transform 1 0 40572 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_441
timestamp 1
transform 1 0 41676 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_447
timestamp 1
transform 1 0 42228 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_449
timestamp 1636968456
transform 1 0 42412 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_461
timestamp 1636968456
transform 1 0 43516 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_473
timestamp 1636968456
transform 1 0 44620 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_485
timestamp 1636968456
transform 1 0 45724 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_497
timestamp 1
transform 1 0 46828 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_503
timestamp 1
transform 1 0 47380 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_505
timestamp 1636968456
transform 1 0 47564 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_517
timestamp 1636968456
transform 1 0 48668 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_529
timestamp 1636968456
transform 1 0 49772 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_541
timestamp 1636968456
transform 1 0 50876 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_553
timestamp 1
transform 1 0 51980 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_559
timestamp 1
transform 1 0 52532 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_561
timestamp 1636968456
transform 1 0 52716 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_573
timestamp 1636968456
transform 1 0 53820 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_585
timestamp 1636968456
transform 1 0 54924 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_597
timestamp 1636968456
transform 1 0 56028 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_609
timestamp 1
transform 1 0 57132 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_615
timestamp 1
transform 1 0 57684 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_617
timestamp 1636968456
transform 1 0 57868 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_629
timestamp 1636968456
transform 1 0 58972 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_641
timestamp 1636968456
transform 1 0 60076 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_653
timestamp 1636968456
transform 1 0 61180 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_665
timestamp 1
transform 1 0 62284 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_671
timestamp 1
transform 1 0 62836 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_673
timestamp 1636968456
transform 1 0 63020 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_685
timestamp 1636968456
transform 1 0 64124 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_697
timestamp 1636968456
transform 1 0 65228 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_709
timestamp 1636968456
transform 1 0 66332 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_721
timestamp 1
transform 1 0 67436 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_727
timestamp 1
transform 1 0 67988 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_729
timestamp 1636968456
transform 1 0 68172 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_741
timestamp 1636968456
transform 1 0 69276 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_753
timestamp 1636968456
transform 1 0 70380 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_765
timestamp 1636968456
transform 1 0 71484 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_777
timestamp 1
transform 1 0 72588 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_783
timestamp 1
transform 1 0 73140 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_785
timestamp 1636968456
transform 1 0 73324 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_797
timestamp 1636968456
transform 1 0 74428 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_809
timestamp 1636968456
transform 1 0 75532 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_821
timestamp 1636968456
transform 1 0 76636 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_833
timestamp 1
transform 1 0 77740 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_839
timestamp 1
transform 1 0 78292 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_841
timestamp 1636968456
transform 1 0 78476 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_853
timestamp 1636968456
transform 1 0 79580 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_865
timestamp 1636968456
transform 1 0 80684 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_877
timestamp 1636968456
transform 1 0 81788 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_889
timestamp 1
transform 1 0 82892 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_895
timestamp 1
transform 1 0 83444 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_897
timestamp 1636968456
transform 1 0 83628 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_909
timestamp 1636968456
transform 1 0 84732 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_921
timestamp 1636968456
transform 1 0 85836 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_933
timestamp 1636968456
transform 1 0 86940 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_945
timestamp 1
transform 1 0 88044 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_951
timestamp 1
transform 1 0 88596 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_953
timestamp 1636968456
transform 1 0 88780 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_965
timestamp 1636968456
transform 1 0 89884 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_977
timestamp 1636968456
transform 1 0 90988 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_989
timestamp 1636968456
transform 1 0 92092 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_1001
timestamp 1
transform 1 0 93196 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_1007
timestamp 1
transform 1 0 93748 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1009
timestamp 1636968456
transform 1 0 93932 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1021
timestamp 1636968456
transform 1 0 95036 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1033
timestamp 1636968456
transform 1 0 96140 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1045
timestamp 1636968456
transform 1 0 97244 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_1057
timestamp 1
transform 1 0 98348 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_1063
timestamp 1
transform 1 0 98900 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1065
timestamp 1636968456
transform 1 0 99084 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1077
timestamp 1636968456
transform 1 0 100188 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1089
timestamp 1636968456
transform 1 0 101292 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1101
timestamp 1636968456
transform 1 0 102396 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_1113
timestamp 1
transform 1 0 103500 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_1119
timestamp 1
transform 1 0 104052 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1121
timestamp 1636968456
transform 1 0 104236 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1133
timestamp 1636968456
transform 1 0 105340 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1145
timestamp 1636968456
transform 1 0 106444 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_257_1157
timestamp 1
transform 1 0 107548 0 -1 142528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_257_1165
timestamp 1
transform 1 0 108284 0 -1 142528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_258_3
timestamp 1636968456
transform 1 0 1380 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_15
timestamp 1636968456
transform 1 0 2484 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_258_27
timestamp 1
transform 1 0 3588 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_29
timestamp 1636968456
transform 1 0 3772 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_41
timestamp 1636968456
transform 1 0 4876 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_53
timestamp 1636968456
transform 1 0 5980 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_65
timestamp 1636968456
transform 1 0 7084 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_77
timestamp 1
transform 1 0 8188 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_83
timestamp 1
transform 1 0 8740 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_85
timestamp 1636968456
transform 1 0 8924 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_97
timestamp 1636968456
transform 1 0 10028 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_109
timestamp 1636968456
transform 1 0 11132 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_121
timestamp 1636968456
transform 1 0 12236 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_133
timestamp 1
transform 1 0 13340 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_139
timestamp 1
transform 1 0 13892 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_141
timestamp 1636968456
transform 1 0 14076 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_153
timestamp 1636968456
transform 1 0 15180 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_165
timestamp 1636968456
transform 1 0 16284 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_177
timestamp 1636968456
transform 1 0 17388 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_189
timestamp 1
transform 1 0 18492 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_195
timestamp 1
transform 1 0 19044 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_197
timestamp 1636968456
transform 1 0 19228 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_209
timestamp 1636968456
transform 1 0 20332 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_221
timestamp 1636968456
transform 1 0 21436 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_233
timestamp 1636968456
transform 1 0 22540 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_245
timestamp 1
transform 1 0 23644 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_251
timestamp 1
transform 1 0 24196 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_253
timestamp 1636968456
transform 1 0 24380 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_265
timestamp 1636968456
transform 1 0 25484 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_277
timestamp 1636968456
transform 1 0 26588 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_289
timestamp 1636968456
transform 1 0 27692 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_301
timestamp 1
transform 1 0 28796 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_307
timestamp 1
transform 1 0 29348 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_309
timestamp 1636968456
transform 1 0 29532 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_321
timestamp 1636968456
transform 1 0 30636 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_333
timestamp 1636968456
transform 1 0 31740 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_345
timestamp 1636968456
transform 1 0 32844 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_357
timestamp 1
transform 1 0 33948 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_363
timestamp 1
transform 1 0 34500 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_365
timestamp 1636968456
transform 1 0 34684 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_377
timestamp 1636968456
transform 1 0 35788 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_389
timestamp 1636968456
transform 1 0 36892 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_401
timestamp 1636968456
transform 1 0 37996 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_413
timestamp 1
transform 1 0 39100 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_419
timestamp 1
transform 1 0 39652 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_421
timestamp 1636968456
transform 1 0 39836 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_433
timestamp 1636968456
transform 1 0 40940 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_445
timestamp 1636968456
transform 1 0 42044 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_457
timestamp 1636968456
transform 1 0 43148 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_469
timestamp 1
transform 1 0 44252 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_475
timestamp 1
transform 1 0 44804 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_477
timestamp 1636968456
transform 1 0 44988 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_489
timestamp 1636968456
transform 1 0 46092 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_501
timestamp 1636968456
transform 1 0 47196 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_513
timestamp 1636968456
transform 1 0 48300 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_525
timestamp 1
transform 1 0 49404 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_531
timestamp 1
transform 1 0 49956 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_533
timestamp 1636968456
transform 1 0 50140 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_545
timestamp 1636968456
transform 1 0 51244 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_557
timestamp 1636968456
transform 1 0 52348 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_569
timestamp 1636968456
transform 1 0 53452 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_581
timestamp 1
transform 1 0 54556 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_587
timestamp 1
transform 1 0 55108 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_589
timestamp 1636968456
transform 1 0 55292 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_601
timestamp 1636968456
transform 1 0 56396 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_613
timestamp 1636968456
transform 1 0 57500 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_625
timestamp 1636968456
transform 1 0 58604 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_637
timestamp 1
transform 1 0 59708 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_643
timestamp 1
transform 1 0 60260 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_645
timestamp 1636968456
transform 1 0 60444 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_657
timestamp 1636968456
transform 1 0 61548 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_669
timestamp 1636968456
transform 1 0 62652 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_681
timestamp 1636968456
transform 1 0 63756 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_693
timestamp 1
transform 1 0 64860 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_699
timestamp 1
transform 1 0 65412 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_701
timestamp 1636968456
transform 1 0 65596 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_713
timestamp 1636968456
transform 1 0 66700 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_725
timestamp 1636968456
transform 1 0 67804 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_737
timestamp 1636968456
transform 1 0 68908 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_749
timestamp 1
transform 1 0 70012 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_755
timestamp 1
transform 1 0 70564 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_757
timestamp 1636968456
transform 1 0 70748 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_769
timestamp 1636968456
transform 1 0 71852 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_781
timestamp 1636968456
transform 1 0 72956 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_793
timestamp 1636968456
transform 1 0 74060 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_805
timestamp 1
transform 1 0 75164 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_811
timestamp 1
transform 1 0 75716 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_813
timestamp 1636968456
transform 1 0 75900 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_825
timestamp 1636968456
transform 1 0 77004 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_837
timestamp 1636968456
transform 1 0 78108 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_849
timestamp 1636968456
transform 1 0 79212 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_861
timestamp 1
transform 1 0 80316 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_867
timestamp 1
transform 1 0 80868 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_869
timestamp 1636968456
transform 1 0 81052 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_881
timestamp 1636968456
transform 1 0 82156 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_893
timestamp 1636968456
transform 1 0 83260 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_905
timestamp 1636968456
transform 1 0 84364 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_917
timestamp 1
transform 1 0 85468 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_923
timestamp 1
transform 1 0 86020 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_925
timestamp 1636968456
transform 1 0 86204 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_937
timestamp 1636968456
transform 1 0 87308 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_949
timestamp 1636968456
transform 1 0 88412 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_961
timestamp 1636968456
transform 1 0 89516 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_973
timestamp 1
transform 1 0 90620 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_979
timestamp 1
transform 1 0 91172 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_981
timestamp 1636968456
transform 1 0 91356 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_993
timestamp 1636968456
transform 1 0 92460 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1005
timestamp 1636968456
transform 1 0 93564 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1017
timestamp 1636968456
transform 1 0 94668 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_1029
timestamp 1
transform 1 0 95772 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_1035
timestamp 1
transform 1 0 96324 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1037
timestamp 1636968456
transform 1 0 96508 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1049
timestamp 1636968456
transform 1 0 97612 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1061
timestamp 1636968456
transform 1 0 98716 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1073
timestamp 1636968456
transform 1 0 99820 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_1085
timestamp 1
transform 1 0 100924 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_1091
timestamp 1
transform 1 0 101476 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1093
timestamp 1636968456
transform 1 0 101660 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1105
timestamp 1636968456
transform 1 0 102764 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1117
timestamp 1636968456
transform 1 0 103868 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1129
timestamp 1636968456
transform 1 0 104972 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_1141
timestamp 1
transform 1 0 106076 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_1147
timestamp 1
transform 1 0 106628 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1149
timestamp 1636968456
transform 1 0 106812 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_1161
timestamp 1
transform 1 0 107916 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_1167
timestamp 1
transform 1 0 108468 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_3
timestamp 1636968456
transform 1 0 1380 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_15
timestamp 1636968456
transform 1 0 2484 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_27
timestamp 1636968456
transform 1 0 3588 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_39
timestamp 1636968456
transform 1 0 4692 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_259_51
timestamp 1
transform 1 0 5796 0 -1 143616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_259_55
timestamp 1
transform 1 0 6164 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_57
timestamp 1636968456
transform 1 0 6348 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_69
timestamp 1636968456
transform 1 0 7452 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_81
timestamp 1636968456
transform 1 0 8556 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_93
timestamp 1636968456
transform 1 0 9660 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_105
timestamp 1
transform 1 0 10764 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_111
timestamp 1
transform 1 0 11316 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_113
timestamp 1636968456
transform 1 0 11500 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_125
timestamp 1636968456
transform 1 0 12604 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_137
timestamp 1636968456
transform 1 0 13708 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_149
timestamp 1636968456
transform 1 0 14812 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_161
timestamp 1
transform 1 0 15916 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_167
timestamp 1
transform 1 0 16468 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_169
timestamp 1636968456
transform 1 0 16652 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_181
timestamp 1636968456
transform 1 0 17756 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_193
timestamp 1636968456
transform 1 0 18860 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_205
timestamp 1636968456
transform 1 0 19964 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_217
timestamp 1
transform 1 0 21068 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_223
timestamp 1
transform 1 0 21620 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_225
timestamp 1636968456
transform 1 0 21804 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_237
timestamp 1636968456
transform 1 0 22908 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_249
timestamp 1636968456
transform 1 0 24012 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_261
timestamp 1636968456
transform 1 0 25116 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_273
timestamp 1
transform 1 0 26220 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_279
timestamp 1
transform 1 0 26772 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_281
timestamp 1636968456
transform 1 0 26956 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_293
timestamp 1636968456
transform 1 0 28060 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_305
timestamp 1636968456
transform 1 0 29164 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_317
timestamp 1636968456
transform 1 0 30268 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_329
timestamp 1
transform 1 0 31372 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_335
timestamp 1
transform 1 0 31924 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_337
timestamp 1636968456
transform 1 0 32108 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_349
timestamp 1636968456
transform 1 0 33212 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_361
timestamp 1636968456
transform 1 0 34316 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_373
timestamp 1636968456
transform 1 0 35420 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_385
timestamp 1
transform 1 0 36524 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_391
timestamp 1
transform 1 0 37076 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_393
timestamp 1636968456
transform 1 0 37260 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_405
timestamp 1636968456
transform 1 0 38364 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_417
timestamp 1636968456
transform 1 0 39468 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_429
timestamp 1636968456
transform 1 0 40572 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_441
timestamp 1
transform 1 0 41676 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_447
timestamp 1
transform 1 0 42228 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_449
timestamp 1636968456
transform 1 0 42412 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_461
timestamp 1636968456
transform 1 0 43516 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_473
timestamp 1636968456
transform 1 0 44620 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_485
timestamp 1636968456
transform 1 0 45724 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_497
timestamp 1
transform 1 0 46828 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_503
timestamp 1
transform 1 0 47380 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_505
timestamp 1636968456
transform 1 0 47564 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_517
timestamp 1636968456
transform 1 0 48668 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_529
timestamp 1636968456
transform 1 0 49772 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_541
timestamp 1636968456
transform 1 0 50876 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_553
timestamp 1
transform 1 0 51980 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_559
timestamp 1
transform 1 0 52532 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_561
timestamp 1636968456
transform 1 0 52716 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_573
timestamp 1636968456
transform 1 0 53820 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_585
timestamp 1636968456
transform 1 0 54924 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_597
timestamp 1636968456
transform 1 0 56028 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_609
timestamp 1
transform 1 0 57132 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_615
timestamp 1
transform 1 0 57684 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_617
timestamp 1636968456
transform 1 0 57868 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_629
timestamp 1636968456
transform 1 0 58972 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_641
timestamp 1636968456
transform 1 0 60076 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_653
timestamp 1636968456
transform 1 0 61180 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_665
timestamp 1
transform 1 0 62284 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_671
timestamp 1
transform 1 0 62836 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_673
timestamp 1636968456
transform 1 0 63020 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_685
timestamp 1636968456
transform 1 0 64124 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_697
timestamp 1636968456
transform 1 0 65228 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_709
timestamp 1636968456
transform 1 0 66332 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_721
timestamp 1
transform 1 0 67436 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_727
timestamp 1
transform 1 0 67988 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_729
timestamp 1636968456
transform 1 0 68172 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_741
timestamp 1636968456
transform 1 0 69276 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_753
timestamp 1636968456
transform 1 0 70380 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_765
timestamp 1636968456
transform 1 0 71484 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_777
timestamp 1
transform 1 0 72588 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_783
timestamp 1
transform 1 0 73140 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_785
timestamp 1636968456
transform 1 0 73324 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_797
timestamp 1636968456
transform 1 0 74428 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_809
timestamp 1636968456
transform 1 0 75532 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_821
timestamp 1636968456
transform 1 0 76636 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_833
timestamp 1
transform 1 0 77740 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_839
timestamp 1
transform 1 0 78292 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_841
timestamp 1636968456
transform 1 0 78476 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_853
timestamp 1636968456
transform 1 0 79580 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_865
timestamp 1636968456
transform 1 0 80684 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_877
timestamp 1636968456
transform 1 0 81788 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_889
timestamp 1
transform 1 0 82892 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_895
timestamp 1
transform 1 0 83444 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_897
timestamp 1636968456
transform 1 0 83628 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_909
timestamp 1636968456
transform 1 0 84732 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_921
timestamp 1636968456
transform 1 0 85836 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_933
timestamp 1636968456
transform 1 0 86940 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_945
timestamp 1
transform 1 0 88044 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_951
timestamp 1
transform 1 0 88596 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_953
timestamp 1636968456
transform 1 0 88780 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_965
timestamp 1636968456
transform 1 0 89884 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_977
timestamp 1636968456
transform 1 0 90988 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_989
timestamp 1636968456
transform 1 0 92092 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_1001
timestamp 1
transform 1 0 93196 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_1007
timestamp 1
transform 1 0 93748 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1009
timestamp 1636968456
transform 1 0 93932 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1021
timestamp 1636968456
transform 1 0 95036 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1033
timestamp 1636968456
transform 1 0 96140 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1045
timestamp 1636968456
transform 1 0 97244 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_1057
timestamp 1
transform 1 0 98348 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_1063
timestamp 1
transform 1 0 98900 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1065
timestamp 1636968456
transform 1 0 99084 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1077
timestamp 1636968456
transform 1 0 100188 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1089
timestamp 1636968456
transform 1 0 101292 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1101
timestamp 1636968456
transform 1 0 102396 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_1113
timestamp 1
transform 1 0 103500 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_1119
timestamp 1
transform 1 0 104052 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1121
timestamp 1636968456
transform 1 0 104236 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1133
timestamp 1636968456
transform 1 0 105340 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1145
timestamp 1636968456
transform 1 0 106444 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_259_1157
timestamp 1
transform 1 0 107548 0 -1 143616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_259_1165
timestamp 1
transform 1 0 108284 0 -1 143616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_260_3
timestamp 1636968456
transform 1 0 1380 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_15
timestamp 1636968456
transform 1 0 2484 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_260_27
timestamp 1
transform 1 0 3588 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_29
timestamp 1636968456
transform 1 0 3772 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_41
timestamp 1636968456
transform 1 0 4876 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_53
timestamp 1636968456
transform 1 0 5980 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_65
timestamp 1636968456
transform 1 0 7084 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_77
timestamp 1
transform 1 0 8188 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_83
timestamp 1
transform 1 0 8740 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_85
timestamp 1636968456
transform 1 0 8924 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_97
timestamp 1636968456
transform 1 0 10028 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_109
timestamp 1636968456
transform 1 0 11132 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_121
timestamp 1636968456
transform 1 0 12236 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_133
timestamp 1
transform 1 0 13340 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_139
timestamp 1
transform 1 0 13892 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_141
timestamp 1636968456
transform 1 0 14076 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_153
timestamp 1636968456
transform 1 0 15180 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_165
timestamp 1636968456
transform 1 0 16284 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_177
timestamp 1636968456
transform 1 0 17388 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_189
timestamp 1
transform 1 0 18492 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_195
timestamp 1
transform 1 0 19044 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_197
timestamp 1636968456
transform 1 0 19228 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_209
timestamp 1636968456
transform 1 0 20332 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_221
timestamp 1636968456
transform 1 0 21436 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_233
timestamp 1636968456
transform 1 0 22540 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_245
timestamp 1
transform 1 0 23644 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_251
timestamp 1
transform 1 0 24196 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_253
timestamp 1636968456
transform 1 0 24380 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_265
timestamp 1636968456
transform 1 0 25484 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_277
timestamp 1636968456
transform 1 0 26588 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_289
timestamp 1636968456
transform 1 0 27692 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_301
timestamp 1
transform 1 0 28796 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_307
timestamp 1
transform 1 0 29348 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_309
timestamp 1636968456
transform 1 0 29532 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_321
timestamp 1636968456
transform 1 0 30636 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_333
timestamp 1636968456
transform 1 0 31740 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_345
timestamp 1636968456
transform 1 0 32844 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_357
timestamp 1
transform 1 0 33948 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_363
timestamp 1
transform 1 0 34500 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_365
timestamp 1636968456
transform 1 0 34684 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_377
timestamp 1636968456
transform 1 0 35788 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_389
timestamp 1636968456
transform 1 0 36892 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_401
timestamp 1636968456
transform 1 0 37996 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_413
timestamp 1
transform 1 0 39100 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_419
timestamp 1
transform 1 0 39652 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_421
timestamp 1636968456
transform 1 0 39836 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_433
timestamp 1636968456
transform 1 0 40940 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_445
timestamp 1636968456
transform 1 0 42044 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_457
timestamp 1636968456
transform 1 0 43148 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_469
timestamp 1
transform 1 0 44252 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_475
timestamp 1
transform 1 0 44804 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_477
timestamp 1636968456
transform 1 0 44988 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_489
timestamp 1636968456
transform 1 0 46092 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_501
timestamp 1636968456
transform 1 0 47196 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_513
timestamp 1636968456
transform 1 0 48300 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_525
timestamp 1
transform 1 0 49404 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_531
timestamp 1
transform 1 0 49956 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_533
timestamp 1636968456
transform 1 0 50140 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_545
timestamp 1636968456
transform 1 0 51244 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_557
timestamp 1636968456
transform 1 0 52348 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_569
timestamp 1636968456
transform 1 0 53452 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_581
timestamp 1
transform 1 0 54556 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_587
timestamp 1
transform 1 0 55108 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_589
timestamp 1636968456
transform 1 0 55292 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_601
timestamp 1636968456
transform 1 0 56396 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_613
timestamp 1636968456
transform 1 0 57500 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_625
timestamp 1636968456
transform 1 0 58604 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_637
timestamp 1
transform 1 0 59708 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_643
timestamp 1
transform 1 0 60260 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_645
timestamp 1636968456
transform 1 0 60444 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_657
timestamp 1636968456
transform 1 0 61548 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_669
timestamp 1636968456
transform 1 0 62652 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_681
timestamp 1636968456
transform 1 0 63756 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_693
timestamp 1
transform 1 0 64860 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_699
timestamp 1
transform 1 0 65412 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_701
timestamp 1636968456
transform 1 0 65596 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_713
timestamp 1636968456
transform 1 0 66700 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_725
timestamp 1636968456
transform 1 0 67804 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_737
timestamp 1636968456
transform 1 0 68908 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_749
timestamp 1
transform 1 0 70012 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_755
timestamp 1
transform 1 0 70564 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_757
timestamp 1636968456
transform 1 0 70748 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_769
timestamp 1636968456
transform 1 0 71852 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_781
timestamp 1636968456
transform 1 0 72956 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_793
timestamp 1636968456
transform 1 0 74060 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_805
timestamp 1
transform 1 0 75164 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_811
timestamp 1
transform 1 0 75716 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_813
timestamp 1636968456
transform 1 0 75900 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_825
timestamp 1636968456
transform 1 0 77004 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_837
timestamp 1636968456
transform 1 0 78108 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_849
timestamp 1636968456
transform 1 0 79212 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_861
timestamp 1
transform 1 0 80316 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_867
timestamp 1
transform 1 0 80868 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_869
timestamp 1636968456
transform 1 0 81052 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_881
timestamp 1636968456
transform 1 0 82156 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_893
timestamp 1636968456
transform 1 0 83260 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_905
timestamp 1636968456
transform 1 0 84364 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_917
timestamp 1
transform 1 0 85468 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_923
timestamp 1
transform 1 0 86020 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_925
timestamp 1636968456
transform 1 0 86204 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_937
timestamp 1636968456
transform 1 0 87308 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_949
timestamp 1636968456
transform 1 0 88412 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_961
timestamp 1636968456
transform 1 0 89516 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_973
timestamp 1
transform 1 0 90620 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_979
timestamp 1
transform 1 0 91172 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_981
timestamp 1636968456
transform 1 0 91356 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_993
timestamp 1636968456
transform 1 0 92460 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1005
timestamp 1636968456
transform 1 0 93564 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1017
timestamp 1636968456
transform 1 0 94668 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_1029
timestamp 1
transform 1 0 95772 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_1035
timestamp 1
transform 1 0 96324 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1037
timestamp 1636968456
transform 1 0 96508 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1049
timestamp 1636968456
transform 1 0 97612 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1061
timestamp 1636968456
transform 1 0 98716 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1073
timestamp 1636968456
transform 1 0 99820 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_1085
timestamp 1
transform 1 0 100924 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_1091
timestamp 1
transform 1 0 101476 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1093
timestamp 1636968456
transform 1 0 101660 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1105
timestamp 1636968456
transform 1 0 102764 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1117
timestamp 1636968456
transform 1 0 103868 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1129
timestamp 1636968456
transform 1 0 104972 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_1141
timestamp 1
transform 1 0 106076 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_1147
timestamp 1
transform 1 0 106628 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1149
timestamp 1636968456
transform 1 0 106812 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_1161
timestamp 1
transform 1 0 107916 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_1167
timestamp 1
transform 1 0 108468 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_3
timestamp 1636968456
transform 1 0 1380 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_15
timestamp 1636968456
transform 1 0 2484 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_27
timestamp 1636968456
transform 1 0 3588 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_39
timestamp 1636968456
transform 1 0 4692 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_261_51
timestamp 1
transform 1 0 5796 0 -1 144704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_261_55
timestamp 1
transform 1 0 6164 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_57
timestamp 1636968456
transform 1 0 6348 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_69
timestamp 1636968456
transform 1 0 7452 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_81
timestamp 1636968456
transform 1 0 8556 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_93
timestamp 1636968456
transform 1 0 9660 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_105
timestamp 1
transform 1 0 10764 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_111
timestamp 1
transform 1 0 11316 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_113
timestamp 1636968456
transform 1 0 11500 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_125
timestamp 1636968456
transform 1 0 12604 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_137
timestamp 1636968456
transform 1 0 13708 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_149
timestamp 1636968456
transform 1 0 14812 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_161
timestamp 1
transform 1 0 15916 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_167
timestamp 1
transform 1 0 16468 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_169
timestamp 1636968456
transform 1 0 16652 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_181
timestamp 1636968456
transform 1 0 17756 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_193
timestamp 1636968456
transform 1 0 18860 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_205
timestamp 1636968456
transform 1 0 19964 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_217
timestamp 1
transform 1 0 21068 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_223
timestamp 1
transform 1 0 21620 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_225
timestamp 1636968456
transform 1 0 21804 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_237
timestamp 1636968456
transform 1 0 22908 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_249
timestamp 1636968456
transform 1 0 24012 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_261
timestamp 1636968456
transform 1 0 25116 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_273
timestamp 1
transform 1 0 26220 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_279
timestamp 1
transform 1 0 26772 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_281
timestamp 1636968456
transform 1 0 26956 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_293
timestamp 1636968456
transform 1 0 28060 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_305
timestamp 1636968456
transform 1 0 29164 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_317
timestamp 1636968456
transform 1 0 30268 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_329
timestamp 1
transform 1 0 31372 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_335
timestamp 1
transform 1 0 31924 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_337
timestamp 1636968456
transform 1 0 32108 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_349
timestamp 1636968456
transform 1 0 33212 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_361
timestamp 1636968456
transform 1 0 34316 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_373
timestamp 1636968456
transform 1 0 35420 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_385
timestamp 1
transform 1 0 36524 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_391
timestamp 1
transform 1 0 37076 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_393
timestamp 1636968456
transform 1 0 37260 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_405
timestamp 1636968456
transform 1 0 38364 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_417
timestamp 1636968456
transform 1 0 39468 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_429
timestamp 1636968456
transform 1 0 40572 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_441
timestamp 1
transform 1 0 41676 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_447
timestamp 1
transform 1 0 42228 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_449
timestamp 1636968456
transform 1 0 42412 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_461
timestamp 1636968456
transform 1 0 43516 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_473
timestamp 1636968456
transform 1 0 44620 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_485
timestamp 1636968456
transform 1 0 45724 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_497
timestamp 1
transform 1 0 46828 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_503
timestamp 1
transform 1 0 47380 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_505
timestamp 1636968456
transform 1 0 47564 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_517
timestamp 1636968456
transform 1 0 48668 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_529
timestamp 1636968456
transform 1 0 49772 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_541
timestamp 1636968456
transform 1 0 50876 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_553
timestamp 1
transform 1 0 51980 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_559
timestamp 1
transform 1 0 52532 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_561
timestamp 1636968456
transform 1 0 52716 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_573
timestamp 1636968456
transform 1 0 53820 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_585
timestamp 1636968456
transform 1 0 54924 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_597
timestamp 1636968456
transform 1 0 56028 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_609
timestamp 1
transform 1 0 57132 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_615
timestamp 1
transform 1 0 57684 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_617
timestamp 1636968456
transform 1 0 57868 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_629
timestamp 1636968456
transform 1 0 58972 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_641
timestamp 1636968456
transform 1 0 60076 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_653
timestamp 1636968456
transform 1 0 61180 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_665
timestamp 1
transform 1 0 62284 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_671
timestamp 1
transform 1 0 62836 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_673
timestamp 1636968456
transform 1 0 63020 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_685
timestamp 1636968456
transform 1 0 64124 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_697
timestamp 1636968456
transform 1 0 65228 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_709
timestamp 1636968456
transform 1 0 66332 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_721
timestamp 1
transform 1 0 67436 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_727
timestamp 1
transform 1 0 67988 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_729
timestamp 1636968456
transform 1 0 68172 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_741
timestamp 1636968456
transform 1 0 69276 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_753
timestamp 1636968456
transform 1 0 70380 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_765
timestamp 1636968456
transform 1 0 71484 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_777
timestamp 1
transform 1 0 72588 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_783
timestamp 1
transform 1 0 73140 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_785
timestamp 1636968456
transform 1 0 73324 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_797
timestamp 1636968456
transform 1 0 74428 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_809
timestamp 1636968456
transform 1 0 75532 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_821
timestamp 1636968456
transform 1 0 76636 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_833
timestamp 1
transform 1 0 77740 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_839
timestamp 1
transform 1 0 78292 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_841
timestamp 1636968456
transform 1 0 78476 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_853
timestamp 1636968456
transform 1 0 79580 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_865
timestamp 1636968456
transform 1 0 80684 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_877
timestamp 1636968456
transform 1 0 81788 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_889
timestamp 1
transform 1 0 82892 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_895
timestamp 1
transform 1 0 83444 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_897
timestamp 1636968456
transform 1 0 83628 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_909
timestamp 1636968456
transform 1 0 84732 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_921
timestamp 1636968456
transform 1 0 85836 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_933
timestamp 1636968456
transform 1 0 86940 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_945
timestamp 1
transform 1 0 88044 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_951
timestamp 1
transform 1 0 88596 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_953
timestamp 1636968456
transform 1 0 88780 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_965
timestamp 1636968456
transform 1 0 89884 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_977
timestamp 1636968456
transform 1 0 90988 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_989
timestamp 1636968456
transform 1 0 92092 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_1001
timestamp 1
transform 1 0 93196 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_1007
timestamp 1
transform 1 0 93748 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1009
timestamp 1636968456
transform 1 0 93932 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1021
timestamp 1636968456
transform 1 0 95036 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1033
timestamp 1636968456
transform 1 0 96140 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1045
timestamp 1636968456
transform 1 0 97244 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_1057
timestamp 1
transform 1 0 98348 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_1063
timestamp 1
transform 1 0 98900 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1065
timestamp 1636968456
transform 1 0 99084 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1077
timestamp 1636968456
transform 1 0 100188 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1089
timestamp 1636968456
transform 1 0 101292 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1101
timestamp 1636968456
transform 1 0 102396 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_1113
timestamp 1
transform 1 0 103500 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_1119
timestamp 1
transform 1 0 104052 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1121
timestamp 1636968456
transform 1 0 104236 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1133
timestamp 1636968456
transform 1 0 105340 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1145
timestamp 1636968456
transform 1 0 106444 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_261_1157
timestamp 1
transform 1 0 107548 0 -1 144704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_261_1165
timestamp 1
transform 1 0 108284 0 -1 144704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_262_3
timestamp 1636968456
transform 1 0 1380 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_15
timestamp 1636968456
transform 1 0 2484 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_262_27
timestamp 1
transform 1 0 3588 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_29
timestamp 1636968456
transform 1 0 3772 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_41
timestamp 1636968456
transform 1 0 4876 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_53
timestamp 1636968456
transform 1 0 5980 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_65
timestamp 1636968456
transform 1 0 7084 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_77
timestamp 1
transform 1 0 8188 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_83
timestamp 1
transform 1 0 8740 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_85
timestamp 1636968456
transform 1 0 8924 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_97
timestamp 1636968456
transform 1 0 10028 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_109
timestamp 1636968456
transform 1 0 11132 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_121
timestamp 1636968456
transform 1 0 12236 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_133
timestamp 1
transform 1 0 13340 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_139
timestamp 1
transform 1 0 13892 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_141
timestamp 1636968456
transform 1 0 14076 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_153
timestamp 1636968456
transform 1 0 15180 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_165
timestamp 1636968456
transform 1 0 16284 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_177
timestamp 1636968456
transform 1 0 17388 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_189
timestamp 1
transform 1 0 18492 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_195
timestamp 1
transform 1 0 19044 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_197
timestamp 1636968456
transform 1 0 19228 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_209
timestamp 1636968456
transform 1 0 20332 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_221
timestamp 1636968456
transform 1 0 21436 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_233
timestamp 1636968456
transform 1 0 22540 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_245
timestamp 1
transform 1 0 23644 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_251
timestamp 1
transform 1 0 24196 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_253
timestamp 1636968456
transform 1 0 24380 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_265
timestamp 1636968456
transform 1 0 25484 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_277
timestamp 1636968456
transform 1 0 26588 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_289
timestamp 1636968456
transform 1 0 27692 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_301
timestamp 1
transform 1 0 28796 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_307
timestamp 1
transform 1 0 29348 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_309
timestamp 1636968456
transform 1 0 29532 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_321
timestamp 1636968456
transform 1 0 30636 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_333
timestamp 1636968456
transform 1 0 31740 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_345
timestamp 1636968456
transform 1 0 32844 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_357
timestamp 1
transform 1 0 33948 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_363
timestamp 1
transform 1 0 34500 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_365
timestamp 1636968456
transform 1 0 34684 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_377
timestamp 1636968456
transform 1 0 35788 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_389
timestamp 1636968456
transform 1 0 36892 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_401
timestamp 1636968456
transform 1 0 37996 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_413
timestamp 1
transform 1 0 39100 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_419
timestamp 1
transform 1 0 39652 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_421
timestamp 1636968456
transform 1 0 39836 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_433
timestamp 1636968456
transform 1 0 40940 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_445
timestamp 1636968456
transform 1 0 42044 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_457
timestamp 1636968456
transform 1 0 43148 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_469
timestamp 1
transform 1 0 44252 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_475
timestamp 1
transform 1 0 44804 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_477
timestamp 1636968456
transform 1 0 44988 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_489
timestamp 1636968456
transform 1 0 46092 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_501
timestamp 1636968456
transform 1 0 47196 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_513
timestamp 1636968456
transform 1 0 48300 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_525
timestamp 1
transform 1 0 49404 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_531
timestamp 1
transform 1 0 49956 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_533
timestamp 1636968456
transform 1 0 50140 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_545
timestamp 1636968456
transform 1 0 51244 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_557
timestamp 1636968456
transform 1 0 52348 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_569
timestamp 1636968456
transform 1 0 53452 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_581
timestamp 1
transform 1 0 54556 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_587
timestamp 1
transform 1 0 55108 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_589
timestamp 1636968456
transform 1 0 55292 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_601
timestamp 1636968456
transform 1 0 56396 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_613
timestamp 1636968456
transform 1 0 57500 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_625
timestamp 1636968456
transform 1 0 58604 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_637
timestamp 1
transform 1 0 59708 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_643
timestamp 1
transform 1 0 60260 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_645
timestamp 1636968456
transform 1 0 60444 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_657
timestamp 1636968456
transform 1 0 61548 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_669
timestamp 1636968456
transform 1 0 62652 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_681
timestamp 1636968456
transform 1 0 63756 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_693
timestamp 1
transform 1 0 64860 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_699
timestamp 1
transform 1 0 65412 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_701
timestamp 1636968456
transform 1 0 65596 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_713
timestamp 1636968456
transform 1 0 66700 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_725
timestamp 1636968456
transform 1 0 67804 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_737
timestamp 1636968456
transform 1 0 68908 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_749
timestamp 1
transform 1 0 70012 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_755
timestamp 1
transform 1 0 70564 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_757
timestamp 1636968456
transform 1 0 70748 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_769
timestamp 1636968456
transform 1 0 71852 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_781
timestamp 1636968456
transform 1 0 72956 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_793
timestamp 1636968456
transform 1 0 74060 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_805
timestamp 1
transform 1 0 75164 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_811
timestamp 1
transform 1 0 75716 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_813
timestamp 1636968456
transform 1 0 75900 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_825
timestamp 1636968456
transform 1 0 77004 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_837
timestamp 1636968456
transform 1 0 78108 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_849
timestamp 1636968456
transform 1 0 79212 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_861
timestamp 1
transform 1 0 80316 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_867
timestamp 1
transform 1 0 80868 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_869
timestamp 1636968456
transform 1 0 81052 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_881
timestamp 1636968456
transform 1 0 82156 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_893
timestamp 1636968456
transform 1 0 83260 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_905
timestamp 1636968456
transform 1 0 84364 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_917
timestamp 1
transform 1 0 85468 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_923
timestamp 1
transform 1 0 86020 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_925
timestamp 1636968456
transform 1 0 86204 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_937
timestamp 1636968456
transform 1 0 87308 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_949
timestamp 1636968456
transform 1 0 88412 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_961
timestamp 1636968456
transform 1 0 89516 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_973
timestamp 1
transform 1 0 90620 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_979
timestamp 1
transform 1 0 91172 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_981
timestamp 1636968456
transform 1 0 91356 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_993
timestamp 1636968456
transform 1 0 92460 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1005
timestamp 1636968456
transform 1 0 93564 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1017
timestamp 1636968456
transform 1 0 94668 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_1029
timestamp 1
transform 1 0 95772 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_1035
timestamp 1
transform 1 0 96324 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1037
timestamp 1636968456
transform 1 0 96508 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1049
timestamp 1636968456
transform 1 0 97612 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1061
timestamp 1636968456
transform 1 0 98716 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1073
timestamp 1636968456
transform 1 0 99820 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_1085
timestamp 1
transform 1 0 100924 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_1091
timestamp 1
transform 1 0 101476 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1093
timestamp 1636968456
transform 1 0 101660 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1105
timestamp 1636968456
transform 1 0 102764 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1117
timestamp 1636968456
transform 1 0 103868 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1129
timestamp 1636968456
transform 1 0 104972 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_1141
timestamp 1
transform 1 0 106076 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_1147
timestamp 1
transform 1 0 106628 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1149
timestamp 1636968456
transform 1 0 106812 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_1161
timestamp 1
transform 1 0 107916 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_1167
timestamp 1
transform 1 0 108468 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_3
timestamp 1636968456
transform 1 0 1380 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_15
timestamp 1636968456
transform 1 0 2484 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_27
timestamp 1636968456
transform 1 0 3588 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_39
timestamp 1636968456
transform 1 0 4692 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_263_51
timestamp 1
transform 1 0 5796 0 -1 145792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_263_55
timestamp 1
transform 1 0 6164 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_57
timestamp 1636968456
transform 1 0 6348 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_69
timestamp 1636968456
transform 1 0 7452 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_81
timestamp 1636968456
transform 1 0 8556 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_93
timestamp 1636968456
transform 1 0 9660 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_105
timestamp 1
transform 1 0 10764 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_111
timestamp 1
transform 1 0 11316 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_113
timestamp 1636968456
transform 1 0 11500 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_125
timestamp 1636968456
transform 1 0 12604 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_137
timestamp 1636968456
transform 1 0 13708 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_149
timestamp 1636968456
transform 1 0 14812 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_161
timestamp 1
transform 1 0 15916 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_167
timestamp 1
transform 1 0 16468 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_169
timestamp 1636968456
transform 1 0 16652 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_181
timestamp 1636968456
transform 1 0 17756 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_193
timestamp 1636968456
transform 1 0 18860 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_205
timestamp 1636968456
transform 1 0 19964 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_217
timestamp 1
transform 1 0 21068 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_223
timestamp 1
transform 1 0 21620 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_225
timestamp 1636968456
transform 1 0 21804 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_237
timestamp 1636968456
transform 1 0 22908 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_249
timestamp 1636968456
transform 1 0 24012 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_261
timestamp 1636968456
transform 1 0 25116 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_273
timestamp 1
transform 1 0 26220 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_279
timestamp 1
transform 1 0 26772 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_281
timestamp 1636968456
transform 1 0 26956 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_293
timestamp 1636968456
transform 1 0 28060 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_305
timestamp 1636968456
transform 1 0 29164 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_317
timestamp 1636968456
transform 1 0 30268 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_329
timestamp 1
transform 1 0 31372 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_335
timestamp 1
transform 1 0 31924 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_337
timestamp 1636968456
transform 1 0 32108 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_349
timestamp 1636968456
transform 1 0 33212 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_361
timestamp 1636968456
transform 1 0 34316 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_373
timestamp 1636968456
transform 1 0 35420 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_385
timestamp 1
transform 1 0 36524 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_391
timestamp 1
transform 1 0 37076 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_393
timestamp 1636968456
transform 1 0 37260 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_405
timestamp 1636968456
transform 1 0 38364 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_417
timestamp 1636968456
transform 1 0 39468 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_429
timestamp 1636968456
transform 1 0 40572 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_441
timestamp 1
transform 1 0 41676 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_447
timestamp 1
transform 1 0 42228 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_449
timestamp 1636968456
transform 1 0 42412 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_461
timestamp 1636968456
transform 1 0 43516 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_473
timestamp 1636968456
transform 1 0 44620 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_485
timestamp 1636968456
transform 1 0 45724 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_497
timestamp 1
transform 1 0 46828 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_503
timestamp 1
transform 1 0 47380 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_505
timestamp 1636968456
transform 1 0 47564 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_517
timestamp 1636968456
transform 1 0 48668 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_529
timestamp 1636968456
transform 1 0 49772 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_541
timestamp 1636968456
transform 1 0 50876 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_553
timestamp 1
transform 1 0 51980 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_559
timestamp 1
transform 1 0 52532 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_561
timestamp 1636968456
transform 1 0 52716 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_573
timestamp 1636968456
transform 1 0 53820 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_585
timestamp 1636968456
transform 1 0 54924 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_597
timestamp 1636968456
transform 1 0 56028 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_609
timestamp 1
transform 1 0 57132 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_615
timestamp 1
transform 1 0 57684 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_617
timestamp 1636968456
transform 1 0 57868 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_629
timestamp 1636968456
transform 1 0 58972 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_641
timestamp 1636968456
transform 1 0 60076 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_653
timestamp 1636968456
transform 1 0 61180 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_665
timestamp 1
transform 1 0 62284 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_671
timestamp 1
transform 1 0 62836 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_673
timestamp 1636968456
transform 1 0 63020 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_685
timestamp 1636968456
transform 1 0 64124 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_697
timestamp 1636968456
transform 1 0 65228 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_709
timestamp 1636968456
transform 1 0 66332 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_721
timestamp 1
transform 1 0 67436 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_727
timestamp 1
transform 1 0 67988 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_729
timestamp 1636968456
transform 1 0 68172 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_741
timestamp 1636968456
transform 1 0 69276 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_753
timestamp 1636968456
transform 1 0 70380 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_765
timestamp 1636968456
transform 1 0 71484 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_777
timestamp 1
transform 1 0 72588 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_783
timestamp 1
transform 1 0 73140 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_785
timestamp 1636968456
transform 1 0 73324 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_797
timestamp 1636968456
transform 1 0 74428 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_809
timestamp 1636968456
transform 1 0 75532 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_821
timestamp 1636968456
transform 1 0 76636 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_833
timestamp 1
transform 1 0 77740 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_839
timestamp 1
transform 1 0 78292 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_841
timestamp 1636968456
transform 1 0 78476 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_853
timestamp 1636968456
transform 1 0 79580 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_865
timestamp 1636968456
transform 1 0 80684 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_877
timestamp 1636968456
transform 1 0 81788 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_889
timestamp 1
transform 1 0 82892 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_895
timestamp 1
transform 1 0 83444 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_897
timestamp 1636968456
transform 1 0 83628 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_909
timestamp 1636968456
transform 1 0 84732 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_921
timestamp 1636968456
transform 1 0 85836 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_933
timestamp 1636968456
transform 1 0 86940 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_945
timestamp 1
transform 1 0 88044 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_951
timestamp 1
transform 1 0 88596 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_953
timestamp 1636968456
transform 1 0 88780 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_965
timestamp 1636968456
transform 1 0 89884 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_977
timestamp 1636968456
transform 1 0 90988 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_989
timestamp 1636968456
transform 1 0 92092 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_1001
timestamp 1
transform 1 0 93196 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_1007
timestamp 1
transform 1 0 93748 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1009
timestamp 1636968456
transform 1 0 93932 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1021
timestamp 1636968456
transform 1 0 95036 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1033
timestamp 1636968456
transform 1 0 96140 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1045
timestamp 1636968456
transform 1 0 97244 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_1057
timestamp 1
transform 1 0 98348 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_1063
timestamp 1
transform 1 0 98900 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1065
timestamp 1636968456
transform 1 0 99084 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1077
timestamp 1636968456
transform 1 0 100188 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1089
timestamp 1636968456
transform 1 0 101292 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1101
timestamp 1636968456
transform 1 0 102396 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_1113
timestamp 1
transform 1 0 103500 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_1119
timestamp 1
transform 1 0 104052 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1121
timestamp 1636968456
transform 1 0 104236 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1133
timestamp 1636968456
transform 1 0 105340 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1145
timestamp 1636968456
transform 1 0 106444 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_263_1157
timestamp 1
transform 1 0 107548 0 -1 145792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_263_1165
timestamp 1
transform 1 0 108284 0 -1 145792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_264_3
timestamp 1636968456
transform 1 0 1380 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_15
timestamp 1636968456
transform 1 0 2484 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_264_27
timestamp 1
transform 1 0 3588 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_29
timestamp 1636968456
transform 1 0 3772 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_41
timestamp 1636968456
transform 1 0 4876 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_53
timestamp 1636968456
transform 1 0 5980 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_65
timestamp 1636968456
transform 1 0 7084 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_77
timestamp 1
transform 1 0 8188 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_83
timestamp 1
transform 1 0 8740 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_85
timestamp 1636968456
transform 1 0 8924 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_97
timestamp 1636968456
transform 1 0 10028 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_109
timestamp 1636968456
transform 1 0 11132 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_121
timestamp 1636968456
transform 1 0 12236 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_133
timestamp 1
transform 1 0 13340 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_139
timestamp 1
transform 1 0 13892 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_141
timestamp 1636968456
transform 1 0 14076 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_153
timestamp 1636968456
transform 1 0 15180 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_165
timestamp 1636968456
transform 1 0 16284 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_177
timestamp 1636968456
transform 1 0 17388 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_189
timestamp 1
transform 1 0 18492 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_195
timestamp 1
transform 1 0 19044 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_197
timestamp 1636968456
transform 1 0 19228 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_209
timestamp 1636968456
transform 1 0 20332 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_221
timestamp 1636968456
transform 1 0 21436 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_233
timestamp 1636968456
transform 1 0 22540 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_245
timestamp 1
transform 1 0 23644 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_251
timestamp 1
transform 1 0 24196 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_253
timestamp 1636968456
transform 1 0 24380 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_265
timestamp 1636968456
transform 1 0 25484 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_277
timestamp 1636968456
transform 1 0 26588 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_289
timestamp 1636968456
transform 1 0 27692 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_301
timestamp 1
transform 1 0 28796 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_307
timestamp 1
transform 1 0 29348 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_309
timestamp 1636968456
transform 1 0 29532 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_321
timestamp 1636968456
transform 1 0 30636 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_333
timestamp 1636968456
transform 1 0 31740 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_345
timestamp 1636968456
transform 1 0 32844 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_357
timestamp 1
transform 1 0 33948 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_363
timestamp 1
transform 1 0 34500 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_365
timestamp 1636968456
transform 1 0 34684 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_377
timestamp 1636968456
transform 1 0 35788 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_389
timestamp 1636968456
transform 1 0 36892 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_401
timestamp 1636968456
transform 1 0 37996 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_413
timestamp 1
transform 1 0 39100 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_419
timestamp 1
transform 1 0 39652 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_421
timestamp 1636968456
transform 1 0 39836 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_433
timestamp 1636968456
transform 1 0 40940 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_445
timestamp 1636968456
transform 1 0 42044 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_457
timestamp 1636968456
transform 1 0 43148 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_469
timestamp 1
transform 1 0 44252 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_475
timestamp 1
transform 1 0 44804 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_477
timestamp 1636968456
transform 1 0 44988 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_489
timestamp 1636968456
transform 1 0 46092 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_501
timestamp 1636968456
transform 1 0 47196 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_513
timestamp 1636968456
transform 1 0 48300 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_525
timestamp 1
transform 1 0 49404 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_531
timestamp 1
transform 1 0 49956 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_533
timestamp 1636968456
transform 1 0 50140 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_545
timestamp 1636968456
transform 1 0 51244 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_557
timestamp 1636968456
transform 1 0 52348 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_569
timestamp 1636968456
transform 1 0 53452 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_581
timestamp 1
transform 1 0 54556 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_587
timestamp 1
transform 1 0 55108 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_589
timestamp 1636968456
transform 1 0 55292 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_601
timestamp 1636968456
transform 1 0 56396 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_613
timestamp 1636968456
transform 1 0 57500 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_625
timestamp 1636968456
transform 1 0 58604 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_637
timestamp 1
transform 1 0 59708 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_643
timestamp 1
transform 1 0 60260 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_645
timestamp 1636968456
transform 1 0 60444 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_657
timestamp 1636968456
transform 1 0 61548 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_669
timestamp 1636968456
transform 1 0 62652 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_681
timestamp 1636968456
transform 1 0 63756 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_693
timestamp 1
transform 1 0 64860 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_699
timestamp 1
transform 1 0 65412 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_701
timestamp 1636968456
transform 1 0 65596 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_713
timestamp 1636968456
transform 1 0 66700 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_725
timestamp 1636968456
transform 1 0 67804 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_737
timestamp 1636968456
transform 1 0 68908 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_749
timestamp 1
transform 1 0 70012 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_755
timestamp 1
transform 1 0 70564 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_757
timestamp 1636968456
transform 1 0 70748 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_769
timestamp 1636968456
transform 1 0 71852 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_781
timestamp 1636968456
transform 1 0 72956 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_793
timestamp 1636968456
transform 1 0 74060 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_805
timestamp 1
transform 1 0 75164 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_811
timestamp 1
transform 1 0 75716 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_813
timestamp 1636968456
transform 1 0 75900 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_825
timestamp 1636968456
transform 1 0 77004 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_837
timestamp 1636968456
transform 1 0 78108 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_849
timestamp 1636968456
transform 1 0 79212 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_861
timestamp 1
transform 1 0 80316 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_867
timestamp 1
transform 1 0 80868 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_869
timestamp 1636968456
transform 1 0 81052 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_881
timestamp 1636968456
transform 1 0 82156 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_893
timestamp 1636968456
transform 1 0 83260 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_905
timestamp 1636968456
transform 1 0 84364 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_917
timestamp 1
transform 1 0 85468 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_923
timestamp 1
transform 1 0 86020 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_925
timestamp 1636968456
transform 1 0 86204 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_937
timestamp 1636968456
transform 1 0 87308 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_949
timestamp 1636968456
transform 1 0 88412 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_961
timestamp 1636968456
transform 1 0 89516 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_973
timestamp 1
transform 1 0 90620 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_979
timestamp 1
transform 1 0 91172 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_981
timestamp 1636968456
transform 1 0 91356 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_993
timestamp 1636968456
transform 1 0 92460 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1005
timestamp 1636968456
transform 1 0 93564 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1017
timestamp 1636968456
transform 1 0 94668 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_1029
timestamp 1
transform 1 0 95772 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_1035
timestamp 1
transform 1 0 96324 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1037
timestamp 1636968456
transform 1 0 96508 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1049
timestamp 1636968456
transform 1 0 97612 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1061
timestamp 1636968456
transform 1 0 98716 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1073
timestamp 1636968456
transform 1 0 99820 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_1085
timestamp 1
transform 1 0 100924 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_1091
timestamp 1
transform 1 0 101476 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1093
timestamp 1636968456
transform 1 0 101660 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1105
timestamp 1636968456
transform 1 0 102764 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1117
timestamp 1636968456
transform 1 0 103868 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1129
timestamp 1636968456
transform 1 0 104972 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_1141
timestamp 1
transform 1 0 106076 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_1147
timestamp 1
transform 1 0 106628 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1149
timestamp 1636968456
transform 1 0 106812 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_1161
timestamp 1
transform 1 0 107916 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_1167
timestamp 1
transform 1 0 108468 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_3
timestamp 1636968456
transform 1 0 1380 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_15
timestamp 1636968456
transform 1 0 2484 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_27
timestamp 1636968456
transform 1 0 3588 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_39
timestamp 1636968456
transform 1 0 4692 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_265_51
timestamp 1
transform 1 0 5796 0 -1 146880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_265_55
timestamp 1
transform 1 0 6164 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_57
timestamp 1636968456
transform 1 0 6348 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_69
timestamp 1636968456
transform 1 0 7452 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_81
timestamp 1636968456
transform 1 0 8556 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_93
timestamp 1636968456
transform 1 0 9660 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_105
timestamp 1
transform 1 0 10764 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_111
timestamp 1
transform 1 0 11316 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_113
timestamp 1636968456
transform 1 0 11500 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_125
timestamp 1636968456
transform 1 0 12604 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_137
timestamp 1636968456
transform 1 0 13708 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_149
timestamp 1636968456
transform 1 0 14812 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_161
timestamp 1
transform 1 0 15916 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_167
timestamp 1
transform 1 0 16468 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_169
timestamp 1636968456
transform 1 0 16652 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_181
timestamp 1636968456
transform 1 0 17756 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_193
timestamp 1636968456
transform 1 0 18860 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_205
timestamp 1636968456
transform 1 0 19964 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_217
timestamp 1
transform 1 0 21068 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_223
timestamp 1
transform 1 0 21620 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_225
timestamp 1636968456
transform 1 0 21804 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_237
timestamp 1636968456
transform 1 0 22908 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_249
timestamp 1636968456
transform 1 0 24012 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_261
timestamp 1636968456
transform 1 0 25116 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_273
timestamp 1
transform 1 0 26220 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_279
timestamp 1
transform 1 0 26772 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_281
timestamp 1636968456
transform 1 0 26956 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_293
timestamp 1636968456
transform 1 0 28060 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_305
timestamp 1636968456
transform 1 0 29164 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_317
timestamp 1636968456
transform 1 0 30268 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_329
timestamp 1
transform 1 0 31372 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_335
timestamp 1
transform 1 0 31924 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_337
timestamp 1636968456
transform 1 0 32108 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_349
timestamp 1636968456
transform 1 0 33212 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_361
timestamp 1636968456
transform 1 0 34316 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_373
timestamp 1636968456
transform 1 0 35420 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_385
timestamp 1
transform 1 0 36524 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_391
timestamp 1
transform 1 0 37076 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_393
timestamp 1636968456
transform 1 0 37260 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_405
timestamp 1636968456
transform 1 0 38364 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_417
timestamp 1636968456
transform 1 0 39468 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_429
timestamp 1636968456
transform 1 0 40572 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_441
timestamp 1
transform 1 0 41676 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_447
timestamp 1
transform 1 0 42228 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_449
timestamp 1636968456
transform 1 0 42412 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_461
timestamp 1636968456
transform 1 0 43516 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_473
timestamp 1636968456
transform 1 0 44620 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_485
timestamp 1636968456
transform 1 0 45724 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_497
timestamp 1
transform 1 0 46828 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_503
timestamp 1
transform 1 0 47380 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_505
timestamp 1636968456
transform 1 0 47564 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_517
timestamp 1636968456
transform 1 0 48668 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_529
timestamp 1636968456
transform 1 0 49772 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_541
timestamp 1636968456
transform 1 0 50876 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_553
timestamp 1
transform 1 0 51980 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_559
timestamp 1
transform 1 0 52532 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_561
timestamp 1636968456
transform 1 0 52716 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_573
timestamp 1636968456
transform 1 0 53820 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_585
timestamp 1636968456
transform 1 0 54924 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_597
timestamp 1636968456
transform 1 0 56028 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_609
timestamp 1
transform 1 0 57132 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_615
timestamp 1
transform 1 0 57684 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_617
timestamp 1636968456
transform 1 0 57868 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_629
timestamp 1636968456
transform 1 0 58972 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_641
timestamp 1636968456
transform 1 0 60076 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_653
timestamp 1636968456
transform 1 0 61180 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_665
timestamp 1
transform 1 0 62284 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_671
timestamp 1
transform 1 0 62836 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_673
timestamp 1636968456
transform 1 0 63020 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_685
timestamp 1636968456
transform 1 0 64124 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_697
timestamp 1636968456
transform 1 0 65228 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_709
timestamp 1636968456
transform 1 0 66332 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_721
timestamp 1
transform 1 0 67436 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_727
timestamp 1
transform 1 0 67988 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_729
timestamp 1636968456
transform 1 0 68172 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_741
timestamp 1636968456
transform 1 0 69276 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_753
timestamp 1636968456
transform 1 0 70380 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_765
timestamp 1636968456
transform 1 0 71484 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_777
timestamp 1
transform 1 0 72588 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_783
timestamp 1
transform 1 0 73140 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_785
timestamp 1636968456
transform 1 0 73324 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_797
timestamp 1636968456
transform 1 0 74428 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_809
timestamp 1636968456
transform 1 0 75532 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_821
timestamp 1636968456
transform 1 0 76636 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_833
timestamp 1
transform 1 0 77740 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_839
timestamp 1
transform 1 0 78292 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_841
timestamp 1636968456
transform 1 0 78476 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_853
timestamp 1636968456
transform 1 0 79580 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_865
timestamp 1636968456
transform 1 0 80684 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_877
timestamp 1636968456
transform 1 0 81788 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_889
timestamp 1
transform 1 0 82892 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_895
timestamp 1
transform 1 0 83444 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_897
timestamp 1636968456
transform 1 0 83628 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_909
timestamp 1636968456
transform 1 0 84732 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_921
timestamp 1636968456
transform 1 0 85836 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_933
timestamp 1636968456
transform 1 0 86940 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_945
timestamp 1
transform 1 0 88044 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_951
timestamp 1
transform 1 0 88596 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_953
timestamp 1636968456
transform 1 0 88780 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_965
timestamp 1636968456
transform 1 0 89884 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_977
timestamp 1636968456
transform 1 0 90988 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_989
timestamp 1636968456
transform 1 0 92092 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_1001
timestamp 1
transform 1 0 93196 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_1007
timestamp 1
transform 1 0 93748 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1009
timestamp 1636968456
transform 1 0 93932 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1021
timestamp 1636968456
transform 1 0 95036 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1033
timestamp 1636968456
transform 1 0 96140 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1045
timestamp 1636968456
transform 1 0 97244 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_1057
timestamp 1
transform 1 0 98348 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_1063
timestamp 1
transform 1 0 98900 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1065
timestamp 1636968456
transform 1 0 99084 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1077
timestamp 1636968456
transform 1 0 100188 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1089
timestamp 1636968456
transform 1 0 101292 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1101
timestamp 1636968456
transform 1 0 102396 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_1113
timestamp 1
transform 1 0 103500 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_1119
timestamp 1
transform 1 0 104052 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1121
timestamp 1636968456
transform 1 0 104236 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1133
timestamp 1636968456
transform 1 0 105340 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1145
timestamp 1636968456
transform 1 0 106444 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_265_1157
timestamp 1
transform 1 0 107548 0 -1 146880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_265_1165
timestamp 1
transform 1 0 108284 0 -1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_3
timestamp 1636968456
transform 1 0 1380 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_15
timestamp 1636968456
transform 1 0 2484 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_266_27
timestamp 1
transform 1 0 3588 0 1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_266_29
timestamp 1636968456
transform 1 0 3772 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_41
timestamp 1636968456
transform 1 0 4876 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_53
timestamp 1
transform 1 0 5980 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_57
timestamp 1636968456
transform 1 0 6348 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_69
timestamp 1636968456
transform 1 0 7452 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_81
timestamp 1
transform 1 0 8556 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_85
timestamp 1636968456
transform 1 0 8924 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_97
timestamp 1636968456
transform 1 0 10028 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_109
timestamp 1
transform 1 0 11132 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_113
timestamp 1636968456
transform 1 0 11500 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_125
timestamp 1636968456
transform 1 0 12604 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_137
timestamp 1
transform 1 0 13708 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_141
timestamp 1636968456
transform 1 0 14076 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_153
timestamp 1636968456
transform 1 0 15180 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_165
timestamp 1
transform 1 0 16284 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_169
timestamp 1636968456
transform 1 0 16652 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_181
timestamp 1636968456
transform 1 0 17756 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_193
timestamp 1
transform 1 0 18860 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_197
timestamp 1636968456
transform 1 0 19228 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_209
timestamp 1636968456
transform 1 0 20332 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_221
timestamp 1
transform 1 0 21436 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_225
timestamp 1636968456
transform 1 0 21804 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_237
timestamp 1636968456
transform 1 0 22908 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_249
timestamp 1
transform 1 0 24012 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_253
timestamp 1636968456
transform 1 0 24380 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_265
timestamp 1636968456
transform 1 0 25484 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_277
timestamp 1
transform 1 0 26588 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_281
timestamp 1636968456
transform 1 0 26956 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_293
timestamp 1636968456
transform 1 0 28060 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_305
timestamp 1
transform 1 0 29164 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_309
timestamp 1636968456
transform 1 0 29532 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_321
timestamp 1636968456
transform 1 0 30636 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_333
timestamp 1
transform 1 0 31740 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_337
timestamp 1636968456
transform 1 0 32108 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_349
timestamp 1636968456
transform 1 0 33212 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_361
timestamp 1
transform 1 0 34316 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_365
timestamp 1636968456
transform 1 0 34684 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_377
timestamp 1636968456
transform 1 0 35788 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_389
timestamp 1
transform 1 0 36892 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_393
timestamp 1636968456
transform 1 0 37260 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_405
timestamp 1636968456
transform 1 0 38364 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_417
timestamp 1
transform 1 0 39468 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_421
timestamp 1636968456
transform 1 0 39836 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_433
timestamp 1636968456
transform 1 0 40940 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_445
timestamp 1
transform 1 0 42044 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_449
timestamp 1636968456
transform 1 0 42412 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_461
timestamp 1636968456
transform 1 0 43516 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_473
timestamp 1
transform 1 0 44620 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_477
timestamp 1636968456
transform 1 0 44988 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_489
timestamp 1636968456
transform 1 0 46092 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_501
timestamp 1
transform 1 0 47196 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_505
timestamp 1636968456
transform 1 0 47564 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_517
timestamp 1636968456
transform 1 0 48668 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_529
timestamp 1
transform 1 0 49772 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_533
timestamp 1636968456
transform 1 0 50140 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_545
timestamp 1636968456
transform 1 0 51244 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_557
timestamp 1
transform 1 0 52348 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_561
timestamp 1636968456
transform 1 0 52716 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_573
timestamp 1636968456
transform 1 0 53820 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_585
timestamp 1
transform 1 0 54924 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_589
timestamp 1636968456
transform 1 0 55292 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_601
timestamp 1636968456
transform 1 0 56396 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_613
timestamp 1
transform 1 0 57500 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_617
timestamp 1636968456
transform 1 0 57868 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_629
timestamp 1636968456
transform 1 0 58972 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_641
timestamp 1
transform 1 0 60076 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_645
timestamp 1636968456
transform 1 0 60444 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_657
timestamp 1636968456
transform 1 0 61548 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_669
timestamp 1
transform 1 0 62652 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_673
timestamp 1636968456
transform 1 0 63020 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_685
timestamp 1636968456
transform 1 0 64124 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_697
timestamp 1
transform 1 0 65228 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_701
timestamp 1636968456
transform 1 0 65596 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_713
timestamp 1636968456
transform 1 0 66700 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_725
timestamp 1
transform 1 0 67804 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_729
timestamp 1636968456
transform 1 0 68172 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_741
timestamp 1636968456
transform 1 0 69276 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_753
timestamp 1
transform 1 0 70380 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_757
timestamp 1636968456
transform 1 0 70748 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_769
timestamp 1636968456
transform 1 0 71852 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_781
timestamp 1
transform 1 0 72956 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_785
timestamp 1636968456
transform 1 0 73324 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_797
timestamp 1636968456
transform 1 0 74428 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_809
timestamp 1
transform 1 0 75532 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_813
timestamp 1636968456
transform 1 0 75900 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_825
timestamp 1636968456
transform 1 0 77004 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_837
timestamp 1
transform 1 0 78108 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_841
timestamp 1636968456
transform 1 0 78476 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_853
timestamp 1636968456
transform 1 0 79580 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_865
timestamp 1
transform 1 0 80684 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_869
timestamp 1636968456
transform 1 0 81052 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_881
timestamp 1636968456
transform 1 0 82156 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_893
timestamp 1
transform 1 0 83260 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_897
timestamp 1636968456
transform 1 0 83628 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_909
timestamp 1636968456
transform 1 0 84732 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_921
timestamp 1
transform 1 0 85836 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_925
timestamp 1636968456
transform 1 0 86204 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_937
timestamp 1636968456
transform 1 0 87308 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_949
timestamp 1
transform 1 0 88412 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_953
timestamp 1636968456
transform 1 0 88780 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_965
timestamp 1636968456
transform 1 0 89884 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_977
timestamp 1
transform 1 0 90988 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_981
timestamp 1636968456
transform 1 0 91356 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_993
timestamp 1636968456
transform 1 0 92460 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1005
timestamp 1
transform 1 0 93564 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1009
timestamp 1636968456
transform 1 0 93932 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1021
timestamp 1636968456
transform 1 0 95036 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1033
timestamp 1
transform 1 0 96140 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1037
timestamp 1636968456
transform 1 0 96508 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1049
timestamp 1636968456
transform 1 0 97612 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1061
timestamp 1
transform 1 0 98716 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1065
timestamp 1636968456
transform 1 0 99084 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1077
timestamp 1636968456
transform 1 0 100188 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1089
timestamp 1
transform 1 0 101292 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1093
timestamp 1636968456
transform 1 0 101660 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1105
timestamp 1636968456
transform 1 0 102764 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1117
timestamp 1
transform 1 0 103868 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1121
timestamp 1636968456
transform 1 0 104236 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1133
timestamp 1636968456
transform 1 0 105340 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1145
timestamp 1
transform 1 0 106444 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1149
timestamp 1636968456
transform 1 0 106812 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_266_1161
timestamp 1
transform 1 0 107916 0 1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_266_1167
timestamp 1
transform 1 0 108468 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1
transform -1 0 2300 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1
transform 1 0 1380 0 -1 89216
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1
transform 1 0 1380 0 1 80512
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1
transform -1 0 1656 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1
transform -1 0 1656 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1
transform -1 0 1656 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1
transform -1 0 1656 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1
transform -1 0 1656 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1
transform -1 0 1656 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1
transform -1 0 1656 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1
transform 1 0 37444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1
transform 1 0 38732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1
transform 1 0 40020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1
transform 1 0 41308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1
transform -1 0 42228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1
transform 1 0 31648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1
transform 1 0 34224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1
transform 1 0 1380 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1
transform 1 0 1380 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1
transform 1 0 1380 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1
transform 1 0 1380 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1
transform 1 0 1380 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1
transform 1 0 1380 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1
transform 1 0 1380 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1
transform 1 0 1380 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1
transform 1 0 1380 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1
transform 1 0 1380 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1
transform 1 0 1380 0 -1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1
transform 1 0 1380 0 1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1
transform 1 0 1380 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1
transform 1 0 1380 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1
transform 1 0 1380 0 1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1
transform 1 0 1380 0 -1 88128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1
transform 1 0 108284 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew85
timestamp 1
transform 1 0 91816 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  load_slew86
timestamp 1
transform 1 0 89240 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  load_slew87
timestamp 1
transform 1 0 90620 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew88
timestamp 1
transform 1 0 91356 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew89
timestamp 1
transform -1 0 90988 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew90
timestamp 1
transform -1 0 90620 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  load_slew91
timestamp 1
transform 1 0 89608 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew92
timestamp 1
transform 1 0 90988 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew93
timestamp 1
transform -1 0 88872 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  load_slew94
timestamp 1
transform 1 0 89608 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew95
timestamp 1
transform 1 0 89976 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew96
timestamp 1
transform -1 0 89976 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew97
timestamp 1
transform 1 0 89332 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  load_slew98
timestamp 1
transform 1 0 92368 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  load_slew99
timestamp 1
transform 1 0 92368 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  load_slew100
timestamp 1
transform 1 0 90712 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  load_slew101
timestamp 1
transform 1 0 91816 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew102
timestamp 1
transform 1 0 90712 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew103
timestamp 1
transform -1 0 86572 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  load_slew104
timestamp 1
transform -1 0 86664 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  load_slew105
timestamp 1
transform 1 0 86848 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  load_slew106
timestamp 1
transform 1 0 85928 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew107
timestamp 1
transform -1 0 84364 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew108
timestamp 1
transform 1 0 90528 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew109
timestamp 1
transform -1 0 90620 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew110
timestamp 1
transform -1 0 84088 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mem_i0_114
timestamp 1
transform -1 0 104604 0 1 59840
box -38 -48 314 592
use ram_256x16  mem_i0
timestamp 0
transform 1 0 10000 0 1 10000
box 0 0 1 1
use sky130_fd_sc_hd__conb_1  mem_i1_115
timestamp 1
transform -1 0 104604 0 1 129472
box -38 -48 314 592
use ram_256x16  mem_i1
timestamp 0
transform 1 0 10000 0 1 80000
box 0 0 1 1
use sky130_fd_sc_hd__clkbuf_1  output52
timestamp 1
transform 1 0 1380 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output53
timestamp 1
transform -1 0 108560 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output54
timestamp 1
transform -1 0 108560 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output55
timestamp 1
transform -1 0 108560 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output56
timestamp 1
transform -1 0 108560 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output57
timestamp 1
transform -1 0 108560 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output58
timestamp 1
transform -1 0 108560 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output59
timestamp 1
transform 1 0 1380 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output60
timestamp 1
transform 1 0 1380 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output61
timestamp 1
transform 1 0 1380 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output62
timestamp 1
transform 1 0 1380 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output63
timestamp 1
transform 1 0 1380 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output64
timestamp 1
transform -1 0 108560 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output65
timestamp 1
transform -1 0 108560 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output66
timestamp 1
transform -1 0 108560 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output67
timestamp 1
transform -1 0 108560 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_267
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 108836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_268
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 108836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_269
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 108836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_270
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 108836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_271
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 108836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_272
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 108836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_273
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 108836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_274
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 108836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_275
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 108836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_276
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 108836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_533
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_747
timestamp 1
transform -1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_534
timestamp 1
transform 1 0 104052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_53
timestamp 1
transform -1 0 108836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_277
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_641
timestamp 1
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_535
timestamp 1
transform 1 0 104052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_54
timestamp 1
transform -1 0 108836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_278
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_642
timestamp 1
transform -1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_536
timestamp 1
transform 1 0 104052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_55
timestamp 1
transform -1 0 108836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_279
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_643
timestamp 1
transform -1 0 7912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_537
timestamp 1
transform 1 0 104052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_56
timestamp 1
transform -1 0 108836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Left_280
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Right_644
timestamp 1
transform -1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_538
timestamp 1
transform 1 0 104052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_57
timestamp 1
transform -1 0 108836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Left_281
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Right_645
timestamp 1
transform -1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_539
timestamp 1
transform 1 0 104052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_58
timestamp 1
transform -1 0 108836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Left_282
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Right_646
timestamp 1
transform -1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_540
timestamp 1
transform 1 0 104052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_59
timestamp 1
transform -1 0 108836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Left_283
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Right_647
timestamp 1
transform -1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_541
timestamp 1
transform 1 0 104052 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_60
timestamp 1
transform -1 0 108836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Left_284
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Right_648
timestamp 1
transform -1 0 7912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_542
timestamp 1
transform 1 0 104052 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_61
timestamp 1
transform -1 0 108836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Left_285
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Right_649
timestamp 1
transform -1 0 7912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_543
timestamp 1
transform 1 0 104052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_62
timestamp 1
transform -1 0 108836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Left_286
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Right_650
timestamp 1
transform -1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_544
timestamp 1
transform 1 0 104052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_63
timestamp 1
transform -1 0 108836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Left_287
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Right_651
timestamp 1
transform -1 0 7912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_545
timestamp 1
transform 1 0 104052 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_64
timestamp 1
transform -1 0 108836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Left_288
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Right_652
timestamp 1
transform -1 0 7912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_546
timestamp 1
transform 1 0 104052 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_65
timestamp 1
transform -1 0 108836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Left_289
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Right_653
timestamp 1
transform -1 0 7912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_547
timestamp 1
transform 1 0 104052 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_66
timestamp 1
transform -1 0 108836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Left_290
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Right_654
timestamp 1
transform -1 0 7912 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_548
timestamp 1
transform 1 0 104052 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_67
timestamp 1
transform -1 0 108836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Left_291
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Right_655
timestamp 1
transform -1 0 7912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_549
timestamp 1
transform 1 0 104052 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_68
timestamp 1
transform -1 0 108836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Left_292
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Right_656
timestamp 1
transform -1 0 7912 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_550
timestamp 1
transform 1 0 104052 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_69
timestamp 1
transform -1 0 108836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Left_293
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Right_657
timestamp 1
transform -1 0 7912 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_551
timestamp 1
transform 1 0 104052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_70
timestamp 1
transform -1 0 108836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Left_294
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Right_658
timestamp 1
transform -1 0 7912 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_552
timestamp 1
transform 1 0 104052 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_71
timestamp 1
transform -1 0 108836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Left_295
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Right_659
timestamp 1
transform -1 0 7912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_553
timestamp 1
transform 1 0 104052 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_72
timestamp 1
transform -1 0 108836 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Left_296
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Right_660
timestamp 1
transform -1 0 7912 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_554
timestamp 1
transform 1 0 104052 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_73
timestamp 1
transform -1 0 108836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Left_297
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Right_661
timestamp 1
transform -1 0 7912 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_555
timestamp 1
transform 1 0 104052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_74
timestamp 1
transform -1 0 108836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Left_298
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Right_662
timestamp 1
transform -1 0 7912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_556
timestamp 1
transform 1 0 104052 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_75
timestamp 1
transform -1 0 108836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Left_299
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Right_663
timestamp 1
transform -1 0 7912 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_557
timestamp 1
transform 1 0 104052 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_76
timestamp 1
transform -1 0 108836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Left_300
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Right_664
timestamp 1
transform -1 0 7912 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_558
timestamp 1
transform 1 0 104052 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_77
timestamp 1
transform -1 0 108836 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Left_301
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Right_665
timestamp 1
transform -1 0 7912 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_559
timestamp 1
transform 1 0 104052 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_78
timestamp 1
transform -1 0 108836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Left_302
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Right_666
timestamp 1
transform -1 0 7912 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_560
timestamp 1
transform 1 0 104052 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_79
timestamp 1
transform -1 0 108836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Left_303
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Right_667
timestamp 1
transform -1 0 7912 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_561
timestamp 1
transform 1 0 104052 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_80
timestamp 1
transform -1 0 108836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Left_304
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Right_668
timestamp 1
transform -1 0 7912 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_562
timestamp 1
transform 1 0 104052 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_81
timestamp 1
transform -1 0 108836 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Left_305
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Right_669
timestamp 1
transform -1 0 7912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_563
timestamp 1
transform 1 0 104052 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_82
timestamp 1
transform -1 0 108836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Left_306
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Right_670
timestamp 1
transform -1 0 7912 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_564
timestamp 1
transform 1 0 104052 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_83
timestamp 1
transform -1 0 108836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Left_307
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Right_671
timestamp 1
transform -1 0 7912 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_565
timestamp 1
transform 1 0 104052 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_84
timestamp 1
transform -1 0 108836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Left_308
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Right_672
timestamp 1
transform -1 0 7912 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_566
timestamp 1
transform 1 0 104052 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_85
timestamp 1
transform -1 0 108836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Left_309
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Right_673
timestamp 1
transform -1 0 7912 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_567
timestamp 1
transform 1 0 104052 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_86
timestamp 1
transform -1 0 108836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Left_310
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Right_674
timestamp 1
transform -1 0 7912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_568
timestamp 1
transform 1 0 104052 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_87
timestamp 1
transform -1 0 108836 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Left_311
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Right_675
timestamp 1
transform -1 0 7912 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_569
timestamp 1
transform 1 0 104052 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_88
timestamp 1
transform -1 0 108836 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Left_312
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Right_676
timestamp 1
transform -1 0 7912 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_570
timestamp 1
transform 1 0 104052 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_89
timestamp 1
transform -1 0 108836 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Left_313
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Right_677
timestamp 1
transform -1 0 7912 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_571
timestamp 1
transform 1 0 104052 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_90
timestamp 1
transform -1 0 108836 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Left_314
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Right_678
timestamp 1
transform -1 0 7912 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_572
timestamp 1
transform 1 0 104052 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_91
timestamp 1
transform -1 0 108836 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Left_315
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Right_679
timestamp 1
transform -1 0 7912 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_573
timestamp 1
transform 1 0 104052 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_92
timestamp 1
transform -1 0 108836 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Left_316
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Right_680
timestamp 1
transform -1 0 7912 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_574
timestamp 1
transform 1 0 104052 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_93
timestamp 1
transform -1 0 108836 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Left_317
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Right_681
timestamp 1
transform -1 0 7912 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_575
timestamp 1
transform 1 0 104052 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_94
timestamp 1
transform -1 0 108836 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Left_318
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Right_682
timestamp 1
transform -1 0 7912 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_576
timestamp 1
transform 1 0 104052 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_95
timestamp 1
transform -1 0 108836 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Left_319
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Right_683
timestamp 1
transform -1 0 7912 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_577
timestamp 1
transform 1 0 104052 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_96
timestamp 1
transform -1 0 108836 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Left_320
timestamp 1
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Right_684
timestamp 1
transform -1 0 7912 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_578
timestamp 1
transform 1 0 104052 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_97
timestamp 1
transform -1 0 108836 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Left_321
timestamp 1
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Right_685
timestamp 1
transform -1 0 7912 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_579
timestamp 1
transform 1 0 104052 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_98
timestamp 1
transform -1 0 108836 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Left_322
timestamp 1
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Right_686
timestamp 1
transform -1 0 7912 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_580
timestamp 1
transform 1 0 104052 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_99
timestamp 1
transform -1 0 108836 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Left_323
timestamp 1
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Right_687
timestamp 1
transform -1 0 7912 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_581
timestamp 1
transform 1 0 104052 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_100
timestamp 1
transform -1 0 108836 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Left_324
timestamp 1
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Right_688
timestamp 1
transform -1 0 7912 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_582
timestamp 1
transform 1 0 104052 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_101
timestamp 1
transform -1 0 108836 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Left_325
timestamp 1
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Right_689
timestamp 1
transform -1 0 7912 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_583
timestamp 1
transform 1 0 104052 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_102
timestamp 1
transform -1 0 108836 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Left_326
timestamp 1
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Right_690
timestamp 1
transform -1 0 7912 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_584
timestamp 1
transform 1 0 104052 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_103
timestamp 1
transform -1 0 108836 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Left_327
timestamp 1
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Right_691
timestamp 1
transform -1 0 7912 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_585
timestamp 1
transform 1 0 104052 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_104
timestamp 1
transform -1 0 108836 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Left_328
timestamp 1
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Right_692
timestamp 1
transform -1 0 7912 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_586
timestamp 1
transform 1 0 104052 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_105
timestamp 1
transform -1 0 108836 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Left_329
timestamp 1
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Right_693
timestamp 1
transform -1 0 7912 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_587
timestamp 1
transform 1 0 104052 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_106
timestamp 1
transform -1 0 108836 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Left_330
timestamp 1
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Right_694
timestamp 1
transform -1 0 7912 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_588
timestamp 1
transform 1 0 104052 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_107
timestamp 1
transform -1 0 108836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Left_331
timestamp 1
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Right_695
timestamp 1
transform -1 0 7912 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_589
timestamp 1
transform 1 0 104052 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_108
timestamp 1
transform -1 0 108836 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Left_332
timestamp 1
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Right_696
timestamp 1
transform -1 0 7912 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_590
timestamp 1
transform 1 0 104052 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_109
timestamp 1
transform -1 0 108836 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Left_333
timestamp 1
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Right_697
timestamp 1
transform -1 0 7912 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Left_591
timestamp 1
transform 1 0 104052 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Right_110
timestamp 1
transform -1 0 108836 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Left_334
timestamp 1
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Right_698
timestamp 1
transform -1 0 7912 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Left_592
timestamp 1
transform 1 0 104052 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Right_111
timestamp 1
transform -1 0 108836 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Left_335
timestamp 1
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Right_699
timestamp 1
transform -1 0 7912 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Left_593
timestamp 1
transform 1 0 104052 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Right_112
timestamp 1
transform -1 0 108836 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Left_336
timestamp 1
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Right_700
timestamp 1
transform -1 0 7912 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Left_594
timestamp 1
transform 1 0 104052 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Right_113
timestamp 1
transform -1 0 108836 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Left_337
timestamp 1
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Right_701
timestamp 1
transform -1 0 7912 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Left_595
timestamp 1
transform 1 0 104052 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Right_114
timestamp 1
transform -1 0 108836 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Left_338
timestamp 1
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Right_702
timestamp 1
transform -1 0 7912 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Left_596
timestamp 1
transform 1 0 104052 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Right_115
timestamp 1
transform -1 0 108836 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Left_339
timestamp 1
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Right_703
timestamp 1
transform -1 0 7912 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Left_597
timestamp 1
transform 1 0 104052 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Right_116
timestamp 1
transform -1 0 108836 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Left_340
timestamp 1
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Right_704
timestamp 1
transform -1 0 7912 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Left_598
timestamp 1
transform 1 0 104052 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Right_117
timestamp 1
transform -1 0 108836 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Left_341
timestamp 1
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Right_705
timestamp 1
transform -1 0 7912 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Left_599
timestamp 1
transform 1 0 104052 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Right_118
timestamp 1
transform -1 0 108836 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Left_342
timestamp 1
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Right_706
timestamp 1
transform -1 0 7912 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Left_600
timestamp 1
transform 1 0 104052 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Right_119
timestamp 1
transform -1 0 108836 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Left_343
timestamp 1
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Right_707
timestamp 1
transform -1 0 7912 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Left_601
timestamp 1
transform 1 0 104052 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Right_120
timestamp 1
transform -1 0 108836 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Left_344
timestamp 1
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Right_708
timestamp 1
transform -1 0 7912 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Left_602
timestamp 1
transform 1 0 104052 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Right_121
timestamp 1
transform -1 0 108836 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Left_345
timestamp 1
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Right_709
timestamp 1
transform -1 0 7912 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Left_603
timestamp 1
transform 1 0 104052 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Right_122
timestamp 1
transform -1 0 108836 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Left_346
timestamp 1
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Right_710
timestamp 1
transform -1 0 7912 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Left_604
timestamp 1
transform 1 0 104052 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Right_123
timestamp 1
transform -1 0 108836 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Left_347
timestamp 1
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Right_711
timestamp 1
transform -1 0 7912 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Left_605
timestamp 1
transform 1 0 104052 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Right_124
timestamp 1
transform -1 0 108836 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Left_348
timestamp 1
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Right_712
timestamp 1
transform -1 0 7912 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Left_606
timestamp 1
transform 1 0 104052 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Right_125
timestamp 1
transform -1 0 108836 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Left_349
timestamp 1
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Right_713
timestamp 1
transform -1 0 7912 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Left_607
timestamp 1
transform 1 0 104052 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Right_126
timestamp 1
transform -1 0 108836 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Left_350
timestamp 1
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Right_714
timestamp 1
transform -1 0 7912 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Left_608
timestamp 1
transform 1 0 104052 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Right_127
timestamp 1
transform -1 0 108836 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Left_351
timestamp 1
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Right_715
timestamp 1
transform -1 0 7912 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Left_609
timestamp 1
transform 1 0 104052 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Right_128
timestamp 1
transform -1 0 108836 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Left_352
timestamp 1
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Right_716
timestamp 1
transform -1 0 7912 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Left_610
timestamp 1
transform 1 0 104052 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Right_129
timestamp 1
transform -1 0 108836 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Left_353
timestamp 1
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Right_717
timestamp 1
transform -1 0 7912 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Left_611
timestamp 1
transform 1 0 104052 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Right_130
timestamp 1
transform -1 0 108836 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Left_354
timestamp 1
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Right_718
timestamp 1
transform -1 0 7912 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Left_612
timestamp 1
transform 1 0 104052 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Right_131
timestamp 1
transform -1 0 108836 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Left_355
timestamp 1
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Right_719
timestamp 1
transform -1 0 7912 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Left_613
timestamp 1
transform 1 0 104052 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Right_132
timestamp 1
transform -1 0 108836 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Left_356
timestamp 1
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Right_720
timestamp 1
transform -1 0 7912 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Left_614
timestamp 1
transform 1 0 104052 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Right_133
timestamp 1
transform -1 0 108836 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Left_357
timestamp 1
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Right_721
timestamp 1
transform -1 0 7912 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Left_615
timestamp 1
transform 1 0 104052 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Right_134
timestamp 1
transform -1 0 108836 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Left_358
timestamp 1
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Right_722
timestamp 1
transform -1 0 7912 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Left_616
timestamp 1
transform 1 0 104052 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Right_135
timestamp 1
transform -1 0 108836 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Left_359
timestamp 1
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Right_723
timestamp 1
transform -1 0 7912 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Left_617
timestamp 1
transform 1 0 104052 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Right_136
timestamp 1
transform -1 0 108836 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Left_360
timestamp 1
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Right_724
timestamp 1
transform -1 0 7912 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Left_618
timestamp 1
transform 1 0 104052 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Right_137
timestamp 1
transform -1 0 108836 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Left_361
timestamp 1
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Right_725
timestamp 1
transform -1 0 7912 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Left_619
timestamp 1
transform 1 0 104052 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Right_138
timestamp 1
transform -1 0 108836 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Left_362
timestamp 1
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Right_726
timestamp 1
transform -1 0 7912 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Left_620
timestamp 1
transform 1 0 104052 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Right_139
timestamp 1
transform -1 0 108836 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Left_363
timestamp 1
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Right_727
timestamp 1
transform -1 0 7912 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Left_621
timestamp 1
transform 1 0 104052 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Right_140
timestamp 1
transform -1 0 108836 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Left_364
timestamp 1
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Right_728
timestamp 1
transform -1 0 7912 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Left_622
timestamp 1
transform 1 0 104052 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Right_141
timestamp 1
transform -1 0 108836 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Left_365
timestamp 1
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Right_729
timestamp 1
transform -1 0 7912 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Left_623
timestamp 1
transform 1 0 104052 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Right_142
timestamp 1
transform -1 0 108836 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Left_366
timestamp 1
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Right_730
timestamp 1
transform -1 0 7912 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Left_624
timestamp 1
transform 1 0 104052 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Right_143
timestamp 1
transform -1 0 108836 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Left_367
timestamp 1
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Right_731
timestamp 1
transform -1 0 7912 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Left_625
timestamp 1
transform 1 0 104052 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Right_144
timestamp 1
transform -1 0 108836 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Left_368
timestamp 1
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Right_732
timestamp 1
transform -1 0 7912 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Left_626
timestamp 1
transform 1 0 104052 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Right_145
timestamp 1
transform -1 0 108836 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Left_369
timestamp 1
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Right_733
timestamp 1
transform -1 0 7912 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Left_627
timestamp 1
transform 1 0 104052 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Right_146
timestamp 1
transform -1 0 108836 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Left_370
timestamp 1
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Right_734
timestamp 1
transform -1 0 7912 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Left_628
timestamp 1
transform 1 0 104052 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Right_147
timestamp 1
transform -1 0 108836 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Left_371
timestamp 1
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Right_735
timestamp 1
transform -1 0 7912 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Left_629
timestamp 1
transform 1 0 104052 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Right_148
timestamp 1
transform -1 0 108836 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Left_372
timestamp 1
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Right_736
timestamp 1
transform -1 0 7912 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Left_630
timestamp 1
transform 1 0 104052 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Right_149
timestamp 1
transform -1 0 108836 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Left_373
timestamp 1
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Right_737
timestamp 1
transform -1 0 7912 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Left_631
timestamp 1
transform 1 0 104052 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Right_150
timestamp 1
transform -1 0 108836 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Left_374
timestamp 1
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Right_738
timestamp 1
transform -1 0 7912 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Left_632
timestamp 1
transform 1 0 104052 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Right_151
timestamp 1
transform -1 0 108836 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Left_375
timestamp 1
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Right_739
timestamp 1
transform -1 0 7912 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Left_633
timestamp 1
transform 1 0 104052 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Right_152
timestamp 1
transform -1 0 108836 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Left_376
timestamp 1
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Right_740
timestamp 1
transform -1 0 7912 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Left_634
timestamp 1
transform 1 0 104052 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Right_153
timestamp 1
transform -1 0 108836 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Left_377
timestamp 1
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Right_741
timestamp 1
transform -1 0 7912 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Left_635
timestamp 1
transform 1 0 104052 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Right_154
timestamp 1
transform -1 0 108836 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Left_378
timestamp 1
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Right_742
timestamp 1
transform -1 0 7912 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Left_636
timestamp 1
transform 1 0 104052 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Right_155
timestamp 1
transform -1 0 108836 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Left_379
timestamp 1
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Right_743
timestamp 1
transform -1 0 7912 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Left_637
timestamp 1
transform 1 0 104052 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Right_156
timestamp 1
transform -1 0 108836 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Left_380
timestamp 1
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Right_744
timestamp 1
transform -1 0 7912 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Left_638
timestamp 1
transform 1 0 104052 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Right_157
timestamp 1
transform -1 0 108836 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Left_381
timestamp 1
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Right_745
timestamp 1
transform -1 0 7912 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Left_639
timestamp 1
transform 1 0 104052 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Right_158
timestamp 1
transform -1 0 108836 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Left_382
timestamp 1
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Right_746
timestamp 1
transform -1 0 7912 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Left_640
timestamp 1
transform 1 0 104052 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Right_159
timestamp 1
transform -1 0 108836 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Left_384
timestamp 1
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Right_10
timestamp 1
transform -1 0 108836 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Left_385
timestamp 1
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Right_11
timestamp 1
transform -1 0 108836 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Left_386
timestamp 1
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Right_12
timestamp 1
transform -1 0 108836 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Left_387
timestamp 1
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Right_13
timestamp 1
transform -1 0 108836 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Left_388
timestamp 1
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Right_14
timestamp 1
transform -1 0 108836 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Left_389
timestamp 1
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Right_15
timestamp 1
transform -1 0 108836 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Left_390
timestamp 1
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Right_16
timestamp 1
transform -1 0 108836 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Left_391
timestamp 1
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Right_17
timestamp 1
transform -1 0 108836 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Left_392
timestamp 1
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Right_18
timestamp 1
transform -1 0 108836 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Left_393
timestamp 1
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Right_19
timestamp 1
transform -1 0 108836 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Left_394
timestamp 1
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Right_20
timestamp 1
transform -1 0 108836 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Left_395
timestamp 1
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Right_21
timestamp 1
transform -1 0 108836 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Left_396
timestamp 1
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Right_22
timestamp 1
transform -1 0 108836 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Left_397
timestamp 1
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Right_23
timestamp 1
transform -1 0 108836 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_Left_398
timestamp 1
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_Right_24
timestamp 1
transform -1 0 108836 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_Left_399
timestamp 1
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_Right_25
timestamp 1
transform -1 0 108836 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_Left_400
timestamp 1
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_Right_26
timestamp 1
transform -1 0 108836 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_Left_401
timestamp 1
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_Right_27
timestamp 1
transform -1 0 108836 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_Left_402
timestamp 1
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_Right_28
timestamp 1
transform -1 0 108836 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_Left_403
timestamp 1
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_Right_29
timestamp 1
transform -1 0 108836 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_Left_404
timestamp 1
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_Right_30
timestamp 1
transform -1 0 108836 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_Left_405
timestamp 1
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_Right_31
timestamp 1
transform -1 0 108836 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Left_383
timestamp 1
transform 1 0 1104 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Right_855
timestamp 1
transform -1 0 7912 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Left_748
timestamp 1
transform 1 0 104052 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Right_160
timestamp 1
transform -1 0 108836 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Left_406
timestamp 1
transform 1 0 1104 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Right_856
timestamp 1
transform -1 0 7912 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Left_749
timestamp 1
transform 1 0 104052 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Right_161
timestamp 1
transform -1 0 108836 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Left_407
timestamp 1
transform 1 0 1104 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Right_857
timestamp 1
transform -1 0 7912 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Left_750
timestamp 1
transform 1 0 104052 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Right_162
timestamp 1
transform -1 0 108836 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Left_408
timestamp 1
transform 1 0 1104 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Right_858
timestamp 1
transform -1 0 7912 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Left_751
timestamp 1
transform 1 0 104052 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Right_163
timestamp 1
transform -1 0 108836 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Left_409
timestamp 1
transform 1 0 1104 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Right_859
timestamp 1
transform -1 0 7912 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Left_752
timestamp 1
transform 1 0 104052 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Right_164
timestamp 1
transform -1 0 108836 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Left_410
timestamp 1
transform 1 0 1104 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Right_860
timestamp 1
transform -1 0 7912 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Left_753
timestamp 1
transform 1 0 104052 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Right_165
timestamp 1
transform -1 0 108836 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Left_411
timestamp 1
transform 1 0 1104 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Right_861
timestamp 1
transform -1 0 7912 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Left_754
timestamp 1
transform 1 0 104052 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Right_166
timestamp 1
transform -1 0 108836 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Left_412
timestamp 1
transform 1 0 1104 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Right_862
timestamp 1
transform -1 0 7912 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Left_755
timestamp 1
transform 1 0 104052 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Right_167
timestamp 1
transform -1 0 108836 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Left_413
timestamp 1
transform 1 0 1104 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Right_863
timestamp 1
transform -1 0 7912 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Left_756
timestamp 1
transform 1 0 104052 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Right_168
timestamp 1
transform -1 0 108836 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Left_414
timestamp 1
transform 1 0 1104 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Right_864
timestamp 1
transform -1 0 7912 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Left_757
timestamp 1
transform 1 0 104052 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Right_169
timestamp 1
transform -1 0 108836 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Left_415
timestamp 1
transform 1 0 1104 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Right_865
timestamp 1
transform -1 0 7912 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Left_758
timestamp 1
transform 1 0 104052 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Right_170
timestamp 1
transform -1 0 108836 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Left_416
timestamp 1
transform 1 0 1104 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Right_866
timestamp 1
transform -1 0 7912 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Left_759
timestamp 1
transform 1 0 104052 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Right_171
timestamp 1
transform -1 0 108836 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Left_417
timestamp 1
transform 1 0 1104 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Right_867
timestamp 1
transform -1 0 7912 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Left_760
timestamp 1
transform 1 0 104052 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Right_172
timestamp 1
transform -1 0 108836 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Left_418
timestamp 1
transform 1 0 1104 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Right_868
timestamp 1
transform -1 0 7912 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Left_761
timestamp 1
transform 1 0 104052 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Right_173
timestamp 1
transform -1 0 108836 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Left_419
timestamp 1
transform 1 0 1104 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Right_869
timestamp 1
transform -1 0 7912 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Left_762
timestamp 1
transform 1 0 104052 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Right_174
timestamp 1
transform -1 0 108836 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Left_420
timestamp 1
transform 1 0 1104 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Right_870
timestamp 1
transform -1 0 7912 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Left_763
timestamp 1
transform 1 0 104052 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Right_175
timestamp 1
transform -1 0 108836 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Left_421
timestamp 1
transform 1 0 1104 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Right_871
timestamp 1
transform -1 0 7912 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Left_764
timestamp 1
transform 1 0 104052 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Right_176
timestamp 1
transform -1 0 108836 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Left_422
timestamp 1
transform 1 0 1104 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Right_872
timestamp 1
transform -1 0 7912 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_2_Left_765
timestamp 1
transform 1 0 104052 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_2_Right_177
timestamp 1
transform -1 0 108836 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Left_423
timestamp 1
transform 1 0 1104 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Right_873
timestamp 1
transform -1 0 7912 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_2_Left_766
timestamp 1
transform 1 0 104052 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_2_Right_178
timestamp 1
transform -1 0 108836 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Left_424
timestamp 1
transform 1 0 1104 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Right_874
timestamp 1
transform -1 0 7912 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_2_Left_767
timestamp 1
transform 1 0 104052 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_2_Right_179
timestamp 1
transform -1 0 108836 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Left_425
timestamp 1
transform 1 0 1104 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Right_875
timestamp 1
transform -1 0 7912 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_2_Left_768
timestamp 1
transform 1 0 104052 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_2_Right_180
timestamp 1
transform -1 0 108836 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Left_426
timestamp 1
transform 1 0 1104 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Right_876
timestamp 1
transform -1 0 7912 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_2_Left_769
timestamp 1
transform 1 0 104052 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_2_Right_181
timestamp 1
transform -1 0 108836 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Left_427
timestamp 1
transform 1 0 1104 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Right_877
timestamp 1
transform -1 0 7912 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_2_Left_770
timestamp 1
transform 1 0 104052 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_2_Right_182
timestamp 1
transform -1 0 108836 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Left_428
timestamp 1
transform 1 0 1104 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Right_878
timestamp 1
transform -1 0 7912 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_2_Left_771
timestamp 1
transform 1 0 104052 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_2_Right_183
timestamp 1
transform -1 0 108836 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Left_429
timestamp 1
transform 1 0 1104 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Right_879
timestamp 1
transform -1 0 7912 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_2_Left_772
timestamp 1
transform 1 0 104052 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_2_Right_184
timestamp 1
transform -1 0 108836 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_1_Left_430
timestamp 1
transform 1 0 1104 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_1_Right_880
timestamp 1
transform -1 0 7912 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_2_Left_773
timestamp 1
transform 1 0 104052 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_2_Right_185
timestamp 1
transform -1 0 108836 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_1_Left_431
timestamp 1
transform 1 0 1104 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_1_Right_881
timestamp 1
transform -1 0 7912 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_2_Left_774
timestamp 1
transform 1 0 104052 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_2_Right_186
timestamp 1
transform -1 0 108836 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_1_Left_432
timestamp 1
transform 1 0 1104 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_1_Right_882
timestamp 1
transform -1 0 7912 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_2_Left_775
timestamp 1
transform 1 0 104052 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_2_Right_187
timestamp 1
transform -1 0 108836 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_1_Left_433
timestamp 1
transform 1 0 1104 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_1_Right_883
timestamp 1
transform -1 0 7912 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_2_Left_776
timestamp 1
transform 1 0 104052 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_2_Right_188
timestamp 1
transform -1 0 108836 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_1_Left_434
timestamp 1
transform 1 0 1104 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_1_Right_884
timestamp 1
transform -1 0 7912 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_2_Left_777
timestamp 1
transform 1 0 104052 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_2_Right_189
timestamp 1
transform -1 0 108836 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_1_Left_435
timestamp 1
transform 1 0 1104 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_1_Right_885
timestamp 1
transform -1 0 7912 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_2_Left_778
timestamp 1
transform 1 0 104052 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_2_Right_190
timestamp 1
transform -1 0 108836 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_1_Left_436
timestamp 1
transform 1 0 1104 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_1_Right_886
timestamp 1
transform -1 0 7912 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_2_Left_779
timestamp 1
transform 1 0 104052 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_2_Right_191
timestamp 1
transform -1 0 108836 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_1_Left_437
timestamp 1
transform 1 0 1104 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_1_Right_887
timestamp 1
transform -1 0 7912 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_2_Left_780
timestamp 1
transform 1 0 104052 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_2_Right_192
timestamp 1
transform -1 0 108836 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_1_Left_438
timestamp 1
transform 1 0 1104 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_1_Right_888
timestamp 1
transform -1 0 7912 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_2_Left_781
timestamp 1
transform 1 0 104052 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_2_Right_193
timestamp 1
transform -1 0 108836 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_1_Left_439
timestamp 1
transform 1 0 1104 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_1_Right_889
timestamp 1
transform -1 0 7912 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_2_Left_782
timestamp 1
transform 1 0 104052 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_2_Right_194
timestamp 1
transform -1 0 108836 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_1_Left_440
timestamp 1
transform 1 0 1104 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_1_Right_890
timestamp 1
transform -1 0 7912 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_2_Left_783
timestamp 1
transform 1 0 104052 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_2_Right_195
timestamp 1
transform -1 0 108836 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_1_Left_441
timestamp 1
transform 1 0 1104 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_1_Right_891
timestamp 1
transform -1 0 7912 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_2_Left_784
timestamp 1
transform 1 0 104052 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_2_Right_196
timestamp 1
transform -1 0 108836 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_1_Left_442
timestamp 1
transform 1 0 1104 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_1_Right_892
timestamp 1
transform -1 0 7912 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_2_Left_785
timestamp 1
transform 1 0 104052 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_2_Right_197
timestamp 1
transform -1 0 108836 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_1_Left_443
timestamp 1
transform 1 0 1104 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_1_Right_893
timestamp 1
transform -1 0 7912 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_2_Left_786
timestamp 1
transform 1 0 104052 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_2_Right_198
timestamp 1
transform -1 0 108836 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_1_Left_444
timestamp 1
transform 1 0 1104 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_1_Right_894
timestamp 1
transform -1 0 7912 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_2_Left_787
timestamp 1
transform 1 0 104052 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_2_Right_199
timestamp 1
transform -1 0 108836 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_1_Left_445
timestamp 1
transform 1 0 1104 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_1_Right_895
timestamp 1
transform -1 0 7912 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_2_Left_788
timestamp 1
transform 1 0 104052 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_2_Right_200
timestamp 1
transform -1 0 108836 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_1_Left_446
timestamp 1
transform 1 0 1104 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_1_Right_896
timestamp 1
transform -1 0 7912 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_2_Left_789
timestamp 1
transform 1 0 104052 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_2_Right_201
timestamp 1
transform -1 0 108836 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_1_Left_447
timestamp 1
transform 1 0 1104 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_1_Right_897
timestamp 1
transform -1 0 7912 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_2_Left_790
timestamp 1
transform 1 0 104052 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_2_Right_202
timestamp 1
transform -1 0 108836 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_1_Left_448
timestamp 1
transform 1 0 1104 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_1_Right_898
timestamp 1
transform -1 0 7912 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_2_Left_791
timestamp 1
transform 1 0 104052 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_2_Right_203
timestamp 1
transform -1 0 108836 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_1_Left_449
timestamp 1
transform 1 0 1104 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_1_Right_899
timestamp 1
transform -1 0 7912 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_2_Left_792
timestamp 1
transform 1 0 104052 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_2_Right_204
timestamp 1
transform -1 0 108836 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_1_Left_450
timestamp 1
transform 1 0 1104 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_1_Right_900
timestamp 1
transform -1 0 7912 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_2_Left_793
timestamp 1
transform 1 0 104052 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_2_Right_205
timestamp 1
transform -1 0 108836 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_1_Left_451
timestamp 1
transform 1 0 1104 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_1_Right_901
timestamp 1
transform -1 0 7912 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_2_Left_794
timestamp 1
transform 1 0 104052 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_2_Right_206
timestamp 1
transform -1 0 108836 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_1_Left_452
timestamp 1
transform 1 0 1104 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_1_Right_902
timestamp 1
transform -1 0 7912 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_2_Left_795
timestamp 1
transform 1 0 104052 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_2_Right_207
timestamp 1
transform -1 0 108836 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_1_Left_453
timestamp 1
transform 1 0 1104 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_1_Right_903
timestamp 1
transform -1 0 7912 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_2_Left_796
timestamp 1
transform 1 0 104052 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_2_Right_208
timestamp 1
transform -1 0 108836 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_1_Left_454
timestamp 1
transform 1 0 1104 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_1_Right_904
timestamp 1
transform -1 0 7912 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_2_Left_797
timestamp 1
transform 1 0 104052 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_2_Right_209
timestamp 1
transform -1 0 108836 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_1_Left_455
timestamp 1
transform 1 0 1104 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_1_Right_905
timestamp 1
transform -1 0 7912 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_2_Left_798
timestamp 1
transform 1 0 104052 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_2_Right_210
timestamp 1
transform -1 0 108836 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_1_Left_456
timestamp 1
transform 1 0 1104 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_1_Right_906
timestamp 1
transform -1 0 7912 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_2_Left_799
timestamp 1
transform 1 0 104052 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_2_Right_211
timestamp 1
transform -1 0 108836 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_1_Left_457
timestamp 1
transform 1 0 1104 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_1_Right_907
timestamp 1
transform -1 0 7912 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_2_Left_800
timestamp 1
transform 1 0 104052 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_2_Right_212
timestamp 1
transform -1 0 108836 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_1_Left_458
timestamp 1
transform 1 0 1104 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_1_Right_908
timestamp 1
transform -1 0 7912 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_2_Left_801
timestamp 1
transform 1 0 104052 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_2_Right_213
timestamp 1
transform -1 0 108836 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_1_Left_459
timestamp 1
transform 1 0 1104 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_1_Right_909
timestamp 1
transform -1 0 7912 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_2_Left_802
timestamp 1
transform 1 0 104052 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_2_Right_214
timestamp 1
transform -1 0 108836 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_1_Left_460
timestamp 1
transform 1 0 1104 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_1_Right_910
timestamp 1
transform -1 0 7912 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_2_Left_803
timestamp 1
transform 1 0 104052 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_2_Right_215
timestamp 1
transform -1 0 108836 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_1_Left_461
timestamp 1
transform 1 0 1104 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_1_Right_911
timestamp 1
transform -1 0 7912 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_2_Left_804
timestamp 1
transform 1 0 104052 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_2_Right_216
timestamp 1
transform -1 0 108836 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_1_Left_462
timestamp 1
transform 1 0 1104 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_1_Right_912
timestamp 1
transform -1 0 7912 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_2_Left_805
timestamp 1
transform 1 0 104052 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_2_Right_217
timestamp 1
transform -1 0 108836 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_1_Left_463
timestamp 1
transform 1 0 1104 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_1_Right_913
timestamp 1
transform -1 0 7912 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_2_Left_806
timestamp 1
transform 1 0 104052 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_2_Right_218
timestamp 1
transform -1 0 108836 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_1_Left_464
timestamp 1
transform 1 0 1104 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_1_Right_914
timestamp 1
transform -1 0 7912 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_2_Left_807
timestamp 1
transform 1 0 104052 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_2_Right_219
timestamp 1
transform -1 0 108836 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_1_Left_465
timestamp 1
transform 1 0 1104 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_1_Right_915
timestamp 1
transform -1 0 7912 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_2_Left_808
timestamp 1
transform 1 0 104052 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_2_Right_220
timestamp 1
transform -1 0 108836 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_1_Left_466
timestamp 1
transform 1 0 1104 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_1_Right_916
timestamp 1
transform -1 0 7912 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_2_Left_809
timestamp 1
transform 1 0 104052 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_2_Right_221
timestamp 1
transform -1 0 108836 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_1_Left_467
timestamp 1
transform 1 0 1104 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_1_Right_917
timestamp 1
transform -1 0 7912 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_2_Left_810
timestamp 1
transform 1 0 104052 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_2_Right_222
timestamp 1
transform -1 0 108836 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_1_Left_468
timestamp 1
transform 1 0 1104 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_1_Right_918
timestamp 1
transform -1 0 7912 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_2_Left_811
timestamp 1
transform 1 0 104052 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_2_Right_223
timestamp 1
transform -1 0 108836 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_1_Left_469
timestamp 1
transform 1 0 1104 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_1_Right_919
timestamp 1
transform -1 0 7912 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_2_Left_812
timestamp 1
transform 1 0 104052 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_2_Right_224
timestamp 1
transform -1 0 108836 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_1_Left_470
timestamp 1
transform 1 0 1104 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_1_Right_920
timestamp 1
transform -1 0 7912 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_2_Left_813
timestamp 1
transform 1 0 104052 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_2_Right_225
timestamp 1
transform -1 0 108836 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_1_Left_471
timestamp 1
transform 1 0 1104 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_1_Right_921
timestamp 1
transform -1 0 7912 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_2_Left_814
timestamp 1
transform 1 0 104052 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_2_Right_226
timestamp 1
transform -1 0 108836 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_1_Left_472
timestamp 1
transform 1 0 1104 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_1_Right_922
timestamp 1
transform -1 0 7912 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_2_Left_815
timestamp 1
transform 1 0 104052 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_2_Right_227
timestamp 1
transform -1 0 108836 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_1_Left_473
timestamp 1
transform 1 0 1104 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_1_Right_923
timestamp 1
transform -1 0 7912 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_2_Left_816
timestamp 1
transform 1 0 104052 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_2_Right_228
timestamp 1
transform -1 0 108836 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_1_Left_474
timestamp 1
transform 1 0 1104 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_1_Right_924
timestamp 1
transform -1 0 7912 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_2_Left_817
timestamp 1
transform 1 0 104052 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_2_Right_229
timestamp 1
transform -1 0 108836 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_1_Left_475
timestamp 1
transform 1 0 1104 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_1_Right_925
timestamp 1
transform -1 0 7912 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_2_Left_818
timestamp 1
transform 1 0 104052 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_2_Right_230
timestamp 1
transform -1 0 108836 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_1_Left_476
timestamp 1
transform 1 0 1104 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_1_Right_926
timestamp 1
transform -1 0 7912 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_2_Left_819
timestamp 1
transform 1 0 104052 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_2_Right_231
timestamp 1
transform -1 0 108836 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_1_Left_477
timestamp 1
transform 1 0 1104 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_1_Right_927
timestamp 1
transform -1 0 7912 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_2_Left_820
timestamp 1
transform 1 0 104052 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_2_Right_232
timestamp 1
transform -1 0 108836 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_1_Left_478
timestamp 1
transform 1 0 1104 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_1_Right_928
timestamp 1
transform -1 0 7912 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_2_Left_821
timestamp 1
transform 1 0 104052 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_2_Right_233
timestamp 1
transform -1 0 108836 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_1_Left_479
timestamp 1
transform 1 0 1104 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_1_Right_929
timestamp 1
transform -1 0 7912 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_2_Left_822
timestamp 1
transform 1 0 104052 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_2_Right_234
timestamp 1
transform -1 0 108836 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_1_Left_480
timestamp 1
transform 1 0 1104 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_1_Right_930
timestamp 1
transform -1 0 7912 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_2_Left_823
timestamp 1
transform 1 0 104052 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_2_Right_235
timestamp 1
transform -1 0 108836 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_1_Left_481
timestamp 1
transform 1 0 1104 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_1_Right_931
timestamp 1
transform -1 0 7912 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_2_Left_824
timestamp 1
transform 1 0 104052 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_2_Right_236
timestamp 1
transform -1 0 108836 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_1_Left_482
timestamp 1
transform 1 0 1104 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_1_Right_932
timestamp 1
transform -1 0 7912 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_2_Left_825
timestamp 1
transform 1 0 104052 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_2_Right_237
timestamp 1
transform -1 0 108836 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_1_Left_483
timestamp 1
transform 1 0 1104 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_1_Right_933
timestamp 1
transform -1 0 7912 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_2_Left_826
timestamp 1
transform 1 0 104052 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_2_Right_238
timestamp 1
transform -1 0 108836 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_1_Left_484
timestamp 1
transform 1 0 1104 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_1_Right_934
timestamp 1
transform -1 0 7912 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_2_Left_827
timestamp 1
transform 1 0 104052 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_2_Right_239
timestamp 1
transform -1 0 108836 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_1_Left_485
timestamp 1
transform 1 0 1104 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_1_Right_935
timestamp 1
transform -1 0 7912 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_2_Left_828
timestamp 1
transform 1 0 104052 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_2_Right_240
timestamp 1
transform -1 0 108836 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_1_Left_486
timestamp 1
transform 1 0 1104 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_1_Right_936
timestamp 1
transform -1 0 7912 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_2_Left_829
timestamp 1
transform 1 0 104052 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_2_Right_241
timestamp 1
transform -1 0 108836 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_1_Left_487
timestamp 1
transform 1 0 1104 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_1_Right_937
timestamp 1
transform -1 0 7912 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_2_Left_830
timestamp 1
transform 1 0 104052 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_2_Right_242
timestamp 1
transform -1 0 108836 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_1_Left_488
timestamp 1
transform 1 0 1104 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_1_Right_938
timestamp 1
transform -1 0 7912 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_2_Left_831
timestamp 1
transform 1 0 104052 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_2_Right_243
timestamp 1
transform -1 0 108836 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_1_Left_489
timestamp 1
transform 1 0 1104 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_1_Right_939
timestamp 1
transform -1 0 7912 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_2_Left_832
timestamp 1
transform 1 0 104052 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_2_Right_244
timestamp 1
transform -1 0 108836 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_1_Left_490
timestamp 1
transform 1 0 1104 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_1_Right_940
timestamp 1
transform -1 0 7912 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_2_Left_833
timestamp 1
transform 1 0 104052 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_2_Right_245
timestamp 1
transform -1 0 108836 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_1_Left_491
timestamp 1
transform 1 0 1104 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_1_Right_941
timestamp 1
transform -1 0 7912 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_2_Left_834
timestamp 1
transform 1 0 104052 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_2_Right_246
timestamp 1
transform -1 0 108836 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_1_Left_492
timestamp 1
transform 1 0 1104 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_1_Right_942
timestamp 1
transform -1 0 7912 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_2_Left_835
timestamp 1
transform 1 0 104052 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_2_Right_247
timestamp 1
transform -1 0 108836 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_1_Left_493
timestamp 1
transform 1 0 1104 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_1_Right_943
timestamp 1
transform -1 0 7912 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_2_Left_836
timestamp 1
transform 1 0 104052 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_2_Right_248
timestamp 1
transform -1 0 108836 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_228_1_Left_494
timestamp 1
transform 1 0 1104 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_228_1_Right_944
timestamp 1
transform -1 0 7912 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_228_2_Left_837
timestamp 1
transform 1 0 104052 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_228_2_Right_249
timestamp 1
transform -1 0 108836 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_229_1_Left_495
timestamp 1
transform 1 0 1104 0 -1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_229_1_Right_945
timestamp 1
transform -1 0 7912 0 -1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_229_2_Left_838
timestamp 1
transform 1 0 104052 0 -1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_229_2_Right_250
timestamp 1
transform -1 0 108836 0 -1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_230_1_Left_496
timestamp 1
transform 1 0 1104 0 1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_230_1_Right_946
timestamp 1
transform -1 0 7912 0 1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_230_2_Left_839
timestamp 1
transform 1 0 104052 0 1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_230_2_Right_251
timestamp 1
transform -1 0 108836 0 1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_231_1_Left_497
timestamp 1
transform 1 0 1104 0 -1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_231_1_Right_947
timestamp 1
transform -1 0 7912 0 -1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_231_2_Left_840
timestamp 1
transform 1 0 104052 0 -1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_231_2_Right_252
timestamp 1
transform -1 0 108836 0 -1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_232_1_Left_498
timestamp 1
transform 1 0 1104 0 1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_232_1_Right_948
timestamp 1
transform -1 0 7912 0 1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_232_2_Left_841
timestamp 1
transform 1 0 104052 0 1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_232_2_Right_253
timestamp 1
transform -1 0 108836 0 1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_233_1_Left_499
timestamp 1
transform 1 0 1104 0 -1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_233_1_Right_949
timestamp 1
transform -1 0 7912 0 -1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_233_2_Left_842
timestamp 1
transform 1 0 104052 0 -1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_233_2_Right_254
timestamp 1
transform -1 0 108836 0 -1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_234_1_Left_500
timestamp 1
transform 1 0 1104 0 1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_234_1_Right_950
timestamp 1
transform -1 0 7912 0 1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_234_2_Left_843
timestamp 1
transform 1 0 104052 0 1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_234_2_Right_255
timestamp 1
transform -1 0 108836 0 1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_235_1_Left_501
timestamp 1
transform 1 0 1104 0 -1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_235_1_Right_951
timestamp 1
transform -1 0 7912 0 -1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_235_2_Left_844
timestamp 1
transform 1 0 104052 0 -1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_235_2_Right_256
timestamp 1
transform -1 0 108836 0 -1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_236_1_Left_502
timestamp 1
transform 1 0 1104 0 1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_236_1_Right_952
timestamp 1
transform -1 0 7912 0 1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_236_2_Left_845
timestamp 1
transform 1 0 104052 0 1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_236_2_Right_257
timestamp 1
transform -1 0 108836 0 1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_237_1_Left_503
timestamp 1
transform 1 0 1104 0 -1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_237_1_Right_953
timestamp 1
transform -1 0 7912 0 -1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_237_2_Left_846
timestamp 1
transform 1 0 104052 0 -1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_237_2_Right_258
timestamp 1
transform -1 0 108836 0 -1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_238_1_Left_504
timestamp 1
transform 1 0 1104 0 1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_238_1_Right_954
timestamp 1
transform -1 0 7912 0 1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_238_2_Left_847
timestamp 1
transform 1 0 104052 0 1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_238_2_Right_259
timestamp 1
transform -1 0 108836 0 1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_239_1_Left_505
timestamp 1
transform 1 0 1104 0 -1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_239_1_Right_955
timestamp 1
transform -1 0 7912 0 -1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_239_2_Left_848
timestamp 1
transform 1 0 104052 0 -1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_239_2_Right_260
timestamp 1
transform -1 0 108836 0 -1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_240_1_Left_506
timestamp 1
transform 1 0 1104 0 1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_240_1_Right_956
timestamp 1
transform -1 0 7912 0 1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_240_2_Left_849
timestamp 1
transform 1 0 104052 0 1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_240_2_Right_261
timestamp 1
transform -1 0 108836 0 1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_241_1_Left_507
timestamp 1
transform 1 0 1104 0 -1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_241_1_Right_957
timestamp 1
transform -1 0 7912 0 -1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_241_2_Left_850
timestamp 1
transform 1 0 104052 0 -1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_241_2_Right_262
timestamp 1
transform -1 0 108836 0 -1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_242_1_Left_508
timestamp 1
transform 1 0 1104 0 1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_242_1_Right_958
timestamp 1
transform -1 0 7912 0 1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_242_2_Left_851
timestamp 1
transform 1 0 104052 0 1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_242_2_Right_263
timestamp 1
transform -1 0 108836 0 1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_243_1_Left_509
timestamp 1
transform 1 0 1104 0 -1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_243_1_Right_959
timestamp 1
transform -1 0 7912 0 -1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_243_2_Left_852
timestamp 1
transform 1 0 104052 0 -1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_243_2_Right_264
timestamp 1
transform -1 0 108836 0 -1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_244_1_Left_510
timestamp 1
transform 1 0 1104 0 1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_244_1_Right_960
timestamp 1
transform -1 0 7912 0 1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_244_2_Left_853
timestamp 1
transform 1 0 104052 0 1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_244_2_Right_265
timestamp 1
transform -1 0 108836 0 1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_245_1_Left_511
timestamp 1
transform 1 0 1104 0 -1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_245_1_Right_961
timestamp 1
transform -1 0 7912 0 -1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_245_2_Left_854
timestamp 1
transform 1 0 104052 0 -1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_245_2_Right_266
timestamp 1
transform -1 0 108836 0 -1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_246_Left_512
timestamp 1
transform 1 0 1104 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_246_Right_32
timestamp 1
transform -1 0 108836 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_247_Left_513
timestamp 1
transform 1 0 1104 0 -1 137088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_247_Right_33
timestamp 1
transform -1 0 108836 0 -1 137088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_248_Left_514
timestamp 1
transform 1 0 1104 0 1 137088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_248_Right_34
timestamp 1
transform -1 0 108836 0 1 137088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_249_Left_515
timestamp 1
transform 1 0 1104 0 -1 138176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_249_Right_35
timestamp 1
transform -1 0 108836 0 -1 138176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_250_Left_516
timestamp 1
transform 1 0 1104 0 1 138176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_250_Right_36
timestamp 1
transform -1 0 108836 0 1 138176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_251_Left_517
timestamp 1
transform 1 0 1104 0 -1 139264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_251_Right_37
timestamp 1
transform -1 0 108836 0 -1 139264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_252_Left_518
timestamp 1
transform 1 0 1104 0 1 139264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_252_Right_38
timestamp 1
transform -1 0 108836 0 1 139264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_253_Left_519
timestamp 1
transform 1 0 1104 0 -1 140352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_253_Right_39
timestamp 1
transform -1 0 108836 0 -1 140352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_254_Left_520
timestamp 1
transform 1 0 1104 0 1 140352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_254_Right_40
timestamp 1
transform -1 0 108836 0 1 140352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_255_Left_521
timestamp 1
transform 1 0 1104 0 -1 141440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_255_Right_41
timestamp 1
transform -1 0 108836 0 -1 141440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_256_Left_522
timestamp 1
transform 1 0 1104 0 1 141440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_256_Right_42
timestamp 1
transform -1 0 108836 0 1 141440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_257_Left_523
timestamp 1
transform 1 0 1104 0 -1 142528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_257_Right_43
timestamp 1
transform -1 0 108836 0 -1 142528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_258_Left_524
timestamp 1
transform 1 0 1104 0 1 142528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_258_Right_44
timestamp 1
transform -1 0 108836 0 1 142528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_259_Left_525
timestamp 1
transform 1 0 1104 0 -1 143616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_259_Right_45
timestamp 1
transform -1 0 108836 0 -1 143616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_260_Left_526
timestamp 1
transform 1 0 1104 0 1 143616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_260_Right_46
timestamp 1
transform -1 0 108836 0 1 143616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_261_Left_527
timestamp 1
transform 1 0 1104 0 -1 144704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_261_Right_47
timestamp 1
transform -1 0 108836 0 -1 144704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_262_Left_528
timestamp 1
transform 1 0 1104 0 1 144704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_262_Right_48
timestamp 1
transform -1 0 108836 0 1 144704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_263_Left_529
timestamp 1
transform 1 0 1104 0 -1 145792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_263_Right_49
timestamp 1
transform -1 0 108836 0 -1 145792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_264_Left_530
timestamp 1
transform 1 0 1104 0 1 145792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_264_Right_50
timestamp 1
transform -1 0 108836 0 1 145792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_265_Left_531
timestamp 1
transform 1 0 1104 0 -1 146880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_265_Right_51
timestamp 1
transform -1 0 108836 0 -1 146880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_266_Left_532
timestamp 1
transform 1 0 1104 0 1 146880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_266_Right_52
timestamp 1
transform -1 0 108836 0 1 146880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_962
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_963
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_964
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_965
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_966
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_967
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_968
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_969
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_970
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_971
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_972
timestamp 1
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_973
timestamp 1
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_974
timestamp 1
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_975
timestamp 1
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_976
timestamp 1
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_977
timestamp 1
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_978
timestamp 1
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_979
timestamp 1
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_980
timestamp 1
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_981
timestamp 1
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_982
timestamp 1
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_983
timestamp 1
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_984
timestamp 1
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_985
timestamp 1
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_986
timestamp 1
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_987
timestamp 1
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_988
timestamp 1
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_989
timestamp 1
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_990
timestamp 1
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_991
timestamp 1
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_992
timestamp 1
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_993
timestamp 1
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_994
timestamp 1
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_995
timestamp 1
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_996
timestamp 1
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_997
timestamp 1
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_998
timestamp 1
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_999
timestamp 1
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_1000
timestamp 1
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_1001
timestamp 1
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_1002
timestamp 1
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1003
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1004
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1005
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1006
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1007
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1008
timestamp 1
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1009
timestamp 1
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1010
timestamp 1
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1011
timestamp 1
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1012
timestamp 1
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1013
timestamp 1
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1014
timestamp 1
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1015
timestamp 1
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1016
timestamp 1
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1017
timestamp 1
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1018
timestamp 1
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1019
timestamp 1
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1020
timestamp 1
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1021
timestamp 1
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1022
timestamp 1
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1023
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1024
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1025
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1026
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1027
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1028
timestamp 1
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1029
timestamp 1
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1030
timestamp 1
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1031
timestamp 1
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1032
timestamp 1
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1033
timestamp 1
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1034
timestamp 1
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1035
timestamp 1
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1036
timestamp 1
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1037
timestamp 1
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1038
timestamp 1
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1039
timestamp 1
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1040
timestamp 1
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1041
timestamp 1
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1042
timestamp 1
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1043
timestamp 1
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1044
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1045
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1046
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1047
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1048
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1049
timestamp 1
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1050
timestamp 1
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1051
timestamp 1
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1052
timestamp 1
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1053
timestamp 1
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1054
timestamp 1
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1055
timestamp 1
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1056
timestamp 1
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1057
timestamp 1
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1058
timestamp 1
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1059
timestamp 1
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1060
timestamp 1
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1061
timestamp 1
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1062
timestamp 1
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1063
timestamp 1
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1064
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1065
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1066
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1067
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1068
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1069
timestamp 1
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1070
timestamp 1
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1071
timestamp 1
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1072
timestamp 1
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1073
timestamp 1
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1074
timestamp 1
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1075
timestamp 1
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1076
timestamp 1
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1077
timestamp 1
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1078
timestamp 1
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1079
timestamp 1
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1080
timestamp 1
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1081
timestamp 1
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1082
timestamp 1
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1083
timestamp 1
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1084
timestamp 1
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1085
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1086
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1087
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1088
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1089
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1090
timestamp 1
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1091
timestamp 1
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1092
timestamp 1
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1093
timestamp 1
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1094
timestamp 1
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1095
timestamp 1
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1096
timestamp 1
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1097
timestamp 1
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1098
timestamp 1
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1099
timestamp 1
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1100
timestamp 1
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1101
timestamp 1
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1102
timestamp 1
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1103
timestamp 1
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1104
timestamp 1
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1105
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1106
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1107
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1108
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1109
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1110
timestamp 1
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1111
timestamp 1
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1112
timestamp 1
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1113
timestamp 1
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1114
timestamp 1
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1115
timestamp 1
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1116
timestamp 1
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1117
timestamp 1
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1118
timestamp 1
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1119
timestamp 1
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1120
timestamp 1
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1121
timestamp 1
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1122
timestamp 1
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1123
timestamp 1
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1124
timestamp 1
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1125
timestamp 1
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1126
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1127
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1128
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1129
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1130
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1131
timestamp 1
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1132
timestamp 1
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1133
timestamp 1
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1134
timestamp 1
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1135
timestamp 1
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1136
timestamp 1
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1137
timestamp 1
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1138
timestamp 1
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1139
timestamp 1
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1140
timestamp 1
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1141
timestamp 1
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1142
timestamp 1
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1143
timestamp 1
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1144
timestamp 1
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1145
timestamp 1
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1146
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1147
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1148
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1149
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1150
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1151
timestamp 1
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1152
timestamp 1
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1153
timestamp 1
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1154
timestamp 1
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1155
timestamp 1
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1156
timestamp 1
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1157
timestamp 1
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1158
timestamp 1
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1159
timestamp 1
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1160
timestamp 1
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1161
timestamp 1
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1162
timestamp 1
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1163
timestamp 1
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1164
timestamp 1
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1165
timestamp 1
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1166
timestamp 1
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1167
timestamp 1
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1168
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1169
timestamp 1
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1170
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1171
timestamp 1
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1172
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1173
timestamp 1
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1174
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1175
timestamp 1
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1176
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1177
timestamp 1
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1178
timestamp 1
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1179
timestamp 1
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1180
timestamp 1
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1181
timestamp 1
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1182
timestamp 1
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1183
timestamp 1
transform 1 0 44896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1184
timestamp 1
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1185
timestamp 1
transform 1 0 50048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1186
timestamp 1
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1187
timestamp 1
transform 1 0 55200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1188
timestamp 1
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1189
timestamp 1
transform 1 0 60352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1190
timestamp 1
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1191
timestamp 1
transform 1 0 65504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1192
timestamp 1
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1193
timestamp 1
transform 1 0 70656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1194
timestamp 1
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1195
timestamp 1
transform 1 0 75808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1196
timestamp 1
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1197
timestamp 1
transform 1 0 80960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1198
timestamp 1
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1199
timestamp 1
transform 1 0 86112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1200
timestamp 1
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1201
timestamp 1
transform 1 0 91264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1202
timestamp 1
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1203
timestamp 1
transform 1 0 96416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1204
timestamp 1
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1205
timestamp 1
transform 1 0 101568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1206
timestamp 1
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1207
timestamp 1
transform 1 0 106720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_2384
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_2385
timestamp 1
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_1_1208
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_1209
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_2386
timestamp 1
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_1_1210
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_1_1211
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_2387
timestamp 1
transform 1 0 106628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_1_1212
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_1_1213
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_2388
timestamp 1
transform 1 0 106628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_1_1214
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_1_1215
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_2389
timestamp 1
transform 1 0 106628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_1_1216
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_1_1217
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_2390
timestamp 1
transform 1 0 106628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_1_1218
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_1_1219
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_2391
timestamp 1
transform 1 0 106628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_1_1220
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_1_1221
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_2392
timestamp 1
transform 1 0 106628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_1_1222
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_1_1223
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_2393
timestamp 1
transform 1 0 106628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_1_1224
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_1_1225
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_2394
timestamp 1
transform 1 0 106628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_1_1226
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_1_1227
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_2395
timestamp 1
transform 1 0 106628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_1_1228
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_1_1229
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_2396
timestamp 1
transform 1 0 106628 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_1_1230
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_1_1231
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_2397
timestamp 1
transform 1 0 106628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_1_1232
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_1_1233
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_2398
timestamp 1
transform 1 0 106628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_1_1234
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_1_1235
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_2399
timestamp 1
transform 1 0 106628 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_1_1236
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_1_1237
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_2400
timestamp 1
transform 1 0 106628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_1_1238
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_1_1239
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_2401
timestamp 1
transform 1 0 106628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_1_1240
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_1_1241
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_2402
timestamp 1
transform 1 0 106628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_1_1242
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_1_1243
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_2403
timestamp 1
transform 1 0 106628 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_1_1244
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1_1245
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_2404
timestamp 1
transform 1 0 106628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1_1246
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1_1247
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_2405
timestamp 1
transform 1 0 106628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1_1248
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1_1249
timestamp 1
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_2406
timestamp 1
transform 1 0 106628 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1_1250
timestamp 1
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1_1251
timestamp 1
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_2407
timestamp 1
transform 1 0 106628 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1_1252
timestamp 1
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1_1253
timestamp 1
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_2408
timestamp 1
transform 1 0 106628 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1_1254
timestamp 1
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1_1255
timestamp 1
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_2409
timestamp 1
transform 1 0 106628 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1_1256
timestamp 1
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1_1257
timestamp 1
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_2410
timestamp 1
transform 1 0 106628 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1_1258
timestamp 1
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1_1259
timestamp 1
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_2411
timestamp 1
transform 1 0 106628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1_1260
timestamp 1
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1_1261
timestamp 1
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_2412
timestamp 1
transform 1 0 106628 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1_1262
timestamp 1
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1_1263
timestamp 1
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_2413
timestamp 1
transform 1 0 106628 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1_1264
timestamp 1
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1_1265
timestamp 1
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_2414
timestamp 1
transform 1 0 106628 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1_1266
timestamp 1
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1_1267
timestamp 1
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_2415
timestamp 1
transform 1 0 106628 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1_1268
timestamp 1
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1_1269
timestamp 1
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_2416
timestamp 1
transform 1 0 106628 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1_1270
timestamp 1
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1_1271
timestamp 1
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_2417
timestamp 1
transform 1 0 106628 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1_1272
timestamp 1
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1_1273
timestamp 1
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_2418
timestamp 1
transform 1 0 106628 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1_1274
timestamp 1
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1_1275
timestamp 1
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_2419
timestamp 1
transform 1 0 106628 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1_1276
timestamp 1
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1_1277
timestamp 1
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_2420
timestamp 1
transform 1 0 106628 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1_1278
timestamp 1
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1_1279
timestamp 1
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_2421
timestamp 1
transform 1 0 106628 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1_1280
timestamp 1
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1_1281
timestamp 1
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_2422
timestamp 1
transform 1 0 106628 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1_1282
timestamp 1
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1_1283
timestamp 1
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_2423
timestamp 1
transform 1 0 106628 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1_1284
timestamp 1
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1_1285
timestamp 1
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_2424
timestamp 1
transform 1 0 106628 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1_1286
timestamp 1
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1_1287
timestamp 1
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_2425
timestamp 1
transform 1 0 106628 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1_1288
timestamp 1
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1_1289
timestamp 1
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_2426
timestamp 1
transform 1 0 106628 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1_1290
timestamp 1
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1_1291
timestamp 1
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_2427
timestamp 1
transform 1 0 106628 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1_1292
timestamp 1
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1_1293
timestamp 1
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_2428
timestamp 1
transform 1 0 106628 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1_1294
timestamp 1
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1_1295
timestamp 1
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_2429
timestamp 1
transform 1 0 106628 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1_1296
timestamp 1
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1_1297
timestamp 1
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_2430
timestamp 1
transform 1 0 106628 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1_1298
timestamp 1
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1_1299
timestamp 1
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_2431
timestamp 1
transform 1 0 106628 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1_1300
timestamp 1
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1_1301
timestamp 1
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_2432
timestamp 1
transform 1 0 106628 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1_1302
timestamp 1
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1_1303
timestamp 1
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_2433
timestamp 1
transform 1 0 106628 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1_1304
timestamp 1
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1_1305
timestamp 1
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_2434
timestamp 1
transform 1 0 106628 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1_1306
timestamp 1
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1_1307
timestamp 1
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_2435
timestamp 1
transform 1 0 106628 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1_1308
timestamp 1
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1_1309
timestamp 1
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_2436
timestamp 1
transform 1 0 106628 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1_1310
timestamp 1
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1_1311
timestamp 1
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_2437
timestamp 1
transform 1 0 106628 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1_1312
timestamp 1
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1_1313
timestamp 1
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_2438
timestamp 1
transform 1 0 106628 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1315
timestamp 1
transform 1 0 3680 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1316
timestamp 1
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1317
timestamp 1
transform 1 0 8832 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1318
timestamp 1
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1319
timestamp 1
transform 1 0 13984 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1320
timestamp 1
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1321
timestamp 1
transform 1 0 19136 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1322
timestamp 1
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1323
timestamp 1
transform 1 0 24288 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1324
timestamp 1
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1325
timestamp 1
transform 1 0 29440 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1326
timestamp 1
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1327
timestamp 1
transform 1 0 34592 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1328
timestamp 1
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1329
timestamp 1
transform 1 0 39744 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1330
timestamp 1
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1331
timestamp 1
transform 1 0 44896 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1332
timestamp 1
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1333
timestamp 1
transform 1 0 50048 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1334
timestamp 1
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1335
timestamp 1
transform 1 0 55200 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1336
timestamp 1
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1337
timestamp 1
transform 1 0 60352 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1338
timestamp 1
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1339
timestamp 1
transform 1 0 65504 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1340
timestamp 1
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1341
timestamp 1
transform 1 0 70656 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1342
timestamp 1
transform 1 0 73232 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1343
timestamp 1
transform 1 0 75808 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1344
timestamp 1
transform 1 0 78384 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1345
timestamp 1
transform 1 0 80960 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1346
timestamp 1
transform 1 0 83536 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1347
timestamp 1
transform 1 0 86112 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1348
timestamp 1
transform 1 0 88688 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1349
timestamp 1
transform 1 0 91264 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1350
timestamp 1
transform 1 0 93840 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1351
timestamp 1
transform 1 0 96416 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1352
timestamp 1
transform 1 0 98992 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1353
timestamp 1
transform 1 0 101568 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1354
timestamp 1
transform 1 0 104144 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1355
timestamp 1
transform 1 0 106720 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1356
timestamp 1
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1357
timestamp 1
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1358
timestamp 1
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1359
timestamp 1
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1360
timestamp 1
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1361
timestamp 1
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1362
timestamp 1
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1363
timestamp 1
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1364
timestamp 1
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1365
timestamp 1
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1366
timestamp 1
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1367
timestamp 1
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1368
timestamp 1
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1369
timestamp 1
transform 1 0 70656 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1370
timestamp 1
transform 1 0 75808 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1371
timestamp 1
transform 1 0 80960 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1372
timestamp 1
transform 1 0 86112 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1373
timestamp 1
transform 1 0 91264 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1374
timestamp 1
transform 1 0 96416 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1375
timestamp 1
transform 1 0 101568 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1376
timestamp 1
transform 1 0 106720 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1377
timestamp 1
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1378
timestamp 1
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1379
timestamp 1
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1380
timestamp 1
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1381
timestamp 1
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1382
timestamp 1
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1383
timestamp 1
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1384
timestamp 1
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1385
timestamp 1
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1386
timestamp 1
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1387
timestamp 1
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1388
timestamp 1
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1389
timestamp 1
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1390
timestamp 1
transform 1 0 73232 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1391
timestamp 1
transform 1 0 78384 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1392
timestamp 1
transform 1 0 83536 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1393
timestamp 1
transform 1 0 88688 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1394
timestamp 1
transform 1 0 93840 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1395
timestamp 1
transform 1 0 98992 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1396
timestamp 1
transform 1 0 104144 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1397
timestamp 1
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1398
timestamp 1
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1399
timestamp 1
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1400
timestamp 1
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1401
timestamp 1
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1402
timestamp 1
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1403
timestamp 1
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1404
timestamp 1
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1405
timestamp 1
transform 1 0 44896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1406
timestamp 1
transform 1 0 50048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1407
timestamp 1
transform 1 0 55200 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1408
timestamp 1
transform 1 0 60352 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1409
timestamp 1
transform 1 0 65504 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1410
timestamp 1
transform 1 0 70656 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1411
timestamp 1
transform 1 0 75808 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1412
timestamp 1
transform 1 0 80960 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1413
timestamp 1
transform 1 0 86112 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1414
timestamp 1
transform 1 0 91264 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1415
timestamp 1
transform 1 0 96416 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1416
timestamp 1
transform 1 0 101568 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1417
timestamp 1
transform 1 0 106720 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1418
timestamp 1
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1419
timestamp 1
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1420
timestamp 1
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1421
timestamp 1
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1422
timestamp 1
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1423
timestamp 1
transform 1 0 32016 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1424
timestamp 1
transform 1 0 37168 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1425
timestamp 1
transform 1 0 42320 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1426
timestamp 1
transform 1 0 47472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1427
timestamp 1
transform 1 0 52624 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1428
timestamp 1
transform 1 0 57776 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1429
timestamp 1
transform 1 0 62928 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1430
timestamp 1
transform 1 0 68080 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1431
timestamp 1
transform 1 0 73232 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1432
timestamp 1
transform 1 0 78384 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1433
timestamp 1
transform 1 0 83536 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1434
timestamp 1
transform 1 0 88688 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1435
timestamp 1
transform 1 0 93840 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1436
timestamp 1
transform 1 0 98992 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1437
timestamp 1
transform 1 0 104144 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1438
timestamp 1
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1439
timestamp 1
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1440
timestamp 1
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1441
timestamp 1
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1442
timestamp 1
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1443
timestamp 1
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1444
timestamp 1
transform 1 0 34592 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1445
timestamp 1
transform 1 0 39744 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1446
timestamp 1
transform 1 0 44896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1447
timestamp 1
transform 1 0 50048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1448
timestamp 1
transform 1 0 55200 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1449
timestamp 1
transform 1 0 60352 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1450
timestamp 1
transform 1 0 65504 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1451
timestamp 1
transform 1 0 70656 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1452
timestamp 1
transform 1 0 75808 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1453
timestamp 1
transform 1 0 80960 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1454
timestamp 1
transform 1 0 86112 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1455
timestamp 1
transform 1 0 91264 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1456
timestamp 1
transform 1 0 96416 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1457
timestamp 1
transform 1 0 101568 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1458
timestamp 1
transform 1 0 106720 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1459
timestamp 1
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1460
timestamp 1
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1461
timestamp 1
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1462
timestamp 1
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1463
timestamp 1
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1464
timestamp 1
transform 1 0 32016 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1465
timestamp 1
transform 1 0 37168 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1466
timestamp 1
transform 1 0 42320 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1467
timestamp 1
transform 1 0 47472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1468
timestamp 1
transform 1 0 52624 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1469
timestamp 1
transform 1 0 57776 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1470
timestamp 1
transform 1 0 62928 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1471
timestamp 1
transform 1 0 68080 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1472
timestamp 1
transform 1 0 73232 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1473
timestamp 1
transform 1 0 78384 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1474
timestamp 1
transform 1 0 83536 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1475
timestamp 1
transform 1 0 88688 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1476
timestamp 1
transform 1 0 93840 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1477
timestamp 1
transform 1 0 98992 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1478
timestamp 1
transform 1 0 104144 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1479
timestamp 1
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1480
timestamp 1
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1481
timestamp 1
transform 1 0 13984 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1482
timestamp 1
transform 1 0 19136 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1483
timestamp 1
transform 1 0 24288 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1484
timestamp 1
transform 1 0 29440 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1485
timestamp 1
transform 1 0 34592 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1486
timestamp 1
transform 1 0 39744 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1487
timestamp 1
transform 1 0 44896 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1488
timestamp 1
transform 1 0 50048 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1489
timestamp 1
transform 1 0 55200 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1490
timestamp 1
transform 1 0 60352 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1491
timestamp 1
transform 1 0 65504 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1492
timestamp 1
transform 1 0 70656 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1493
timestamp 1
transform 1 0 75808 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1494
timestamp 1
transform 1 0 80960 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1495
timestamp 1
transform 1 0 86112 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1496
timestamp 1
transform 1 0 91264 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1497
timestamp 1
transform 1 0 96416 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1498
timestamp 1
transform 1 0 101568 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1499
timestamp 1
transform 1 0 106720 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1500
timestamp 1
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1501
timestamp 1
transform 1 0 11408 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1502
timestamp 1
transform 1 0 16560 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1503
timestamp 1
transform 1 0 21712 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1504
timestamp 1
transform 1 0 26864 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1505
timestamp 1
transform 1 0 32016 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1506
timestamp 1
transform 1 0 37168 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1507
timestamp 1
transform 1 0 42320 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1508
timestamp 1
transform 1 0 47472 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1509
timestamp 1
transform 1 0 52624 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1510
timestamp 1
transform 1 0 57776 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1511
timestamp 1
transform 1 0 62928 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1512
timestamp 1
transform 1 0 68080 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1513
timestamp 1
transform 1 0 73232 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1514
timestamp 1
transform 1 0 78384 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1515
timestamp 1
transform 1 0 83536 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1516
timestamp 1
transform 1 0 88688 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1517
timestamp 1
transform 1 0 93840 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1518
timestamp 1
transform 1 0 98992 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1519
timestamp 1
transform 1 0 104144 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1520
timestamp 1
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1521
timestamp 1
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1522
timestamp 1
transform 1 0 13984 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1523
timestamp 1
transform 1 0 19136 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1524
timestamp 1
transform 1 0 24288 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1525
timestamp 1
transform 1 0 29440 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1526
timestamp 1
transform 1 0 34592 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1527
timestamp 1
transform 1 0 39744 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1528
timestamp 1
transform 1 0 44896 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1529
timestamp 1
transform 1 0 50048 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1530
timestamp 1
transform 1 0 55200 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1531
timestamp 1
transform 1 0 60352 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1532
timestamp 1
transform 1 0 65504 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1533
timestamp 1
transform 1 0 70656 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1534
timestamp 1
transform 1 0 75808 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1535
timestamp 1
transform 1 0 80960 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1536
timestamp 1
transform 1 0 86112 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1537
timestamp 1
transform 1 0 91264 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1538
timestamp 1
transform 1 0 96416 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1539
timestamp 1
transform 1 0 101568 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1540
timestamp 1
transform 1 0 106720 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1541
timestamp 1
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1542
timestamp 1
transform 1 0 11408 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1543
timestamp 1
transform 1 0 16560 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1544
timestamp 1
transform 1 0 21712 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1545
timestamp 1
transform 1 0 26864 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1546
timestamp 1
transform 1 0 32016 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1547
timestamp 1
transform 1 0 37168 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1548
timestamp 1
transform 1 0 42320 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1549
timestamp 1
transform 1 0 47472 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1550
timestamp 1
transform 1 0 52624 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1551
timestamp 1
transform 1 0 57776 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1552
timestamp 1
transform 1 0 62928 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1553
timestamp 1
transform 1 0 68080 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1554
timestamp 1
transform 1 0 73232 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1555
timestamp 1
transform 1 0 78384 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1556
timestamp 1
transform 1 0 83536 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1557
timestamp 1
transform 1 0 88688 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1558
timestamp 1
transform 1 0 93840 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1559
timestamp 1
transform 1 0 98992 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1560
timestamp 1
transform 1 0 104144 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1561
timestamp 1
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1562
timestamp 1
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1563
timestamp 1
transform 1 0 13984 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1564
timestamp 1
transform 1 0 19136 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1565
timestamp 1
transform 1 0 24288 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1566
timestamp 1
transform 1 0 29440 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1567
timestamp 1
transform 1 0 34592 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1568
timestamp 1
transform 1 0 39744 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1569
timestamp 1
transform 1 0 44896 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1570
timestamp 1
transform 1 0 50048 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1571
timestamp 1
transform 1 0 55200 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1572
timestamp 1
transform 1 0 60352 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1573
timestamp 1
transform 1 0 65504 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1574
timestamp 1
transform 1 0 70656 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1575
timestamp 1
transform 1 0 75808 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1576
timestamp 1
transform 1 0 80960 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1577
timestamp 1
transform 1 0 86112 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1578
timestamp 1
transform 1 0 91264 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1579
timestamp 1
transform 1 0 96416 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1580
timestamp 1
transform 1 0 101568 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1581
timestamp 1
transform 1 0 106720 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1582
timestamp 1
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1583
timestamp 1
transform 1 0 11408 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1584
timestamp 1
transform 1 0 16560 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1585
timestamp 1
transform 1 0 21712 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1586
timestamp 1
transform 1 0 26864 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1587
timestamp 1
transform 1 0 32016 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1588
timestamp 1
transform 1 0 37168 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1589
timestamp 1
transform 1 0 42320 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1590
timestamp 1
transform 1 0 47472 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1591
timestamp 1
transform 1 0 52624 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1592
timestamp 1
transform 1 0 57776 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1593
timestamp 1
transform 1 0 62928 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1594
timestamp 1
transform 1 0 68080 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1595
timestamp 1
transform 1 0 73232 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1596
timestamp 1
transform 1 0 78384 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1597
timestamp 1
transform 1 0 83536 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1598
timestamp 1
transform 1 0 88688 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1599
timestamp 1
transform 1 0 93840 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1600
timestamp 1
transform 1 0 98992 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1601
timestamp 1
transform 1 0 104144 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1602
timestamp 1
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1603
timestamp 1
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1604
timestamp 1
transform 1 0 13984 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1605
timestamp 1
transform 1 0 19136 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1606
timestamp 1
transform 1 0 24288 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1607
timestamp 1
transform 1 0 29440 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1608
timestamp 1
transform 1 0 34592 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1609
timestamp 1
transform 1 0 39744 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1610
timestamp 1
transform 1 0 44896 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1611
timestamp 1
transform 1 0 50048 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1612
timestamp 1
transform 1 0 55200 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1613
timestamp 1
transform 1 0 60352 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1614
timestamp 1
transform 1 0 65504 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1615
timestamp 1
transform 1 0 70656 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1616
timestamp 1
transform 1 0 75808 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1617
timestamp 1
transform 1 0 80960 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1618
timestamp 1
transform 1 0 86112 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1619
timestamp 1
transform 1 0 91264 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1620
timestamp 1
transform 1 0 96416 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1621
timestamp 1
transform 1 0 101568 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1622
timestamp 1
transform 1 0 106720 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1623
timestamp 1
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1624
timestamp 1
transform 1 0 11408 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1625
timestamp 1
transform 1 0 16560 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1626
timestamp 1
transform 1 0 21712 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1627
timestamp 1
transform 1 0 26864 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1628
timestamp 1
transform 1 0 32016 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1629
timestamp 1
transform 1 0 37168 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1630
timestamp 1
transform 1 0 42320 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1631
timestamp 1
transform 1 0 47472 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1632
timestamp 1
transform 1 0 52624 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1633
timestamp 1
transform 1 0 57776 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1634
timestamp 1
transform 1 0 62928 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1635
timestamp 1
transform 1 0 68080 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1636
timestamp 1
transform 1 0 73232 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1637
timestamp 1
transform 1 0 78384 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1638
timestamp 1
transform 1 0 83536 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1639
timestamp 1
transform 1 0 88688 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1640
timestamp 1
transform 1 0 93840 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1641
timestamp 1
transform 1 0 98992 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1642
timestamp 1
transform 1 0 104144 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1643
timestamp 1
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1644
timestamp 1
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1645
timestamp 1
transform 1 0 13984 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1646
timestamp 1
transform 1 0 19136 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1647
timestamp 1
transform 1 0 24288 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1648
timestamp 1
transform 1 0 29440 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1649
timestamp 1
transform 1 0 34592 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1650
timestamp 1
transform 1 0 39744 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1651
timestamp 1
transform 1 0 44896 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1652
timestamp 1
transform 1 0 50048 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1653
timestamp 1
transform 1 0 55200 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1654
timestamp 1
transform 1 0 60352 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1655
timestamp 1
transform 1 0 65504 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1656
timestamp 1
transform 1 0 70656 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1657
timestamp 1
transform 1 0 75808 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1658
timestamp 1
transform 1 0 80960 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1659
timestamp 1
transform 1 0 86112 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1660
timestamp 1
transform 1 0 91264 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1661
timestamp 1
transform 1 0 96416 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1662
timestamp 1
transform 1 0 101568 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1663
timestamp 1
transform 1 0 106720 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1664
timestamp 1
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1665
timestamp 1
transform 1 0 11408 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1666
timestamp 1
transform 1 0 16560 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1667
timestamp 1
transform 1 0 21712 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1668
timestamp 1
transform 1 0 26864 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1669
timestamp 1
transform 1 0 32016 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1670
timestamp 1
transform 1 0 37168 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1671
timestamp 1
transform 1 0 42320 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1672
timestamp 1
transform 1 0 47472 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1673
timestamp 1
transform 1 0 52624 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1674
timestamp 1
transform 1 0 57776 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1675
timestamp 1
transform 1 0 62928 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1676
timestamp 1
transform 1 0 68080 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1677
timestamp 1
transform 1 0 73232 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1678
timestamp 1
transform 1 0 78384 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1679
timestamp 1
transform 1 0 83536 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1680
timestamp 1
transform 1 0 88688 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1681
timestamp 1
transform 1 0 93840 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1682
timestamp 1
transform 1 0 98992 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1683
timestamp 1
transform 1 0 104144 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1684
timestamp 1
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1685
timestamp 1
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1686
timestamp 1
transform 1 0 13984 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1687
timestamp 1
transform 1 0 19136 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1688
timestamp 1
transform 1 0 24288 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1689
timestamp 1
transform 1 0 29440 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1690
timestamp 1
transform 1 0 34592 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1691
timestamp 1
transform 1 0 39744 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1692
timestamp 1
transform 1 0 44896 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1693
timestamp 1
transform 1 0 50048 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1694
timestamp 1
transform 1 0 55200 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1695
timestamp 1
transform 1 0 60352 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1696
timestamp 1
transform 1 0 65504 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1697
timestamp 1
transform 1 0 70656 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1698
timestamp 1
transform 1 0 75808 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1699
timestamp 1
transform 1 0 80960 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1700
timestamp 1
transform 1 0 86112 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1701
timestamp 1
transform 1 0 91264 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1702
timestamp 1
transform 1 0 96416 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1703
timestamp 1
transform 1 0 101568 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1704
timestamp 1
transform 1 0 106720 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1705
timestamp 1
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1706
timestamp 1
transform 1 0 11408 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1707
timestamp 1
transform 1 0 16560 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1708
timestamp 1
transform 1 0 21712 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1709
timestamp 1
transform 1 0 26864 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1710
timestamp 1
transform 1 0 32016 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1711
timestamp 1
transform 1 0 37168 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1712
timestamp 1
transform 1 0 42320 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1713
timestamp 1
transform 1 0 47472 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1714
timestamp 1
transform 1 0 52624 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1715
timestamp 1
transform 1 0 57776 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1716
timestamp 1
transform 1 0 62928 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1717
timestamp 1
transform 1 0 68080 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1718
timestamp 1
transform 1 0 73232 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1719
timestamp 1
transform 1 0 78384 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1720
timestamp 1
transform 1 0 83536 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1721
timestamp 1
transform 1 0 88688 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1722
timestamp 1
transform 1 0 93840 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1723
timestamp 1
transform 1 0 98992 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1724
timestamp 1
transform 1 0 104144 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1725
timestamp 1
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1726
timestamp 1
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1727
timestamp 1
transform 1 0 13984 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1728
timestamp 1
transform 1 0 19136 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1729
timestamp 1
transform 1 0 24288 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1730
timestamp 1
transform 1 0 29440 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1731
timestamp 1
transform 1 0 34592 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1732
timestamp 1
transform 1 0 39744 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1733
timestamp 1
transform 1 0 44896 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1734
timestamp 1
transform 1 0 50048 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1735
timestamp 1
transform 1 0 55200 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1736
timestamp 1
transform 1 0 60352 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1737
timestamp 1
transform 1 0 65504 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1738
timestamp 1
transform 1 0 70656 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1739
timestamp 1
transform 1 0 75808 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1740
timestamp 1
transform 1 0 80960 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1741
timestamp 1
transform 1 0 86112 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1742
timestamp 1
transform 1 0 91264 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1743
timestamp 1
transform 1 0 96416 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1744
timestamp 1
transform 1 0 101568 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1745
timestamp 1
transform 1 0 106720 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1746
timestamp 1
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1747
timestamp 1
transform 1 0 11408 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1748
timestamp 1
transform 1 0 16560 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1749
timestamp 1
transform 1 0 21712 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1750
timestamp 1
transform 1 0 26864 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1751
timestamp 1
transform 1 0 32016 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1752
timestamp 1
transform 1 0 37168 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1753
timestamp 1
transform 1 0 42320 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1754
timestamp 1
transform 1 0 47472 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1755
timestamp 1
transform 1 0 52624 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1756
timestamp 1
transform 1 0 57776 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1757
timestamp 1
transform 1 0 62928 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1758
timestamp 1
transform 1 0 68080 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1759
timestamp 1
transform 1 0 73232 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1760
timestamp 1
transform 1 0 78384 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1761
timestamp 1
transform 1 0 83536 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1762
timestamp 1
transform 1 0 88688 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1763
timestamp 1
transform 1 0 93840 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1764
timestamp 1
transform 1 0 98992 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1765
timestamp 1
transform 1 0 104144 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1766
timestamp 1
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1767
timestamp 1
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1768
timestamp 1
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1769
timestamp 1
transform 1 0 11408 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1770
timestamp 1
transform 1 0 13984 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1771
timestamp 1
transform 1 0 16560 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1772
timestamp 1
transform 1 0 19136 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1773
timestamp 1
transform 1 0 21712 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1774
timestamp 1
transform 1 0 24288 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1775
timestamp 1
transform 1 0 26864 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1776
timestamp 1
transform 1 0 29440 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1777
timestamp 1
transform 1 0 32016 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1778
timestamp 1
transform 1 0 34592 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1779
timestamp 1
transform 1 0 37168 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1780
timestamp 1
transform 1 0 39744 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1781
timestamp 1
transform 1 0 42320 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1782
timestamp 1
transform 1 0 44896 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1783
timestamp 1
transform 1 0 47472 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1784
timestamp 1
transform 1 0 50048 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1785
timestamp 1
transform 1 0 52624 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1786
timestamp 1
transform 1 0 55200 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1787
timestamp 1
transform 1 0 57776 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1788
timestamp 1
transform 1 0 60352 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1789
timestamp 1
transform 1 0 62928 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1790
timestamp 1
transform 1 0 65504 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1791
timestamp 1
transform 1 0 68080 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1792
timestamp 1
transform 1 0 70656 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1793
timestamp 1
transform 1 0 73232 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1794
timestamp 1
transform 1 0 75808 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1795
timestamp 1
transform 1 0 78384 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1796
timestamp 1
transform 1 0 80960 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1797
timestamp 1
transform 1 0 83536 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1798
timestamp 1
transform 1 0 86112 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1799
timestamp 1
transform 1 0 88688 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1800
timestamp 1
transform 1 0 91264 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1801
timestamp 1
transform 1 0 93840 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1802
timestamp 1
transform 1 0 96416 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1803
timestamp 1
transform 1 0 98992 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1804
timestamp 1
transform 1 0 101568 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1805
timestamp 1
transform 1 0 104144 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1806
timestamp 1
transform 1 0 106720 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1_1314
timestamp 1
transform 1 0 6256 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1_1807
timestamp 1
transform 1 0 3680 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_2439
timestamp 1
transform 1 0 106628 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1_1808
timestamp 1
transform 1 0 6256 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1_1809
timestamp 1
transform 1 0 3680 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_2440
timestamp 1
transform 1 0 106628 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1_1810
timestamp 1
transform 1 0 6256 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1_1811
timestamp 1
transform 1 0 3680 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_2441
timestamp 1
transform 1 0 106628 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1_1812
timestamp 1
transform 1 0 6256 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1_1813
timestamp 1
transform 1 0 3680 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_2442
timestamp 1
transform 1 0 106628 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1_1814
timestamp 1
transform 1 0 6256 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1_1815
timestamp 1
transform 1 0 3680 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_2443
timestamp 1
transform 1 0 106628 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1_1816
timestamp 1
transform 1 0 6256 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1_1817
timestamp 1
transform 1 0 3680 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_2444
timestamp 1
transform 1 0 106628 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1_1818
timestamp 1
transform 1 0 6256 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1_1819
timestamp 1
transform 1 0 3680 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_2445
timestamp 1
transform 1 0 106628 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1_1820
timestamp 1
transform 1 0 6256 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1_1821
timestamp 1
transform 1 0 3680 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_2446
timestamp 1
transform 1 0 106628 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1_1822
timestamp 1
transform 1 0 6256 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1_1823
timestamp 1
transform 1 0 3680 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_2_2447
timestamp 1
transform 1 0 106628 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1_1824
timestamp 1
transform 1 0 6256 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1_1825
timestamp 1
transform 1 0 3680 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_2_2448
timestamp 1
transform 1 0 106628 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1_1826
timestamp 1
transform 1 0 6256 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1_1827
timestamp 1
transform 1 0 3680 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_2_2449
timestamp 1
transform 1 0 106628 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1_1828
timestamp 1
transform 1 0 6256 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1_1829
timestamp 1
transform 1 0 3680 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_2_2450
timestamp 1
transform 1 0 106628 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1_1830
timestamp 1
transform 1 0 6256 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1_1831
timestamp 1
transform 1 0 3680 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_2_2451
timestamp 1
transform 1 0 106628 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1_1832
timestamp 1
transform 1 0 6256 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1_1833
timestamp 1
transform 1 0 3680 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_2_2452
timestamp 1
transform 1 0 106628 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1_1834
timestamp 1
transform 1 0 6256 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1_1835
timestamp 1
transform 1 0 3680 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_2_2453
timestamp 1
transform 1 0 106628 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1_1836
timestamp 1
transform 1 0 6256 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1_1837
timestamp 1
transform 1 0 3680 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_2_2454
timestamp 1
transform 1 0 106628 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1_1838
timestamp 1
transform 1 0 6256 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1_1839
timestamp 1
transform 1 0 3680 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_2_2455
timestamp 1
transform 1 0 106628 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1_1840
timestamp 1
transform 1 0 6256 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1_1841
timestamp 1
transform 1 0 3680 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_2_2456
timestamp 1
transform 1 0 106628 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1_1842
timestamp 1
transform 1 0 6256 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1_1843
timestamp 1
transform 1 0 3680 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_2_2457
timestamp 1
transform 1 0 106628 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1_1844
timestamp 1
transform 1 0 6256 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1_1845
timestamp 1
transform 1 0 3680 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_2_2458
timestamp 1
transform 1 0 106628 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1_1846
timestamp 1
transform 1 0 6256 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_1_1847
timestamp 1
transform 1 0 3680 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2_2459
timestamp 1
transform 1 0 106628 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_1_1848
timestamp 1
transform 1 0 6256 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_1_1849
timestamp 1
transform 1 0 3680 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2_2460
timestamp 1
transform 1 0 106628 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_183_1_1850
timestamp 1
transform 1 0 6256 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_184_1_1851
timestamp 1
transform 1 0 3680 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_184_2_2461
timestamp 1
transform 1 0 106628 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_185_1_1852
timestamp 1
transform 1 0 6256 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_186_1_1853
timestamp 1
transform 1 0 3680 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_186_2_2462
timestamp 1
transform 1 0 106628 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_187_1_1854
timestamp 1
transform 1 0 6256 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_188_1_1855
timestamp 1
transform 1 0 3680 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_188_2_2463
timestamp 1
transform 1 0 106628 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_189_1_1856
timestamp 1
transform 1 0 6256 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_190_1_1857
timestamp 1
transform 1 0 3680 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_190_2_2464
timestamp 1
transform 1 0 106628 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_191_1_1858
timestamp 1
transform 1 0 6256 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_192_1_1859
timestamp 1
transform 1 0 3680 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_192_2_2465
timestamp 1
transform 1 0 106628 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_193_1_1860
timestamp 1
transform 1 0 6256 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_194_1_1861
timestamp 1
transform 1 0 3680 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_194_2_2466
timestamp 1
transform 1 0 106628 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_195_1_1862
timestamp 1
transform 1 0 6256 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_196_1_1863
timestamp 1
transform 1 0 3680 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_196_2_2467
timestamp 1
transform 1 0 106628 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_197_1_1864
timestamp 1
transform 1 0 6256 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_198_1_1865
timestamp 1
transform 1 0 3680 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_198_2_2468
timestamp 1
transform 1 0 106628 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_199_1_1866
timestamp 1
transform 1 0 6256 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_200_1_1867
timestamp 1
transform 1 0 3680 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_200_2_2469
timestamp 1
transform 1 0 106628 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_201_1_1868
timestamp 1
transform 1 0 6256 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_202_1_1869
timestamp 1
transform 1 0 3680 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_202_2_2470
timestamp 1
transform 1 0 106628 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_203_1_1870
timestamp 1
transform 1 0 6256 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_204_1_1871
timestamp 1
transform 1 0 3680 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_204_2_2471
timestamp 1
transform 1 0 106628 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_205_1_1872
timestamp 1
transform 1 0 6256 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_206_1_1873
timestamp 1
transform 1 0 3680 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_206_2_2472
timestamp 1
transform 1 0 106628 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_207_1_1874
timestamp 1
transform 1 0 6256 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_208_1_1875
timestamp 1
transform 1 0 3680 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_208_2_2473
timestamp 1
transform 1 0 106628 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_209_1_1876
timestamp 1
transform 1 0 6256 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_210_1_1877
timestamp 1
transform 1 0 3680 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_210_2_2474
timestamp 1
transform 1 0 106628 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_211_1_1878
timestamp 1
transform 1 0 6256 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_212_1_1879
timestamp 1
transform 1 0 3680 0 1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_212_2_2475
timestamp 1
transform 1 0 106628 0 1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_213_1_1880
timestamp 1
transform 1 0 6256 0 -1 118592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_214_1_1881
timestamp 1
transform 1 0 3680 0 1 118592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_214_2_2476
timestamp 1
transform 1 0 106628 0 1 118592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_215_1_1882
timestamp 1
transform 1 0 6256 0 -1 119680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_216_1_1883
timestamp 1
transform 1 0 3680 0 1 119680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_216_2_2477
timestamp 1
transform 1 0 106628 0 1 119680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_217_1_1884
timestamp 1
transform 1 0 6256 0 -1 120768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_218_1_1885
timestamp 1
transform 1 0 3680 0 1 120768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_218_2_2478
timestamp 1
transform 1 0 106628 0 1 120768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_219_1_1886
timestamp 1
transform 1 0 6256 0 -1 121856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_220_1_1887
timestamp 1
transform 1 0 3680 0 1 121856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_220_2_2479
timestamp 1
transform 1 0 106628 0 1 121856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_221_1_1888
timestamp 1
transform 1 0 6256 0 -1 122944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_222_1_1889
timestamp 1
transform 1 0 3680 0 1 122944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_222_2_2480
timestamp 1
transform 1 0 106628 0 1 122944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_223_1_1890
timestamp 1
transform 1 0 6256 0 -1 124032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_224_1_1891
timestamp 1
transform 1 0 3680 0 1 124032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_224_2_2481
timestamp 1
transform 1 0 106628 0 1 124032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_225_1_1892
timestamp 1
transform 1 0 6256 0 -1 125120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_226_1_1893
timestamp 1
transform 1 0 3680 0 1 125120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_226_2_2482
timestamp 1
transform 1 0 106628 0 1 125120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_227_1_1894
timestamp 1
transform 1 0 6256 0 -1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1_1895
timestamp 1
transform 1 0 3680 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_2_2483
timestamp 1
transform 1 0 106628 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1_1896
timestamp 1
transform 1 0 6256 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_230_1_1897
timestamp 1
transform 1 0 3680 0 1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_230_2_2484
timestamp 1
transform 1 0 106628 0 1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_231_1_1898
timestamp 1
transform 1 0 6256 0 -1 128384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_232_1_1899
timestamp 1
transform 1 0 3680 0 1 128384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_232_2_2485
timestamp 1
transform 1 0 106628 0 1 128384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_233_1_1900
timestamp 1
transform 1 0 6256 0 -1 129472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_234_1_1901
timestamp 1
transform 1 0 3680 0 1 129472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_234_2_2486
timestamp 1
transform 1 0 106628 0 1 129472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_235_1_1902
timestamp 1
transform 1 0 6256 0 -1 130560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_236_1_1903
timestamp 1
transform 1 0 3680 0 1 130560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_236_2_2487
timestamp 1
transform 1 0 106628 0 1 130560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_237_1_1904
timestamp 1
transform 1 0 6256 0 -1 131648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_238_1_1905
timestamp 1
transform 1 0 3680 0 1 131648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_238_2_2488
timestamp 1
transform 1 0 106628 0 1 131648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_239_1_1906
timestamp 1
transform 1 0 6256 0 -1 132736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_240_1_1907
timestamp 1
transform 1 0 3680 0 1 132736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_240_2_2489
timestamp 1
transform 1 0 106628 0 1 132736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_241_1_1908
timestamp 1
transform 1 0 6256 0 -1 133824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_242_1_1909
timestamp 1
transform 1 0 3680 0 1 133824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_242_2_2490
timestamp 1
transform 1 0 106628 0 1 133824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_243_1_1910
timestamp 1
transform 1 0 6256 0 -1 134912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_244_1_1911
timestamp 1
transform 1 0 3680 0 1 134912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_244_2_2491
timestamp 1
transform 1 0 106628 0 1 134912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_245_1_1912
timestamp 1
transform 1 0 6256 0 -1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1913
timestamp 1
transform 1 0 3680 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1914
timestamp 1
transform 1 0 6256 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1915
timestamp 1
transform 1 0 8832 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1916
timestamp 1
transform 1 0 11408 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1917
timestamp 1
transform 1 0 13984 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1918
timestamp 1
transform 1 0 16560 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1919
timestamp 1
transform 1 0 19136 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1920
timestamp 1
transform 1 0 21712 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1921
timestamp 1
transform 1 0 24288 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1922
timestamp 1
transform 1 0 26864 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1923
timestamp 1
transform 1 0 29440 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1924
timestamp 1
transform 1 0 32016 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1925
timestamp 1
transform 1 0 34592 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1926
timestamp 1
transform 1 0 37168 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1927
timestamp 1
transform 1 0 39744 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1928
timestamp 1
transform 1 0 42320 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1929
timestamp 1
transform 1 0 44896 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1930
timestamp 1
transform 1 0 47472 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1931
timestamp 1
transform 1 0 50048 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1932
timestamp 1
transform 1 0 52624 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1933
timestamp 1
transform 1 0 55200 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1934
timestamp 1
transform 1 0 57776 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1935
timestamp 1
transform 1 0 60352 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1936
timestamp 1
transform 1 0 62928 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1937
timestamp 1
transform 1 0 65504 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1938
timestamp 1
transform 1 0 68080 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1939
timestamp 1
transform 1 0 70656 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1940
timestamp 1
transform 1 0 73232 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1941
timestamp 1
transform 1 0 75808 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1942
timestamp 1
transform 1 0 78384 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1943
timestamp 1
transform 1 0 80960 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1944
timestamp 1
transform 1 0 83536 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1945
timestamp 1
transform 1 0 86112 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1946
timestamp 1
transform 1 0 88688 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1947
timestamp 1
transform 1 0 91264 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1948
timestamp 1
transform 1 0 93840 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1949
timestamp 1
transform 1 0 96416 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1950
timestamp 1
transform 1 0 98992 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1951
timestamp 1
transform 1 0 101568 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1952
timestamp 1
transform 1 0 104144 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1953
timestamp 1
transform 1 0 106720 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1954
timestamp 1
transform 1 0 6256 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1955
timestamp 1
transform 1 0 11408 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1956
timestamp 1
transform 1 0 16560 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1957
timestamp 1
transform 1 0 21712 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1958
timestamp 1
transform 1 0 26864 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1959
timestamp 1
transform 1 0 32016 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1960
timestamp 1
transform 1 0 37168 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1961
timestamp 1
transform 1 0 42320 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1962
timestamp 1
transform 1 0 47472 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1963
timestamp 1
transform 1 0 52624 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1964
timestamp 1
transform 1 0 57776 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1965
timestamp 1
transform 1 0 62928 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1966
timestamp 1
transform 1 0 68080 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1967
timestamp 1
transform 1 0 73232 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1968
timestamp 1
transform 1 0 78384 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1969
timestamp 1
transform 1 0 83536 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1970
timestamp 1
transform 1 0 88688 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1971
timestamp 1
transform 1 0 93840 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1972
timestamp 1
transform 1 0 98992 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1973
timestamp 1
transform 1 0 104144 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1974
timestamp 1
transform 1 0 3680 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1975
timestamp 1
transform 1 0 8832 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1976
timestamp 1
transform 1 0 13984 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1977
timestamp 1
transform 1 0 19136 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1978
timestamp 1
transform 1 0 24288 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1979
timestamp 1
transform 1 0 29440 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1980
timestamp 1
transform 1 0 34592 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1981
timestamp 1
transform 1 0 39744 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1982
timestamp 1
transform 1 0 44896 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1983
timestamp 1
transform 1 0 50048 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1984
timestamp 1
transform 1 0 55200 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1985
timestamp 1
transform 1 0 60352 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1986
timestamp 1
transform 1 0 65504 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1987
timestamp 1
transform 1 0 70656 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1988
timestamp 1
transform 1 0 75808 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1989
timestamp 1
transform 1 0 80960 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1990
timestamp 1
transform 1 0 86112 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1991
timestamp 1
transform 1 0 91264 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1992
timestamp 1
transform 1 0 96416 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1993
timestamp 1
transform 1 0 101568 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1994
timestamp 1
transform 1 0 106720 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_1995
timestamp 1
transform 1 0 6256 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_1996
timestamp 1
transform 1 0 11408 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_1997
timestamp 1
transform 1 0 16560 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_1998
timestamp 1
transform 1 0 21712 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_1999
timestamp 1
transform 1 0 26864 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2000
timestamp 1
transform 1 0 32016 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2001
timestamp 1
transform 1 0 37168 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2002
timestamp 1
transform 1 0 42320 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2003
timestamp 1
transform 1 0 47472 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2004
timestamp 1
transform 1 0 52624 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2005
timestamp 1
transform 1 0 57776 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2006
timestamp 1
transform 1 0 62928 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2007
timestamp 1
transform 1 0 68080 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2008
timestamp 1
transform 1 0 73232 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2009
timestamp 1
transform 1 0 78384 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2010
timestamp 1
transform 1 0 83536 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2011
timestamp 1
transform 1 0 88688 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2012
timestamp 1
transform 1 0 93840 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2013
timestamp 1
transform 1 0 98992 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2014
timestamp 1
transform 1 0 104144 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2015
timestamp 1
transform 1 0 3680 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2016
timestamp 1
transform 1 0 8832 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2017
timestamp 1
transform 1 0 13984 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2018
timestamp 1
transform 1 0 19136 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2019
timestamp 1
transform 1 0 24288 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2020
timestamp 1
transform 1 0 29440 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2021
timestamp 1
transform 1 0 34592 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2022
timestamp 1
transform 1 0 39744 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2023
timestamp 1
transform 1 0 44896 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2024
timestamp 1
transform 1 0 50048 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2025
timestamp 1
transform 1 0 55200 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2026
timestamp 1
transform 1 0 60352 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2027
timestamp 1
transform 1 0 65504 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2028
timestamp 1
transform 1 0 70656 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2029
timestamp 1
transform 1 0 75808 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2030
timestamp 1
transform 1 0 80960 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2031
timestamp 1
transform 1 0 86112 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2032
timestamp 1
transform 1 0 91264 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2033
timestamp 1
transform 1 0 96416 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2034
timestamp 1
transform 1 0 101568 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2035
timestamp 1
transform 1 0 106720 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2036
timestamp 1
transform 1 0 6256 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2037
timestamp 1
transform 1 0 11408 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2038
timestamp 1
transform 1 0 16560 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2039
timestamp 1
transform 1 0 21712 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2040
timestamp 1
transform 1 0 26864 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2041
timestamp 1
transform 1 0 32016 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2042
timestamp 1
transform 1 0 37168 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2043
timestamp 1
transform 1 0 42320 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2044
timestamp 1
transform 1 0 47472 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2045
timestamp 1
transform 1 0 52624 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2046
timestamp 1
transform 1 0 57776 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2047
timestamp 1
transform 1 0 62928 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2048
timestamp 1
transform 1 0 68080 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2049
timestamp 1
transform 1 0 73232 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2050
timestamp 1
transform 1 0 78384 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2051
timestamp 1
transform 1 0 83536 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2052
timestamp 1
transform 1 0 88688 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2053
timestamp 1
transform 1 0 93840 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2054
timestamp 1
transform 1 0 98992 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2055
timestamp 1
transform 1 0 104144 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2056
timestamp 1
transform 1 0 3680 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2057
timestamp 1
transform 1 0 8832 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2058
timestamp 1
transform 1 0 13984 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2059
timestamp 1
transform 1 0 19136 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2060
timestamp 1
transform 1 0 24288 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2061
timestamp 1
transform 1 0 29440 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2062
timestamp 1
transform 1 0 34592 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2063
timestamp 1
transform 1 0 39744 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2064
timestamp 1
transform 1 0 44896 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2065
timestamp 1
transform 1 0 50048 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2066
timestamp 1
transform 1 0 55200 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2067
timestamp 1
transform 1 0 60352 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2068
timestamp 1
transform 1 0 65504 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2069
timestamp 1
transform 1 0 70656 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2070
timestamp 1
transform 1 0 75808 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2071
timestamp 1
transform 1 0 80960 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2072
timestamp 1
transform 1 0 86112 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2073
timestamp 1
transform 1 0 91264 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2074
timestamp 1
transform 1 0 96416 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2075
timestamp 1
transform 1 0 101568 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2076
timestamp 1
transform 1 0 106720 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2077
timestamp 1
transform 1 0 6256 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2078
timestamp 1
transform 1 0 11408 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2079
timestamp 1
transform 1 0 16560 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2080
timestamp 1
transform 1 0 21712 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2081
timestamp 1
transform 1 0 26864 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2082
timestamp 1
transform 1 0 32016 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2083
timestamp 1
transform 1 0 37168 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2084
timestamp 1
transform 1 0 42320 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2085
timestamp 1
transform 1 0 47472 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2086
timestamp 1
transform 1 0 52624 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2087
timestamp 1
transform 1 0 57776 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2088
timestamp 1
transform 1 0 62928 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2089
timestamp 1
transform 1 0 68080 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2090
timestamp 1
transform 1 0 73232 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2091
timestamp 1
transform 1 0 78384 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2092
timestamp 1
transform 1 0 83536 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2093
timestamp 1
transform 1 0 88688 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2094
timestamp 1
transform 1 0 93840 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2095
timestamp 1
transform 1 0 98992 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2096
timestamp 1
transform 1 0 104144 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2097
timestamp 1
transform 1 0 3680 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2098
timestamp 1
transform 1 0 8832 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2099
timestamp 1
transform 1 0 13984 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2100
timestamp 1
transform 1 0 19136 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2101
timestamp 1
transform 1 0 24288 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2102
timestamp 1
transform 1 0 29440 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2103
timestamp 1
transform 1 0 34592 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2104
timestamp 1
transform 1 0 39744 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2105
timestamp 1
transform 1 0 44896 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2106
timestamp 1
transform 1 0 50048 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2107
timestamp 1
transform 1 0 55200 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2108
timestamp 1
transform 1 0 60352 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2109
timestamp 1
transform 1 0 65504 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2110
timestamp 1
transform 1 0 70656 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2111
timestamp 1
transform 1 0 75808 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2112
timestamp 1
transform 1 0 80960 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2113
timestamp 1
transform 1 0 86112 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2114
timestamp 1
transform 1 0 91264 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2115
timestamp 1
transform 1 0 96416 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2116
timestamp 1
transform 1 0 101568 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2117
timestamp 1
transform 1 0 106720 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2118
timestamp 1
transform 1 0 6256 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2119
timestamp 1
transform 1 0 11408 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2120
timestamp 1
transform 1 0 16560 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2121
timestamp 1
transform 1 0 21712 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2122
timestamp 1
transform 1 0 26864 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2123
timestamp 1
transform 1 0 32016 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2124
timestamp 1
transform 1 0 37168 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2125
timestamp 1
transform 1 0 42320 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2126
timestamp 1
transform 1 0 47472 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2127
timestamp 1
transform 1 0 52624 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2128
timestamp 1
transform 1 0 57776 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2129
timestamp 1
transform 1 0 62928 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2130
timestamp 1
transform 1 0 68080 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2131
timestamp 1
transform 1 0 73232 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2132
timestamp 1
transform 1 0 78384 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2133
timestamp 1
transform 1 0 83536 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2134
timestamp 1
transform 1 0 88688 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2135
timestamp 1
transform 1 0 93840 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2136
timestamp 1
transform 1 0 98992 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2137
timestamp 1
transform 1 0 104144 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2138
timestamp 1
transform 1 0 3680 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2139
timestamp 1
transform 1 0 8832 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2140
timestamp 1
transform 1 0 13984 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2141
timestamp 1
transform 1 0 19136 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2142
timestamp 1
transform 1 0 24288 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2143
timestamp 1
transform 1 0 29440 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2144
timestamp 1
transform 1 0 34592 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2145
timestamp 1
transform 1 0 39744 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2146
timestamp 1
transform 1 0 44896 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2147
timestamp 1
transform 1 0 50048 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2148
timestamp 1
transform 1 0 55200 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2149
timestamp 1
transform 1 0 60352 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2150
timestamp 1
transform 1 0 65504 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2151
timestamp 1
transform 1 0 70656 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2152
timestamp 1
transform 1 0 75808 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2153
timestamp 1
transform 1 0 80960 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2154
timestamp 1
transform 1 0 86112 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2155
timestamp 1
transform 1 0 91264 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2156
timestamp 1
transform 1 0 96416 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2157
timestamp 1
transform 1 0 101568 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2158
timestamp 1
transform 1 0 106720 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2159
timestamp 1
transform 1 0 6256 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2160
timestamp 1
transform 1 0 11408 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2161
timestamp 1
transform 1 0 16560 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2162
timestamp 1
transform 1 0 21712 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2163
timestamp 1
transform 1 0 26864 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2164
timestamp 1
transform 1 0 32016 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2165
timestamp 1
transform 1 0 37168 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2166
timestamp 1
transform 1 0 42320 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2167
timestamp 1
transform 1 0 47472 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2168
timestamp 1
transform 1 0 52624 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2169
timestamp 1
transform 1 0 57776 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2170
timestamp 1
transform 1 0 62928 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2171
timestamp 1
transform 1 0 68080 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2172
timestamp 1
transform 1 0 73232 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2173
timestamp 1
transform 1 0 78384 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2174
timestamp 1
transform 1 0 83536 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2175
timestamp 1
transform 1 0 88688 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2176
timestamp 1
transform 1 0 93840 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2177
timestamp 1
transform 1 0 98992 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2178
timestamp 1
transform 1 0 104144 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2179
timestamp 1
transform 1 0 3680 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2180
timestamp 1
transform 1 0 8832 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2181
timestamp 1
transform 1 0 13984 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2182
timestamp 1
transform 1 0 19136 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2183
timestamp 1
transform 1 0 24288 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2184
timestamp 1
transform 1 0 29440 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2185
timestamp 1
transform 1 0 34592 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2186
timestamp 1
transform 1 0 39744 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2187
timestamp 1
transform 1 0 44896 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2188
timestamp 1
transform 1 0 50048 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2189
timestamp 1
transform 1 0 55200 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2190
timestamp 1
transform 1 0 60352 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2191
timestamp 1
transform 1 0 65504 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2192
timestamp 1
transform 1 0 70656 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2193
timestamp 1
transform 1 0 75808 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2194
timestamp 1
transform 1 0 80960 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2195
timestamp 1
transform 1 0 86112 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2196
timestamp 1
transform 1 0 91264 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2197
timestamp 1
transform 1 0 96416 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2198
timestamp 1
transform 1 0 101568 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2199
timestamp 1
transform 1 0 106720 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2200
timestamp 1
transform 1 0 6256 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2201
timestamp 1
transform 1 0 11408 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2202
timestamp 1
transform 1 0 16560 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2203
timestamp 1
transform 1 0 21712 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2204
timestamp 1
transform 1 0 26864 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2205
timestamp 1
transform 1 0 32016 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2206
timestamp 1
transform 1 0 37168 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2207
timestamp 1
transform 1 0 42320 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2208
timestamp 1
transform 1 0 47472 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2209
timestamp 1
transform 1 0 52624 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2210
timestamp 1
transform 1 0 57776 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2211
timestamp 1
transform 1 0 62928 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2212
timestamp 1
transform 1 0 68080 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2213
timestamp 1
transform 1 0 73232 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2214
timestamp 1
transform 1 0 78384 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2215
timestamp 1
transform 1 0 83536 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2216
timestamp 1
transform 1 0 88688 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2217
timestamp 1
transform 1 0 93840 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2218
timestamp 1
transform 1 0 98992 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2219
timestamp 1
transform 1 0 104144 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2220
timestamp 1
transform 1 0 3680 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2221
timestamp 1
transform 1 0 8832 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2222
timestamp 1
transform 1 0 13984 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2223
timestamp 1
transform 1 0 19136 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2224
timestamp 1
transform 1 0 24288 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2225
timestamp 1
transform 1 0 29440 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2226
timestamp 1
transform 1 0 34592 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2227
timestamp 1
transform 1 0 39744 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2228
timestamp 1
transform 1 0 44896 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2229
timestamp 1
transform 1 0 50048 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2230
timestamp 1
transform 1 0 55200 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2231
timestamp 1
transform 1 0 60352 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2232
timestamp 1
transform 1 0 65504 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2233
timestamp 1
transform 1 0 70656 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2234
timestamp 1
transform 1 0 75808 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2235
timestamp 1
transform 1 0 80960 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2236
timestamp 1
transform 1 0 86112 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2237
timestamp 1
transform 1 0 91264 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2238
timestamp 1
transform 1 0 96416 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2239
timestamp 1
transform 1 0 101568 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2240
timestamp 1
transform 1 0 106720 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2241
timestamp 1
transform 1 0 6256 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2242
timestamp 1
transform 1 0 11408 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2243
timestamp 1
transform 1 0 16560 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2244
timestamp 1
transform 1 0 21712 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2245
timestamp 1
transform 1 0 26864 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2246
timestamp 1
transform 1 0 32016 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2247
timestamp 1
transform 1 0 37168 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2248
timestamp 1
transform 1 0 42320 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2249
timestamp 1
transform 1 0 47472 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2250
timestamp 1
transform 1 0 52624 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2251
timestamp 1
transform 1 0 57776 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2252
timestamp 1
transform 1 0 62928 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2253
timestamp 1
transform 1 0 68080 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2254
timestamp 1
transform 1 0 73232 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2255
timestamp 1
transform 1 0 78384 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2256
timestamp 1
transform 1 0 83536 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2257
timestamp 1
transform 1 0 88688 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2258
timestamp 1
transform 1 0 93840 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2259
timestamp 1
transform 1 0 98992 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2260
timestamp 1
transform 1 0 104144 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2261
timestamp 1
transform 1 0 3680 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2262
timestamp 1
transform 1 0 8832 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2263
timestamp 1
transform 1 0 13984 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2264
timestamp 1
transform 1 0 19136 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2265
timestamp 1
transform 1 0 24288 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2266
timestamp 1
transform 1 0 29440 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2267
timestamp 1
transform 1 0 34592 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2268
timestamp 1
transform 1 0 39744 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2269
timestamp 1
transform 1 0 44896 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2270
timestamp 1
transform 1 0 50048 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2271
timestamp 1
transform 1 0 55200 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2272
timestamp 1
transform 1 0 60352 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2273
timestamp 1
transform 1 0 65504 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2274
timestamp 1
transform 1 0 70656 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2275
timestamp 1
transform 1 0 75808 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2276
timestamp 1
transform 1 0 80960 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2277
timestamp 1
transform 1 0 86112 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2278
timestamp 1
transform 1 0 91264 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2279
timestamp 1
transform 1 0 96416 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2280
timestamp 1
transform 1 0 101568 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2281
timestamp 1
transform 1 0 106720 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2282
timestamp 1
transform 1 0 6256 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2283
timestamp 1
transform 1 0 11408 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2284
timestamp 1
transform 1 0 16560 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2285
timestamp 1
transform 1 0 21712 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2286
timestamp 1
transform 1 0 26864 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2287
timestamp 1
transform 1 0 32016 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2288
timestamp 1
transform 1 0 37168 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2289
timestamp 1
transform 1 0 42320 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2290
timestamp 1
transform 1 0 47472 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2291
timestamp 1
transform 1 0 52624 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2292
timestamp 1
transform 1 0 57776 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2293
timestamp 1
transform 1 0 62928 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2294
timestamp 1
transform 1 0 68080 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2295
timestamp 1
transform 1 0 73232 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2296
timestamp 1
transform 1 0 78384 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2297
timestamp 1
transform 1 0 83536 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2298
timestamp 1
transform 1 0 88688 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2299
timestamp 1
transform 1 0 93840 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2300
timestamp 1
transform 1 0 98992 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2301
timestamp 1
transform 1 0 104144 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2302
timestamp 1
transform 1 0 3680 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2303
timestamp 1
transform 1 0 8832 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2304
timestamp 1
transform 1 0 13984 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2305
timestamp 1
transform 1 0 19136 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2306
timestamp 1
transform 1 0 24288 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2307
timestamp 1
transform 1 0 29440 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2308
timestamp 1
transform 1 0 34592 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2309
timestamp 1
transform 1 0 39744 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2310
timestamp 1
transform 1 0 44896 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2311
timestamp 1
transform 1 0 50048 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2312
timestamp 1
transform 1 0 55200 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2313
timestamp 1
transform 1 0 60352 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2314
timestamp 1
transform 1 0 65504 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2315
timestamp 1
transform 1 0 70656 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2316
timestamp 1
transform 1 0 75808 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2317
timestamp 1
transform 1 0 80960 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2318
timestamp 1
transform 1 0 86112 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2319
timestamp 1
transform 1 0 91264 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2320
timestamp 1
transform 1 0 96416 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2321
timestamp 1
transform 1 0 101568 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2322
timestamp 1
transform 1 0 106720 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2323
timestamp 1
transform 1 0 6256 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2324
timestamp 1
transform 1 0 11408 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2325
timestamp 1
transform 1 0 16560 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2326
timestamp 1
transform 1 0 21712 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2327
timestamp 1
transform 1 0 26864 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2328
timestamp 1
transform 1 0 32016 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2329
timestamp 1
transform 1 0 37168 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2330
timestamp 1
transform 1 0 42320 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2331
timestamp 1
transform 1 0 47472 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2332
timestamp 1
transform 1 0 52624 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2333
timestamp 1
transform 1 0 57776 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2334
timestamp 1
transform 1 0 62928 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2335
timestamp 1
transform 1 0 68080 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2336
timestamp 1
transform 1 0 73232 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2337
timestamp 1
transform 1 0 78384 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2338
timestamp 1
transform 1 0 83536 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2339
timestamp 1
transform 1 0 88688 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2340
timestamp 1
transform 1 0 93840 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2341
timestamp 1
transform 1 0 98992 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2342
timestamp 1
transform 1 0 104144 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2343
timestamp 1
transform 1 0 3680 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2344
timestamp 1
transform 1 0 6256 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2345
timestamp 1
transform 1 0 8832 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2346
timestamp 1
transform 1 0 11408 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2347
timestamp 1
transform 1 0 13984 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2348
timestamp 1
transform 1 0 16560 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2349
timestamp 1
transform 1 0 19136 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2350
timestamp 1
transform 1 0 21712 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2351
timestamp 1
transform 1 0 24288 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2352
timestamp 1
transform 1 0 26864 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2353
timestamp 1
transform 1 0 29440 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2354
timestamp 1
transform 1 0 32016 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2355
timestamp 1
transform 1 0 34592 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2356
timestamp 1
transform 1 0 37168 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2357
timestamp 1
transform 1 0 39744 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2358
timestamp 1
transform 1 0 42320 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2359
timestamp 1
transform 1 0 44896 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2360
timestamp 1
transform 1 0 47472 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2361
timestamp 1
transform 1 0 50048 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2362
timestamp 1
transform 1 0 52624 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2363
timestamp 1
transform 1 0 55200 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2364
timestamp 1
transform 1 0 57776 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2365
timestamp 1
transform 1 0 60352 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2366
timestamp 1
transform 1 0 62928 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2367
timestamp 1
transform 1 0 65504 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2368
timestamp 1
transform 1 0 68080 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2369
timestamp 1
transform 1 0 70656 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2370
timestamp 1
transform 1 0 73232 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2371
timestamp 1
transform 1 0 75808 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2372
timestamp 1
transform 1 0 78384 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2373
timestamp 1
transform 1 0 80960 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2374
timestamp 1
transform 1 0 83536 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2375
timestamp 1
transform 1 0 86112 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2376
timestamp 1
transform 1 0 88688 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2377
timestamp 1
transform 1 0 91264 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2378
timestamp 1
transform 1 0 93840 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2379
timestamp 1
transform 1 0 96416 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2380
timestamp 1
transform 1 0 98992 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2381
timestamp 1
transform 1 0 101568 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2382
timestamp 1
transform 1 0 104144 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2383
timestamp 1
transform 1 0 106720 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  wire68
timestamp 1
transform 1 0 60536 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire69
timestamp 1
transform 1 0 58052 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire70
timestamp 1
transform 1 0 55660 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire71
timestamp 1
transform 1 0 53452 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire72
timestamp 1
transform -1 0 47932 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire73
timestamp 1
transform -1 0 45448 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire74
timestamp 1
transform -1 0 43148 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire75
timestamp 1
transform -1 0 40848 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire76
timestamp 1
transform -1 0 38364 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire77
timestamp 1
transform 1 0 74060 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire78
timestamp 1
transform 1 0 72036 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire79
timestamp 1
transform 1 0 69644 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire80
timestamp 1
transform 1 0 67436 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire81
timestamp 1
transform 1 0 64860 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire82
timestamp 1
transform 1 0 63020 0 1 136000
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 addr00[0]
port 0 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 addr00[1]
port 1 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 addr00[2]
port 2 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 addr00[3]
port 3 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 addr00[4]
port 4 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 addr00[5]
port 5 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 addr00[6]
port 6 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 addr00[7]
port 7 nsew signal input
flabel metal3 s 0 88408 800 88528 0 FreeSans 480 0 0 0 addr01[0]
port 8 nsew signal input
flabel metal3 s 0 80248 800 80368 0 FreeSans 480 0 0 0 addr01[1]
port 9 nsew signal input
flabel metal3 s 0 104048 800 104168 0 FreeSans 480 0 0 0 addr01[2]
port 10 nsew signal input
flabel metal3 s 0 105408 800 105528 0 FreeSans 480 0 0 0 addr01[3]
port 11 nsew signal input
flabel metal3 s 0 106768 800 106888 0 FreeSans 480 0 0 0 addr01[4]
port 12 nsew signal input
flabel metal3 s 0 108128 800 108248 0 FreeSans 480 0 0 0 addr01[5]
port 13 nsew signal input
flabel metal3 s 0 109488 800 109608 0 FreeSans 480 0 0 0 addr01[6]
port 14 nsew signal input
flabel metal3 s 0 110848 800 110968 0 FreeSans 480 0 0 0 addr01[7]
port 15 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 clk
port 16 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 csb00
port 17 nsew signal input
flabel metal3 s 0 85688 800 85808 0 FreeSans 480 0 0 0 csb01
port 18 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 din00[0]
port 19 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 din00[10]
port 20 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 din00[11]
port 21 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 din00[12]
port 22 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 din00[13]
port 23 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 din00[14]
port 24 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 din00[15]
port 25 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 din00[1]
port 26 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 din00[2]
port 27 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 din00[3]
port 28 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 din00[4]
port 29 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 din00[5]
port 30 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 din00[6]
port 31 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 din00[7]
port 32 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 din00[8]
port 33 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 din00[9]
port 34 nsew signal input
flabel metal3 s 0 80928 800 81048 0 FreeSans 480 0 0 0 din01[0]
port 35 nsew signal input
flabel metal3 s 0 79568 800 79688 0 FreeSans 480 0 0 0 din01[10]
port 36 nsew signal input
flabel metal3 s 0 81608 800 81728 0 FreeSans 480 0 0 0 din01[11]
port 37 nsew signal input
flabel metal3 s 0 82288 800 82408 0 FreeSans 480 0 0 0 din01[12]
port 38 nsew signal input
flabel metal3 s 0 82968 800 83088 0 FreeSans 480 0 0 0 din01[13]
port 39 nsew signal input
flabel metal3 s 0 78888 800 79008 0 FreeSans 480 0 0 0 din01[14]
port 40 nsew signal input
flabel metal3 s 0 76848 800 76968 0 FreeSans 480 0 0 0 din01[15]
port 41 nsew signal input
flabel metal3 s 0 84328 800 84448 0 FreeSans 480 0 0 0 din01[1]
port 42 nsew signal input
flabel metal3 s 0 72088 800 72208 0 FreeSans 480 0 0 0 din01[2]
port 43 nsew signal input
flabel metal3 s 0 78208 800 78328 0 FreeSans 480 0 0 0 din01[3]
port 44 nsew signal input
flabel metal3 s 0 86368 800 86488 0 FreeSans 480 0 0 0 din01[4]
port 45 nsew signal input
flabel metal3 s 0 83648 800 83768 0 FreeSans 480 0 0 0 din01[5]
port 46 nsew signal input
flabel metal3 s 0 85008 800 85128 0 FreeSans 480 0 0 0 din01[6]
port 47 nsew signal input
flabel metal3 s 0 77528 800 77648 0 FreeSans 480 0 0 0 din01[7]
port 48 nsew signal input
flabel metal3 s 0 87048 800 87168 0 FreeSans 480 0 0 0 din01[8]
port 49 nsew signal input
flabel metal3 s 0 87728 800 87848 0 FreeSans 480 0 0 0 din01[9]
port 50 nsew signal input
flabel metal3 s 109200 67328 110000 67448 0 FreeSans 480 0 0 0 rst
port 51 nsew signal input
flabel metal3 s 0 76168 800 76288 0 FreeSans 480 0 0 0 sine_out[0]
port 52 nsew signal output
flabel metal3 s 109200 72768 110000 72888 0 FreeSans 480 0 0 0 sine_out[10]
port 53 nsew signal output
flabel metal3 s 109200 78888 110000 79008 0 FreeSans 480 0 0 0 sine_out[11]
port 54 nsew signal output
flabel metal3 s 109200 78208 110000 78328 0 FreeSans 480 0 0 0 sine_out[12]
port 55 nsew signal output
flabel metal3 s 109200 77528 110000 77648 0 FreeSans 480 0 0 0 sine_out[13]
port 56 nsew signal output
flabel metal3 s 109200 76168 110000 76288 0 FreeSans 480 0 0 0 sine_out[14]
port 57 nsew signal output
flabel metal3 s 109200 76848 110000 76968 0 FreeSans 480 0 0 0 sine_out[15]
port 58 nsew signal output
flabel metal3 s 0 72768 800 72888 0 FreeSans 480 0 0 0 sine_out[1]
port 59 nsew signal output
flabel metal3 s 0 73448 800 73568 0 FreeSans 480 0 0 0 sine_out[2]
port 60 nsew signal output
flabel metal3 s 0 74128 800 74248 0 FreeSans 480 0 0 0 sine_out[3]
port 61 nsew signal output
flabel metal3 s 0 74808 800 74928 0 FreeSans 480 0 0 0 sine_out[4]
port 62 nsew signal output
flabel metal3 s 0 75488 800 75608 0 FreeSans 480 0 0 0 sine_out[5]
port 63 nsew signal output
flabel metal3 s 109200 73448 110000 73568 0 FreeSans 480 0 0 0 sine_out[6]
port 64 nsew signal output
flabel metal3 s 109200 74128 110000 74248 0 FreeSans 480 0 0 0 sine_out[7]
port 65 nsew signal output
flabel metal3 s 109200 74808 110000 74928 0 FreeSans 480 0 0 0 sine_out[8]
port 66 nsew signal output
flabel metal3 s 109200 75488 110000 75608 0 FreeSans 480 0 0 0 sine_out[9]
port 67 nsew signal output
flabel metal4 s 4208 2128 4528 147472 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 34928 2128 35248 7880 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 34928 65650 35248 77880 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 34928 135650 35248 147472 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 65648 2128 65968 8064 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 65648 65776 65968 78064 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 65648 135834 65968 147472 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 96368 2128 96688 8064 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 96368 65650 96688 78064 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 96368 135650 96688 147472 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal5 s 1056 5346 108884 5666 0 FreeSans 2560 0 0 0 vccd1
port 68 nsew power bidirectional
flabel metal5 s 1056 35982 108884 36302 0 FreeSans 2560 0 0 0 vccd1
port 68 nsew power bidirectional
flabel metal5 s 1056 66618 108884 66938 0 FreeSans 2560 0 0 0 vccd1
port 68 nsew power bidirectional
flabel metal5 s 1056 97254 108884 97574 0 FreeSans 2560 0 0 0 vccd1
port 68 nsew power bidirectional
flabel metal5 s 1056 127890 108884 128210 0 FreeSans 2560 0 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 105916 7024 106236 66416 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 105916 77200 106236 136592 0 FreeSans 1920 90 0 0 vccd1
port 68 nsew power bidirectional
flabel metal5 s 4208 140940 108884 141260 0 FreeSans 2560 0 0 0 vccd1
port 68 nsew power bidirectional
flabel metal4 s 4868 2128 5188 147472 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 8064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 35588 65650 35908 78064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 35588 135650 35908 147472 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 66308 2128 66628 8064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 66308 65650 66628 78064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 66308 135650 66628 147472 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 97028 2128 97348 8064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 97028 65650 97348 78064 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 97028 135650 97348 147472 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal5 s 1056 6006 108884 6326 0 FreeSans 2560 0 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal5 s 1056 36642 108884 36962 0 FreeSans 2560 0 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal5 s 1056 67278 108884 67598 0 FreeSans 2560 0 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal5 s 1056 97914 108884 98234 0 FreeSans 2560 0 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal5 s 1056 128550 108884 128870 0 FreeSans 2560 0 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 106652 7024 106972 66416 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal4 s 106652 77200 106972 136592 0 FreeSans 1920 90 0 0 vssd1
port 69 nsew ground bidirectional
flabel metal5 s 4208 141620 108884 141940 0 FreeSans 2560 0 0 0 vssd1
port 69 nsew ground bidirectional
rlabel via4 101806 128050 101806 128050 0 vccd1
rlabel via4 101110 128710 101110 128710 0 vssd1
rlabel metal2 21298 77690 21298 77690 0 _000_
rlabel metal2 70426 77792 70426 77792 0 _001_
rlabel metal2 71990 78030 71990 78030 0 _002_
rlabel metal2 74474 77894 74474 77894 0 _003_
rlabel metal2 76682 78064 76682 78064 0 _004_
rlabel metal2 79258 78098 79258 78098 0 _005_
rlabel metal2 80914 77792 80914 77792 0 _006_
rlabel metal2 32706 76908 32706 76908 0 _007_
rlabel metal1 25254 78234 25254 78234 0 _008_
rlabel metal2 24334 76466 24334 76466 0 _009_
rlabel metal2 30498 76993 30498 76993 0 _010_
rlabel metal2 39974 77367 39974 77367 0 _011_
rlabel metal1 62652 77350 62652 77350 0 _012_
rlabel metal2 63986 77894 63986 77894 0 _013_
rlabel metal1 68954 77418 68954 77418 0 _014_
rlabel metal2 69138 77826 69138 77826 0 _015_
rlabel metal1 83536 77146 83536 77146 0 _016_
rlabel metal1 85974 77554 85974 77554 0 _017_
rlabel metal2 89010 72080 89010 72080 0 _018_
rlabel metal1 90298 67320 90298 67320 0 _019_
rlabel metal2 88918 66776 88918 66776 0 _020_
rlabel metal1 90160 66810 90160 66810 0 _021_
rlabel metal1 88550 65960 88550 65960 0 _022_
rlabel metal1 84778 66266 84778 66266 0 _023_
rlabel metal1 77326 70414 77326 70414 0 _024_
rlabel metal1 84403 75990 84403 75990 0 _025_
rlabel metal1 86296 75378 86296 75378 0 _026_
rlabel metal1 86894 75446 86894 75446 0 _027_
rlabel metal2 85790 76840 85790 76840 0 _028_
rlabel metal1 88964 76534 88964 76534 0 _029_
rlabel metal2 88550 76840 88550 76840 0 _030_
rlabel metal1 91264 76602 91264 76602 0 _031_
rlabel metal2 95266 77248 95266 77248 0 _032_
rlabel metal2 81558 77282 81558 77282 0 _033_
rlabel metal2 84318 77010 84318 77010 0 _034_
rlabel metal1 88550 70822 88550 70822 0 _035_
rlabel metal2 90758 67694 90758 67694 0 _036_
rlabel metal1 86848 68102 86848 68102 0 _037_
rlabel metal1 86710 67626 86710 67626 0 _038_
rlabel metal1 85054 67014 85054 67014 0 _039_
rlabel metal1 84134 67014 84134 67014 0 _040_
rlabel metal1 74152 72250 74152 72250 0 _041_
rlabel metal2 20838 77724 20838 77724 0 _042_
rlabel metal1 26135 76330 26135 76330 0 _043_
rlabel metal1 23874 77595 23874 77595 0 _044_
rlabel metal2 24794 76806 24794 76806 0 _045_
rlabel metal1 29532 76602 29532 76602 0 _046_
rlabel metal2 26082 77826 26082 77826 0 _047_
rlabel metal1 82570 75174 82570 75174 0 _048_
rlabel metal1 82800 76330 82800 76330 0 _049_
rlabel via1 90482 73134 90482 73134 0 _050_
rlabel metal1 90252 75718 90252 75718 0 _051_
rlabel metal1 90942 67728 90942 67728 0 _052_
rlabel metal2 91126 68170 91126 68170 0 _053_
rlabel metal1 91034 65926 91034 65926 0 _054_
rlabel viali 91037 66606 91037 66606 0 _055_
rlabel metal1 88918 66198 88918 66198 0 _056_
rlabel metal1 81788 70414 81788 70414 0 _057_
rlabel metal1 86066 65994 86066 65994 0 _058_
rlabel metal1 1426 5202 1426 5202 0 addr00[0]
rlabel metal2 1978 8143 1978 8143 0 addr00[1]
rlabel metal1 1426 10642 1426 10642 0 addr00[2]
rlabel metal1 1380 11730 1380 11730 0 addr00[3]
rlabel metal2 1518 12563 1518 12563 0 addr00[4]
rlabel metal1 1426 13226 1426 13226 0 addr00[5]
rlabel metal2 1518 10999 1518 10999 0 addr00[6]
rlabel metal2 1518 13787 1518 13787 0 addr00[7]
rlabel metal1 1426 88978 1426 88978 0 addr01[0]
rlabel metal1 1380 80342 1380 80342 0 addr01[1]
rlabel metal1 1380 104210 1380 104210 0 addr01[2]
rlabel metal1 1380 105774 1380 105774 0 addr01[3]
rlabel metal1 1334 106862 1334 106862 0 addr01[4]
rlabel metal1 1380 108562 1380 108562 0 addr01[5]
rlabel metal1 1380 109650 1380 109650 0 addr01[6]
rlabel metal1 1380 111214 1380 111214 0 addr01[7]
rlabel metal1 55982 71978 55982 71978 0 clk
rlabel metal1 44666 72760 44666 72760 0 clknet_0_clk
rlabel metal2 83674 76908 83674 76908 0 clknet_2_0__leaf_clk
rlabel metal1 94898 77554 94898 77554 0 clknet_2_1__leaf_clk
rlabel metal2 6854 60180 6854 60180 0 clknet_2_2__leaf_clk
rlabel metal2 24610 76772 24610 76772 0 clknet_2_3__leaf_clk
rlabel metal2 1426 5593 1426 5593 0 csb00
rlabel metal1 1380 86190 1380 86190 0 csb01
rlabel metal1 1380 6290 1380 6290 0 din00[0]
rlabel metal2 37398 1520 37398 1520 0 din00[10]
rlabel metal2 38686 1520 38686 1520 0 din00[11]
rlabel metal2 39974 1520 39974 1520 0 din00[12]
rlabel metal2 41262 1520 41262 1520 0 din00[13]
rlabel metal2 41906 1520 41906 1520 0 din00[14]
rlabel metal2 43194 1520 43194 1520 0 din00[15]
rlabel metal1 1426 8874 1426 8874 0 din00[1]
rlabel metal3 1004 6868 1004 6868 0 din00[2]
rlabel metal2 1518 9775 1518 9775 0 din00[3]
rlabel metal1 1426 7786 1426 7786 0 din00[4]
rlabel metal2 31602 1520 31602 1520 0 din00[5]
rlabel metal2 32890 1520 32890 1520 0 din00[6]
rlabel metal2 34178 1520 34178 1520 0 din00[7]
rlabel metal2 35466 1520 35466 1520 0 din00[8]
rlabel metal2 36110 1520 36110 1520 0 din00[9]
rlabel metal1 1426 81362 1426 81362 0 din01[0]
rlabel metal1 1380 79594 1380 79594 0 din01[10]
rlabel metal1 1380 81770 1380 81770 0 din01[11]
rlabel metal1 1380 82450 1380 82450 0 din01[12]
rlabel metal1 1426 83538 1426 83538 0 din01[13]
rlabel metal1 1426 79186 1426 79186 0 din01[14]
rlabel metal1 1380 77010 1380 77010 0 din01[15]
rlabel metal1 1426 84626 1426 84626 0 din01[1]
rlabel metal1 1334 72658 1334 72658 0 din01[2]
rlabel metal1 1426 78506 1426 78506 0 din01[3]
rlabel metal1 1426 86802 1426 86802 0 din01[4]
rlabel metal1 1426 83946 1426 83946 0 din01[5]
rlabel metal1 1380 85034 1380 85034 0 din01[6]
rlabel metal1 1426 78098 1426 78098 0 din01[7]
rlabel metal1 1380 87210 1380 87210 0 din01[8]
rlabel metal1 1380 87890 1380 87890 0 din01[9]
rlabel metal1 1794 5066 1794 5066 0 net1
rlabel metal1 4002 80614 4002 80614 0 net10
rlabel metal3 102095 95060 102095 95060 0 net100
rlabel via2 102279 25060 102279 25060 0 net101
rlabel metal1 90704 75174 90704 75174 0 net102
rlabel metal4 86174 63983 86174 63983 0 net103
rlabel metal2 102626 106012 102626 106012 0 net104
rlabel metal1 86848 75990 86848 75990 0 net105
rlabel metal2 102258 105230 102258 105230 0 net106
rlabel metal1 85790 77010 85790 77010 0 net107
rlabel metal1 89148 71910 89148 71910 0 net108
rlabel metal1 90850 75276 90850 75276 0 net109
rlabel metal2 8418 104023 8418 104023 0 net11
rlabel metal2 84042 77078 84042 77078 0 net110
rlabel metal1 85974 76398 85974 76398 0 net111
rlabel metal2 83950 76500 83950 76500 0 net112
rlabel metal1 31510 76398 31510 76398 0 net113
rlabel metal3 102279 59738 102279 59738 0 net114
rlabel metal3 102279 129738 102279 129738 0 net115
rlabel metal2 8418 105757 8418 105757 0 net12
rlabel metal2 8418 106845 8418 106845 0 net13
rlabel via2 8418 108443 8418 108443 0 net14
rlabel via2 8418 109531 8418 109531 0 net15
rlabel metal2 8418 111265 8418 111265 0 net16
rlabel metal1 1702 5882 1702 5882 0 net17
rlabel metal2 6026 85765 6026 85765 0 net18
rlabel metal1 1794 6154 1794 6154 0 net19
rlabel metal1 1978 8364 1978 8364 0 net2
rlabel metal4 37486 9934 37486 9934 0 net20
rlabel metal4 38654 9934 38654 9934 0 net21
rlabel metal1 40020 2618 40020 2618 0 net22
rlabel metal4 40990 9934 40990 9934 0 net23
rlabel metal4 42158 9934 42158 9934 0 net24
rlabel metal3 43401 8228 43401 8228 0 net25
rlabel metal1 1794 8874 1794 8874 0 net26
rlabel metal1 1794 7242 1794 7242 0 net27
rlabel metal1 1794 9962 1794 9962 0 net28
rlabel metal1 1794 7786 1794 7786 0 net29
rlabel metal1 1702 10778 1702 10778 0 net3
rlabel via3 31717 8228 31717 8228 0 net30
rlabel metal4 32814 9866 32814 9866 0 net31
rlabel metal4 33982 9866 33982 9866 0 net32
rlabel metal1 35512 2618 35512 2618 0 net33
rlabel metal4 36318 9934 36318 9934 0 net34
rlabel metal1 3726 81158 3726 81158 0 net35
rlabel metal1 1794 79594 1794 79594 0 net36
rlabel metal2 1886 81464 1886 81464 0 net37
rlabel metal1 2162 82246 2162 82246 0 net38
rlabel metal1 2208 83334 2208 83334 0 net39
rlabel metal1 1702 11866 1702 11866 0 net4
rlabel metal1 1794 79050 1794 79050 0 net40
rlabel metal1 1794 76874 1794 76874 0 net41
rlabel metal1 1748 84490 1748 84490 0 net42
rlabel metal1 1794 72522 1794 72522 0 net43
rlabel metal1 1794 78506 1794 78506 0 net44
rlabel metal1 1794 86666 1794 86666 0 net45
rlabel metal1 1794 83946 1794 83946 0 net46
rlabel metal2 1886 83485 1886 83485 0 net47
rlabel metal1 1794 77962 1794 77962 0 net48
rlabel metal2 1886 86632 1886 86632 0 net49
rlabel metal1 1748 12886 1748 12886 0 net5
rlabel metal1 1794 87754 1794 87754 0 net50
rlabel metal2 107962 68272 107962 68272 0 net51
rlabel metal1 1702 76398 1702 76398 0 net52
rlabel metal1 89654 75786 89654 75786 0 net53
rlabel metal2 88918 78064 88918 78064 0 net54
rlabel metal2 99682 77724 99682 77724 0 net55
rlabel metal1 91310 76874 91310 76874 0 net56
rlabel metal2 93150 77826 93150 77826 0 net57
rlabel metal1 99590 77520 99590 77520 0 net58
rlabel metal2 23506 76874 23506 76874 0 net59
rlabel metal1 1748 13498 1748 13498 0 net6
rlabel metal1 22816 77350 22816 77350 0 net60
rlabel metal1 23874 76534 23874 76534 0 net61
rlabel metal1 1702 75310 1702 75310 0 net62
rlabel metal1 2070 76058 2070 76058 0 net63
rlabel metal2 102166 74256 102166 74256 0 net64
rlabel metal1 85284 76262 85284 76262 0 net65
rlabel metal1 87722 75310 87722 75310 0 net66
rlabel metal1 87998 76296 87998 76296 0 net67
rlabel metal2 61042 135932 61042 135932 0 net68
rlabel metal2 58558 135966 58558 135966 0 net69
rlabel metal1 1748 11322 1748 11322 0 net7
rlabel metal2 63342 78013 63342 78013 0 net70
rlabel metal2 61134 78404 61134 78404 0 net71
rlabel metal2 42918 77469 42918 77469 0 net72
rlabel metal2 45218 136000 45218 136000 0 net73
rlabel metal2 42918 135966 42918 135966 0 net74
rlabel metal2 40618 135932 40618 135932 0 net75
rlabel metal2 38134 135898 38134 135898 0 net76
rlabel metal1 80454 77622 80454 77622 0 net77
rlabel metal2 78798 77979 78798 77979 0 net78
rlabel metal2 76222 77911 76222 77911 0 net79
rlabel metal1 2668 14042 2668 14042 0 net8
rlabel metal2 74014 77843 74014 77843 0 net80
rlabel metal2 70978 77843 70978 77843 0 net81
rlabel metal2 63526 135898 63526 135898 0 net82
rlabel metal1 61456 77554 61456 77554 0 net83
rlabel metal1 75072 77486 75072 77486 0 net84
rlabel metal4 90846 9934 90846 9934 0 net85
rlabel metal4 90846 79954 90846 79954 0 net86
rlabel metal2 102166 37876 102166 37876 0 net87
rlabel metal1 90758 66504 90758 66504 0 net88
rlabel metal3 90827 79492 90827 79492 0 net89
rlabel metal4 23460 79410 23460 79410 0 net9
rlabel metal4 90559 79954 90559 79954 0 net90
rlabel metal4 90559 9866 90559 9866 0 net91
rlabel metal1 89378 66266 89378 66266 0 net92
rlabel metal2 90574 66130 90574 66130 0 net93
rlabel metal3 102164 22232 102164 22232 0 net94
rlabel metal1 89102 66028 89102 66028 0 net95
rlabel metal1 90114 66606 90114 66606 0 net96
rlabel metal3 102279 92232 102279 92232 0 net97
rlabel via1 103086 93857 103086 93857 0 net98
rlabel metal3 102026 23360 102026 23360 0 net99
rlabel metal2 108514 67541 108514 67541 0 rst
rlabel metal3 751 76228 751 76228 0 sine_out[0]
rlabel metal2 108514 72913 108514 72913 0 sine_out[10]
rlabel via2 108514 78965 108514 78965 0 sine_out[11]
rlabel metal2 108514 78353 108514 78353 0 sine_out[12]
rlabel metal2 108514 77741 108514 77741 0 sine_out[13]
rlabel via2 108514 76245 108514 76245 0 sine_out[14]
rlabel via2 108514 76891 108514 76891 0 sine_out[15]
rlabel metal3 751 72828 751 72828 0 sine_out[1]
rlabel metal3 751 73508 751 73508 0 sine_out[2]
rlabel metal3 751 74188 751 74188 0 sine_out[3]
rlabel metal3 751 74868 751 74868 0 sine_out[4]
rlabel metal3 1050 75548 1050 75548 0 sine_out[5]
rlabel via2 108514 73525 108514 73525 0 sine_out[6]
rlabel metal2 108514 74137 108514 74137 0 sine_out[7]
rlabel metal2 108514 75021 108514 75021 0 sine_out[8]
rlabel metal2 108514 75803 108514 75803 0 sine_out[9]
rlabel metal4 36107 63983 36107 63983 0 sine_out_temp0\[0\]
rlabel metal4 61134 64260 61134 64260 0 sine_out_temp0\[10\]
rlabel via3 63595 66164 63595 66164 0 sine_out_temp0\[11\]
rlabel metal4 66059 63983 66059 63983 0 sine_out_temp0\[12\]
rlabel metal1 76084 77146 76084 77146 0 sine_out_temp0\[13\]
rlabel metal1 78890 77554 78890 77554 0 sine_out_temp0\[14\]
rlabel metal2 80086 77996 80086 77996 0 sine_out_temp0\[15\]
rlabel metal4 38575 64260 38575 64260 0 sine_out_temp0\[1\]
rlabel metal4 41099 63983 41099 63983 0 sine_out_temp0\[2\]
rlabel metal4 43654 64260 43654 64260 0 sine_out_temp0\[3\]
rlabel via3 46115 66164 46115 66164 0 sine_out_temp0\[4\]
rlabel metal1 43102 77418 43102 77418 0 sine_out_temp0\[5\]
rlabel metal1 60996 77418 60996 77418 0 sine_out_temp0\[6\]
rlabel metal2 62514 77792 62514 77792 0 sine_out_temp0\[7\]
rlabel metal4 56051 64260 56051 64260 0 sine_out_temp0\[8\]
rlabel metal4 58571 63983 58571 63983 0 sine_out_temp0\[9\]
rlabel metal2 36110 135014 36110 135014 0 sine_out_temp1\[0\]
rlabel metal4 61088 134003 61088 134003 0 sine_out_temp1\[10\]
rlabel metal2 64446 135643 64446 135643 0 sine_out_temp1\[11\]
rlabel metal4 66059 134003 66059 134003 0 sine_out_temp1\[12\]
rlabel metal4 68540 134479 68540 134479 0 sine_out_temp1\[13\]
rlabel metal4 71051 134003 71051 134003 0 sine_out_temp1\[14\]
rlabel metal4 73547 133935 73547 133935 0 sine_out_temp1\[15\]
rlabel metal4 38603 133935 38603 133935 0 sine_out_temp1\[1\]
rlabel metal4 41099 133935 41099 133935 0 sine_out_temp1\[2\]
rlabel metal4 43595 133799 43595 133799 0 sine_out_temp1\[3\]
rlabel metal4 46091 133799 46091 133799 0 sine_out_temp1\[4\]
rlabel metal4 48576 133799 48576 133799 0 sine_out_temp1\[5\]
rlabel metal4 51083 133935 51083 133935 0 sine_out_temp1\[6\]
rlabel metal2 55798 135099 55798 135099 0 sine_out_temp1\[7\]
rlabel metal4 56075 133935 56075 133935 0 sine_out_temp1\[8\]
rlabel metal4 58571 134003 58571 134003 0 sine_out_temp1\[9\]
rlabel metal1 83858 77520 83858 77520 0 tcout\[0\]
rlabel metal2 86526 77452 86526 77452 0 tcout\[1\]
rlabel metal1 91034 71570 91034 71570 0 tcout\[2\]
rlabel metal1 92184 71978 92184 71978 0 tcout\[3\]
rlabel metal1 89056 67218 89056 67218 0 tcout\[4\]
rlabel metal2 91218 65892 91218 65892 0 tcout\[5\]
rlabel metal2 90390 65926 90390 65926 0 tcout\[6\]
rlabel metal2 89378 66640 89378 66640 0 tcout\[7\]
rlabel metal2 75118 71774 75118 71774 0 tcout\[8\]
<< properties >>
string FIXED_BBOX 0 0 110000 150000
<< end >>
