logic [0:255] [15:0] sine_table1 = {
16'h0000,
16'hfe6e,
16'hfcdc,
16'hfb4a,
16'hf9b8,
16'hf827,
16'hf696,
16'hf505,
16'hf374,
16'hf1e4,
16'hf055,
16'heec6,
16'hed38,
16'hebab,
16'hea1e,
16'he892,
16'he707,
16'he57e,
16'he3f5,
16'he26d,
16'he0e6,
16'hdf61,
16'hdddd,
16'hdc5a,
16'hdad8,
16'hd958,
16'hd7da,
16'hd65d,
16'hd4e1,
16'hd367,
16'hd1ef,
16'hd079,
16'hcf05,
16'hcd92,
16'hcc21,
16'hcab3,
16'hc946,
16'hc7dc,
16'hc674,
16'hc50e,
16'hc3aa,
16'hc248,
16'hc0e9,
16'hbf8d,
16'hbe32,
16'hbcdb,
16'hbb86,
16'hba33,
16'hb8e4,
16'hb797,
16'hb64c,
16'hb505,
16'hb3c1,
16'hb27f,
16'hb141,
16'hb005,
16'haecd,
16'had98,
16'hac65,
16'hab37,
16'haa0b,
16'ha8e3,
16'ha7be,
16'ha69c,
16'ha57e,
16'ha464,
16'ha34d,
16'ha239,
16'ha129,
16'ha01d,
16'h9f15,
16'h9e10,
16'h9d0f,
16'h9c12,
16'h9b18,
16'h9a23,
16'h9931,
16'h9844,
16'h975a,
16'h9675,
16'h9593,
16'h94b6,
16'h93dd,
16'h9308,
16'h9237,
16'h916a,
16'h90a2,
16'h8fde,
16'h8f1e,
16'h8e63,
16'h8dac,
16'h8cf9,
16'h8c4b,
16'h8ba1,
16'h8afc,
16'h8a5b,
16'h89bf,
16'h8928,
16'h8895,
16'h8806,
16'h877c,
16'h86f7,
16'h8677,
16'h85fb,
16'h8584,
16'h8512,
16'h84a4,
16'h843b,
16'h83d7,
16'h8378,
16'h831d,
16'h82c7,
16'h8277,
16'h822b,
16'h81e3,
16'h81a1,
16'h8164,
16'h812b,
16'h80f7,
16'h80c9,
16'h809f,
16'h807a,
16'h805a,
16'h803f,
16'h8028,
16'h8017,
16'h800b,
16'h8003,
16'h8001,
16'h8003,
16'h800b,
16'h8017,
16'h8028,
16'h803f,
16'h805a,
16'h807a,
16'h809f,
16'h80c9,
16'h80f7,
16'h812b,
16'h8164,
16'h81a1,
16'h81e3,
16'h822b,
16'h8277,
16'h82c7,
16'h831d,
16'h8378,
16'h83d7,
16'h843b,
16'h84a4,
16'h8512,
16'h8584,
16'h85fb,
16'h8677,
16'h86f7,
16'h877c,
16'h8806,
16'h8895,
16'h8928,
16'h89bf,
16'h8a5b,
16'h8afc,
16'h8ba1,
16'h8c4b,
16'h8cf9,
16'h8dac,
16'h8e63,
16'h8f1e,
16'h8fde,
16'h90a2,
16'h916a,
16'h9237,
16'h9308,
16'h93dd,
16'h94b6,
16'h9593,
16'h9675,
16'h975a,
16'h9844,
16'h9931,
16'h9a23,
16'h9b18,
16'h9c12,
16'h9d0f,
16'h9e10,
16'h9f15,
16'ha01d,
16'ha129,
16'ha239,
16'ha34d,
16'ha464,
16'ha57e,
16'ha69c,
16'ha7be,
16'ha8e3,
16'haa0b,
16'hab37,
16'hac65,
16'had98,
16'haecd,
16'hb005,
16'hb141,
16'hb27f,
16'hb3c1,
16'hb505,
16'hb64c,
16'hb797,
16'hb8e4,
16'hba33,
16'hbb86,
16'hbcdb,
16'hbe32,
16'hbf8d,
16'hc0e9,
16'hc248,
16'hc3aa,
16'hc50e,
16'hc674,
16'hc7dc,
16'hc946,
16'hcab3,
16'hcc21,
16'hcd92,
16'hcf05,
16'hd079,
16'hd1ef,
16'hd367,
16'hd4e1,
16'hd65d,
16'hd7da,
16'hd958,
16'hdad8,
16'hdc5a,
16'hdddd,
16'hdf61,
16'he0e6,
16'he26d,
16'he3f5,
16'he57e,
16'he707,
16'he892,
16'hea1e,
16'hebab,
16'hed38,
16'heec6,
16'hf055,
16'hf1e4,
16'hf374,
16'hf505,
16'hf696,
16'hf827,
16'hf9b8,
16'hfb4a,
16'hfcdc,
16'hfe6e
};
