module counter (clk,
    csb00,
    csb01,
    rst,
    addr00,
    addr01,
    din00,
    din01,
    sine_out);
 input clk;
 input csb00;
 input csb01;
 input rst;
 input [7:0] addr00;
 input [7:0] addr01;
 input [15:0] din00;
 input [15:0] din01;
 output [15:0] sine_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire net135;
 wire clknet_0_clk;
 wire \sine_out_temp0[0] ;
 wire \sine_out_temp0[10] ;
 wire \sine_out_temp0[11] ;
 wire \sine_out_temp0[12] ;
 wire \sine_out_temp0[13] ;
 wire \sine_out_temp0[14] ;
 wire \sine_out_temp0[15] ;
 wire \sine_out_temp0[1] ;
 wire \sine_out_temp0[2] ;
 wire \sine_out_temp0[3] ;
 wire \sine_out_temp0[4] ;
 wire \sine_out_temp0[5] ;
 wire \sine_out_temp0[6] ;
 wire \sine_out_temp0[7] ;
 wire \sine_out_temp0[8] ;
 wire \sine_out_temp0[9] ;
 wire \sine_out_temp1[0] ;
 wire \sine_out_temp1[10] ;
 wire \sine_out_temp1[11] ;
 wire \sine_out_temp1[12] ;
 wire \sine_out_temp1[13] ;
 wire \sine_out_temp1[14] ;
 wire \sine_out_temp1[15] ;
 wire \sine_out_temp1[1] ;
 wire \sine_out_temp1[2] ;
 wire \sine_out_temp1[3] ;
 wire \sine_out_temp1[4] ;
 wire \sine_out_temp1[5] ;
 wire \sine_out_temp1[6] ;
 wire \sine_out_temp1[7] ;
 wire \sine_out_temp1[8] ;
 wire \sine_out_temp1[9] ;
 wire \tcout[0] ;
 wire \tcout[1] ;
 wire \tcout[2] ;
 wire \tcout[3] ;
 wire \tcout[4] ;
 wire \tcout[5] ;
 wire \tcout[6] ;
 wire \tcout[7] ;
 wire \tcout[8] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire net136;
 wire net137;

 sky130_fd_sc_hd__inv_2 _061_ (.A(net130),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _062_ (.A(net131),
    .Y(_025_));
 sky130_fd_sc_hd__mux2_1 _063_ (.A0(net99),
    .A1(net83),
    .S(net100),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _064_ (.A0(net92),
    .A1(net76),
    .S(net100),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _065_ (.A0(net91),
    .A1(net75),
    .S(net100),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _066_ (.A0(net90),
    .A1(net74),
    .S(net100),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _067_ (.A0(net89),
    .A1(net73),
    .S(net100),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _068_ (.A0(net88),
    .A1(net72),
    .S(net100),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _069_ (.A0(net87),
    .A1(net71),
    .S(net100),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _070_ (.A0(net86),
    .A1(net70),
    .S(net100),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _071_ (.A0(net85),
    .A1(net69),
    .S(net100),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _072_ (.A0(net84),
    .A1(net68),
    .S(net100),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _073_ (.A0(net98),
    .A1(net82),
    .S(net101),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _074_ (.A0(net97),
    .A1(net81),
    .S(net101),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _075_ (.A0(net96),
    .A1(net80),
    .S(net101),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _076_ (.A0(net95),
    .A1(net79),
    .S(net101),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _077_ (.A0(net94),
    .A1(net78),
    .S(net101),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _078_ (.A0(net93),
    .A1(net77),
    .S(net101),
    .X(_006_));
 sky130_fd_sc_hd__xor2_1 _079_ (.A(net129),
    .B(net125),
    .X(_017_));
 sky130_fd_sc_hd__and3_1 _080_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .C(\tcout[2] ),
    .X(_050_));
 sky130_fd_sc_hd__a21oi_1 _081_ (.A1(\tcout[0] ),
    .A2(\tcout[1] ),
    .B1(\tcout[2] ),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_1 _082_ (.A(_050_),
    .B(_051_),
    .Y(_018_));
 sky130_fd_sc_hd__and4_2 _083_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .C(net120),
    .D(\tcout[3] ),
    .X(_052_));
 sky130_fd_sc_hd__nor2_1 _084_ (.A(\tcout[3] ),
    .B(_050_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_1 _085_ (.A(_052_),
    .B(_053_),
    .Y(_019_));
 sky130_fd_sc_hd__xor2_1 _086_ (.A(net137),
    .B(_052_),
    .X(_020_));
 sky130_fd_sc_hd__and3_1 _087_ (.A(net115),
    .B(\tcout[5] ),
    .C(_052_),
    .X(_054_));
 sky130_fd_sc_hd__a21oi_1 _088_ (.A1(net115),
    .A2(_052_),
    .B1(\tcout[5] ),
    .Y(_055_));
 sky130_fd_sc_hd__nor2_1 _089_ (.A(_054_),
    .B(_055_),
    .Y(_021_));
 sky130_fd_sc_hd__xor2_1 _090_ (.A(net136),
    .B(_054_),
    .X(_022_));
 sky130_fd_sc_hd__and2_1 _091_ (.A(net106),
    .B(net103),
    .X(_056_));
 sky130_fd_sc_hd__and4_1 _092_ (.A(net113),
    .B(\tcout[5] ),
    .C(_052_),
    .D(_056_),
    .X(_057_));
 sky130_fd_sc_hd__a41o_1 _093_ (.A1(net115),
    .A2(net110),
    .A3(net107),
    .A4(_052_),
    .B1(\tcout[7] ),
    .X(_058_));
 sky130_fd_sc_hd__and2b_1 _094_ (.A_N(_057_),
    .B(_058_),
    .X(_023_));
 sky130_fd_sc_hd__xor2_1 _095_ (.A(net101),
    .B(_057_),
    .X(_024_));
 sky130_fd_sc_hd__inv_2 _096_ (.A(net131),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _097_ (.A(net131),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _098_ (.A(net131),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _099_ (.A(net131),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _100_ (.A(net131),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _101_ (.A(net131),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _102_ (.A(net133),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _103_ (.A(net133),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _104_ (.A(net133),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _105_ (.A(net133),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _106_ (.A(net133),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _107_ (.A(net132),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _108_ (.A(net131),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _109_ (.A(net131),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _110_ (.A(net131),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _111_ (.A(net133),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _112_ (.A(net132),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _113_ (.A(net132),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _114_ (.A(net132),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _115_ (.A(net132),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _116_ (.A(net132),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _117_ (.A(net132),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _118_ (.A(net132),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _119_ (.A(net132),
    .Y(_049_));
 sky130_fd_sc_hd__dfrtp_1 _120_ (.CLK(clknet_2_0_0_clk),
    .D(_014_),
    .RESET_B(_025_),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_1 _121_ (.CLK(clknet_2_0_0_clk),
    .D(_015_),
    .RESET_B(_026_),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _122_ (.CLK(clknet_2_3_0_clk),
    .D(_001_),
    .RESET_B(_027_),
    .Q(net53));
 sky130_fd_sc_hd__dfrtp_1 _123_ (.CLK(clknet_2_3_0_clk),
    .D(_002_),
    .RESET_B(_028_),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_1 _124_ (.CLK(clknet_2_3_0_clk),
    .D(_003_),
    .RESET_B(_029_),
    .Q(net55));
 sky130_fd_sc_hd__dfrtp_1 _125_ (.CLK(clknet_2_3_0_clk),
    .D(_004_),
    .RESET_B(_030_),
    .Q(net56));
 sky130_fd_sc_hd__dfrtp_1 _126_ (.CLK(clknet_2_2_0_clk),
    .D(_005_),
    .RESET_B(_031_),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _127_ (.CLK(clknet_2_2_0_clk),
    .D(_006_),
    .RESET_B(_032_),
    .Q(net58));
 sky130_fd_sc_hd__dfrtp_1 _128_ (.CLK(clknet_2_3_0_clk),
    .D(_016_),
    .RESET_B(_033_),
    .Q(\tcout[0] ));
 sky130_fd_sc_hd__dfrtp_1 _129_ (.CLK(clknet_2_3_0_clk),
    .D(_017_),
    .RESET_B(_034_),
    .Q(\tcout[1] ));
 sky130_fd_sc_hd__dfrtp_1 _130_ (.CLK(clknet_2_3_0_clk),
    .D(_018_),
    .RESET_B(_035_),
    .Q(\tcout[2] ));
 sky130_fd_sc_hd__dfrtp_1 _131_ (.CLK(clknet_2_3_0_clk),
    .D(_019_),
    .RESET_B(_036_),
    .Q(\tcout[3] ));
 sky130_fd_sc_hd__dfrtp_1 _132_ (.CLK(clknet_2_2_0_clk),
    .D(_020_),
    .RESET_B(_037_),
    .Q(\tcout[4] ));
 sky130_fd_sc_hd__dfrtp_1 _133_ (.CLK(clknet_2_2_0_clk),
    .D(_021_),
    .RESET_B(_038_),
    .Q(\tcout[5] ));
 sky130_fd_sc_hd__dfrtp_1 _134_ (.CLK(clknet_2_2_0_clk),
    .D(_022_),
    .RESET_B(_039_),
    .Q(\tcout[6] ));
 sky130_fd_sc_hd__dfrtp_1 _135_ (.CLK(clknet_2_2_0_clk),
    .D(_023_),
    .RESET_B(_040_),
    .Q(\tcout[7] ));
 sky130_fd_sc_hd__dfrtp_1 _136_ (.CLK(clknet_2_3_0_clk),
    .D(_024_),
    .RESET_B(_041_),
    .Q(\tcout[8] ));
 sky130_fd_sc_hd__dfrtp_1 _137_ (.CLK(clknet_2_1_0_clk),
    .D(_000_),
    .RESET_B(_042_),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_1 _138_ (.CLK(clknet_2_1_0_clk),
    .D(_007_),
    .RESET_B(_043_),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_1 _139_ (.CLK(clknet_2_0_0_clk),
    .D(_008_),
    .RESET_B(_044_),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _140_ (.CLK(clknet_2_1_0_clk),
    .D(_009_),
    .RESET_B(_045_),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_1 _141_ (.CLK(clknet_2_1_0_clk),
    .D(_010_),
    .RESET_B(_046_),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_1 _142_ (.CLK(clknet_2_1_0_clk),
    .D(_011_),
    .RESET_B(_047_),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_1 _143_ (.CLK(clknet_2_1_0_clk),
    .D(_012_),
    .RESET_B(_048_),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _144_ (.CLK(clknet_2_0_0_clk),
    .D(_013_),
    .RESET_B(_049_),
    .Q(net65));
 sky130_fd_sc_hd__conb_1 mem_i1_135 (.LO(net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 ram_256x16 mem_i0 (.csb0(net17),
    .csb1(net134),
    .clk0(clknet_2_0_0_clk),
    .clk1(clknet_2_1_0_clk),
    .addr0({net8,
    net7,
    net6,
    net5,
    net4,
    net3,
    net2,
    net1}),
    .addr1({net104,
    net108,
    net111,
    net114,
    net117,
    net121,
    net123,
    net127}),
    .din0({net25,
    net24,
    net23,
    net22,
    net21,
    net20,
    net34,
    net33,
    net32,
    net31,
    net30,
    net29,
    net28,
    net27,
    net26,
    net19}),
    .dout1({\sine_out_temp0[15] ,
    \sine_out_temp0[14] ,
    \sine_out_temp0[13] ,
    \sine_out_temp0[12] ,
    \sine_out_temp0[11] ,
    \sine_out_temp0[10] ,
    \sine_out_temp0[9] ,
    \sine_out_temp0[8] ,
    \sine_out_temp0[7] ,
    \sine_out_temp0[6] ,
    \sine_out_temp0[5] ,
    \sine_out_temp0[4] ,
    \sine_out_temp0[3] ,
    \sine_out_temp0[2] ,
    \sine_out_temp0[1] ,
    \sine_out_temp0[0] }));
 ram_256x16 mem_i1 (.csb0(net18),
    .csb1(net135),
    .clk0(clknet_2_2_0_clk),
    .clk1(clknet_2_3_0_clk),
    .addr0({net16,
    net15,
    net14,
    net13,
    net12,
    net11,
    net10,
    net9}),
    .addr1({net102,
    net105,
    net109,
    net112,
    net116,
    net119,
    net122,
    net126}),
    .din0({net41,
    net40,
    net39,
    net38,
    net37,
    net36,
    net50,
    net49,
    net48,
    net47,
    net46,
    net45,
    net44,
    net43,
    net42,
    net35}),
    .dout1({\sine_out_temp1[15] ,
    \sine_out_temp1[14] ,
    \sine_out_temp1[13] ,
    \sine_out_temp1[12] ,
    \sine_out_temp1[11] ,
    \sine_out_temp1[10] ,
    \sine_out_temp1[9] ,
    \sine_out_temp1[8] ,
    \sine_out_temp1[7] ,
    \sine_out_temp1[6] ,
    \sine_out_temp1[5] ,
    \sine_out_temp1[4] ,
    \sine_out_temp1[3] ,
    \sine_out_temp1[2] ,
    \sine_out_temp1[1] ,
    \sine_out_temp1[0] }));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_246_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_247_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_248_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_249_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_250_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_251_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_252_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_253_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_254_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_255_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_256_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_257_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_258_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_259_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_260_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_261_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_262_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_263_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_264_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_265_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_266_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_267_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_268_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_269_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_270_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_271_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_272_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_273_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_274_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_275_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_276_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_277_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_278_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_279_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_280_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_281_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_282_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_283_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_284_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_285_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_3_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_3_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_3_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_3_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_3_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_3_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_3_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_3_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_3_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_3_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_3_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_3_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_3_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_3_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_3_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_3_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_3_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_3_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_3_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_3_Right_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_3_Right_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_3_Right_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_3_Right_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_3_Right_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_3_Right_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_3_Right_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_3_Right_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_3_Right_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_3_Right_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_3_Right_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_3_Right_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_3_Right_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_3_Right_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_3_Right_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_3_Right_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_3_Right_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_3_Right_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_3_Right_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_3_Right_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_3_Right_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_3_Right_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_3_Right_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_3_Right_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_3_Right_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_3_Right_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_3_Right_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_3_Right_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_3_Right_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_3_Right_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_3_Right_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_3_Right_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_3_Right_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_3_Right_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_3_Right_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_3_Right_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_3_Right_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_3_Right_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_3_Right_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_3_Right_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_3_Right_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_3_Right_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_3_Right_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_3_Right_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_3_Right_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_3_Right_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_3_Right_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_3_Right_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_3_Right_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_3_Right_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_3_Right_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_3_Right_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_3_Right_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_3_Right_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_3_Right_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_3_Right_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_3_Right_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_3_Right_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_3_Right_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_3_Right_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_3_Right_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_3_Right_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_3_Right_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_3_Right_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_3_Right_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_3_Right_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_3_Right_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_3_Right_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_3_Right_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_3_Right_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_3_Right_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_3_Right_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_3_Right_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_3_Right_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_3_Right_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_3_Right_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_3_Right_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_3_Right_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_3_Right_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_3_Right_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_3_Right_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_3_Right_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_3_Right_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_3_Right_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_3_Right_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_3_Right_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_3_Right_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_3_Right_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_444 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_445 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_446 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_447 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_448 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_449 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_450 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_451 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_452 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_453 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_454 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_455 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_456 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_457 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_458 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_459 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Left_460 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Left_461 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Left_462 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Left_463 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Left_464 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Left_465 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Left_466 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Left_467 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Left_468 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Left_469 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Left_470 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Left_471 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Left_472 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Left_473 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Left_474 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Left_475 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Left_476 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Left_477 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Left_478 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Left_479 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Left_480 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Left_481 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Left_482 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Left_483 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Left_484 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Left_485 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Left_486 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Left_487 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Left_488 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Left_489 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Left_490 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Left_491 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Left_492 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Left_493 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Left_494 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Left_495 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Left_496 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Left_497 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Left_498 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Left_499 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Left_500 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Left_501 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Left_502 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Left_503 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Left_504 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Left_505 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Left_506 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_Left_507 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_Left_508 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_Left_509 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_Left_510 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_Left_511 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_Left_512 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_Left_513 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_Left_514 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_Left_515 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_Left_516 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_Left_517 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_Left_518 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_Left_519 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_Left_520 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_Left_521 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_Left_522 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_Left_523 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_Left_524 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_Left_525 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_Left_526 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_Left_527 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_Left_528 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_Left_529 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_Left_530 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_246_Left_531 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_247_Left_532 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_248_Left_533 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_249_Left_534 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_250_Left_535 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_251_Left_536 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_252_Left_537 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_253_Left_538 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_254_Left_539 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_255_Left_540 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_256_Left_541 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_257_Left_542 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_258_Left_543 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_259_Left_544 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_260_Left_545 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_261_Left_546 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_262_Left_547 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_263_Left_548 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_264_Left_549 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_265_Left_550 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_266_Left_551 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_267_Left_552 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_268_Left_553 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_269_Left_554 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_270_Left_555 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_271_Left_556 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_272_Left_557 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_273_Left_558 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_274_Left_559 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_275_Left_560 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_276_Left_561 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_277_Left_562 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_278_Left_563 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_279_Left_564 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_280_Left_565 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_281_Left_566 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_282_Left_567 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_283_Left_568 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_284_Left_569 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_285_Left_570 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Left_571 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_572 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_573 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_574 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_575 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_576 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_577 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_578 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_579 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_580 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_581 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_582 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_583 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_584 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_585 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_586 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_587 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_588 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_589 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_590 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_591 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_592 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_593 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_594 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_595 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_596 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_597 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_598 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_599 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_600 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_601 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_602 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_603 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_604 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_605 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_606 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_607 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_608 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_609 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_610 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_611 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_612 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_613 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_614 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_615 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_616 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_617 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_618 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_619 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_620 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_621 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_622 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_623 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_624 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_625 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_626 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_627 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_628 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Left_629 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Left_630 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Left_631 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Left_632 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Left_633 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Left_634 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Left_635 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Left_636 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Left_637 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Left_638 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Left_639 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Left_640 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Left_641 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Left_642 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Left_643 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Left_644 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Left_645 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Left_646 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Left_647 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Left_648 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Left_649 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Left_650 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Left_651 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Left_652 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Left_653 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Left_654 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Left_655 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Left_656 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Left_657 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Left_658 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Left_659 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Left_660 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Left_661 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Left_662 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Left_663 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Left_664 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Left_665 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Left_666 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Left_667 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Left_668 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Left_669 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Left_670 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Left_671 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Left_672 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Left_673 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Left_674 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Left_675 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Left_676 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Left_677 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Left_678 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Right_679 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Right_680 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Right_681 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Right_682 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Right_683 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Right_684 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Right_685 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Right_686 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Right_687 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Right_688 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Right_689 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Right_690 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Right_691 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Right_692 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Right_693 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Right_694 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Right_695 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Right_696 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Right_697 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Right_698 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Right_699 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Right_700 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Right_701 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Right_702 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Right_703 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Right_704 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Right_705 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Right_706 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Right_707 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Right_708 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Right_709 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Right_710 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Right_711 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Right_712 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Right_713 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Right_714 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Right_715 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Right_716 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Right_717 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Right_718 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Right_719 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Right_720 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Right_721 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Right_722 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Right_723 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Right_724 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Right_725 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Right_726 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Right_727 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Right_728 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Right_729 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Right_730 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Right_731 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Right_732 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Right_733 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Right_734 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Right_735 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Right_736 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Right_737 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Right_738 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Right_739 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Right_740 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Right_741 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Right_742 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Right_743 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Right_744 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Right_745 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Right_746 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Right_747 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Right_748 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Right_749 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Right_750 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Right_751 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Right_752 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Right_753 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Right_754 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Right_755 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Right_756 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Right_757 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Right_758 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Right_759 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Right_760 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Right_761 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Right_762 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Right_763 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Right_764 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Right_765 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Right_766 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Right_767 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Right_768 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Right_769 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Right_770 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Right_771 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Right_772 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Right_773 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Right_774 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Right_775 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Right_776 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Right_777 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Right_778 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Right_779 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Right_780 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Right_781 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Right_782 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Right_783 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Right_784 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Right_785 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_3_Left_786 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_3_Left_787 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_3_Left_788 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_3_Left_789 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_3_Left_790 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_3_Left_791 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_3_Left_792 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_3_Left_793 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_3_Left_794 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_3_Left_795 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_3_Left_796 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_3_Left_797 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_3_Left_798 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_3_Left_799 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_3_Left_800 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_3_Left_801 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_3_Left_802 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_3_Left_803 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_3_Left_804 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_3_Left_805 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_3_Left_806 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_3_Left_807 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_3_Left_808 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_3_Left_809 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_3_Left_810 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_3_Left_811 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_3_Left_812 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_3_Left_813 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_3_Left_814 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_3_Left_815 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_3_Left_816 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_3_Left_817 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_3_Left_818 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_3_Left_819 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_3_Left_820 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_3_Left_821 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_3_Left_822 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_3_Left_823 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_3_Left_824 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_3_Left_825 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_3_Left_826 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_3_Left_827 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_3_Left_828 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_3_Left_829 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_3_Left_830 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_3_Left_831 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_3_Left_832 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_3_Left_833 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_3_Left_834 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_3_Left_835 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_3_Left_836 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_3_Left_837 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_3_Left_838 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_3_Left_839 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_3_Left_840 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_3_Left_841 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_3_Left_842 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_3_Left_843 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_3_Left_844 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_3_Left_845 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_3_Left_846 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_3_Left_847 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_3_Left_848 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_3_Left_849 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_3_Left_850 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_3_Left_851 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_3_Left_852 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_3_Left_853 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_3_Left_854 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_3_Left_855 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_3_Left_856 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_3_Left_857 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_3_Left_858 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_3_Left_859 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_3_Left_860 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_3_Left_861 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_3_Left_862 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_3_Left_863 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_3_Left_864 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_3_Left_865 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_3_Left_866 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_3_Left_867 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_3_Left_868 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_3_Left_869 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_3_Left_870 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_3_Left_871 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_3_Left_872 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_3_Left_873 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_3_Left_874 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_3_Left_875 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_3_Left_876 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_3_Left_877 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_3_Left_878 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_3_Left_879 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_3_Left_880 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_3_Left_881 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_3_Left_882 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_3_Left_883 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_3_Left_884 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_3_Left_885 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_3_Left_886 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_3_Left_887 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_3_Left_888 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_3_Left_889 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_3_Left_890 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_3_Left_891 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_3_Left_892 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_893 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_894 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_895 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_896 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_897 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_898 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_899 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_900 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_901 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_902 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_903 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_904 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_905 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_906 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_907 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_908 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_909 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_910 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_911 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_912 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_913 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_914 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_915 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_916 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_917 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_918 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_919 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_920 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_921 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_922 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_923 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_924 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_925 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_926 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_927 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_928 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_929 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_930 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_931 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_932 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_933 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_934 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_935 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_936 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_937 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_938 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_939 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_940 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_941 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_942 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_943 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_944 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_945 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_946 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_947 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_948 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_949 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Right_950 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Right_951 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Right_952 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Right_953 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Right_954 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Right_955 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Right_956 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Right_957 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Right_958 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Right_959 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Right_960 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Right_961 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Right_962 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Right_963 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Right_964 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Right_965 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Right_966 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Right_967 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Right_968 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Right_969 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Right_970 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Right_971 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Right_972 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Right_973 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Right_974 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Right_975 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Right_976 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Right_977 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Right_978 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Right_979 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Right_980 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Right_981 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Right_982 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Right_983 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Right_984 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Right_985 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Right_986 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Right_987 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Right_988 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Right_989 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Right_990 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Right_991 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Right_992 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Right_993 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Right_994 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Right_995 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Right_996 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Right_997 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Right_998 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Right_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_267_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_268_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_269_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_270_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_271_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_272_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_273_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_274_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_275_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_276_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_277_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_278_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_279_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_280_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_281_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_282_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_283_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_284_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_285_9523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_9524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_9525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_9526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_9527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_9528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_9529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_3_9530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_3_9531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_3_9532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_2_9533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_2_9534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_2_9535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_2_9536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_3_9537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_3_9538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_9539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_9540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_9541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_9542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_9543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_3_9544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_3_9545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_3_9546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_2_9547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_2_9548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_2_9549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_2_9550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_3_9551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_3_9552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_9553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_9554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_9555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_9556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_9557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_3_9558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_3_9559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_3_9560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_2_9561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_2_9562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_2_9563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_2_9564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_3_9565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_3_9566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_9567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_9568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_9569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_9570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_9571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_3_9572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_3_9573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_3_9574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_2_9575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_2_9576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_2_9577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_2_9578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_3_9579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_3_9580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_9581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_9582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_9583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_9584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_9585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_3_9586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_3_9587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_3_9588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_2_9589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_2_9590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_2_9591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_2_9592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_3_9593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_3_9594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_9595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_9596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_9597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_9598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_9599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_3_9600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_3_9601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_3_9602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_2_9603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_2_9604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_2_9605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_2_9606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_3_9607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_3_9608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_9609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_9610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_9611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_9612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_9613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_3_9614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_3_9615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_3_9616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_2_9617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_2_9618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_2_9619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_2_9620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_3_9621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_3_9622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_9623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_9624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_9625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_9626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_9627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_3_9628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_3_9629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_3_9630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_2_9631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_2_9632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_2_9633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_2_9634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_3_9635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_3_9636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_9637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_9638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_9639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_9640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_9641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_3_9642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_3_9643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_3_9644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_2_9645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_2_9646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_2_9647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_2_9648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_3_9649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_3_9650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_9651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_9652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_9653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_9654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_9655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_3_9656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_3_9657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_3_9658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_2_9659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_2_9660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_2_9661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_2_9662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_3_9663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_3_9664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_9665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_9666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_9667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_9668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_9669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_3_9670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_3_9671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_3_9672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2_9673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2_9674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2_9675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2_9676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_3_9677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_3_9678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_9679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_9680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_9681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_9682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_9683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_3_9684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_3_9685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_3_9686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2_9687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2_9688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2_9689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2_9690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_3_9691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_3_9692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_9693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_9694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_9695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_9696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_9697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_3_9698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_3_9699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_3_9700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_2_9701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_2_9702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_2_9703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_2_9704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_3_9705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_3_9706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_9707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_9708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_9709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_9710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_9711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_3_9712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_3_9713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_3_9714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_2_9715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_2_9716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_2_9717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_2_9718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_3_9719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_3_9720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_9721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_9722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_9723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_9724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_9725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_3_9726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_3_9727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_3_9728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_2_9729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_2_9730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_2_9731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_2_9732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_3_9733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_3_9734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_9735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_9736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_9737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_9738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_9739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_3_9740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_3_9741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_3_9742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_2_9743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_2_9744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_2_9745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_2_9746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_3_9747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_3_9748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_9749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_9750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_9751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_9752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_9753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_3_9754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_3_9755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_3_9756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_2_9757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_2_9758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_2_9759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_2_9760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_3_9761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_3_9762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_9763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_9764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_9765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_9766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_9767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_3_9768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_3_9769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_3_9770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_2_9771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_2_9772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_2_9773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_2_9774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_3_9775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_3_9776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_9777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_9778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_9779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_9780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_9781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_3_9782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_3_9783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_3_9784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_2_9785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_2_9786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_2_9787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_2_9788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_3_9789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_3_9790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_9791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_9792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_9793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_9794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_9795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_3_9796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_3_9797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_3_9798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_2_9799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_2_9800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_2_9801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_2_9802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_3_9803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_3_9804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_9805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_9806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_9807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_9808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_9809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_3_9810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_3_9811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_3_9812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_2_9813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_2_9814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_2_9815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_2_9816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_3_9817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_3_9818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_9819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_9820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_9821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_9822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_9823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_3_9824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_3_9825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_3_9826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_2_9827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_2_9828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_2_9829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_2_9830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_3_9831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_3_9832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_9833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_9834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_9835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_9836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_9837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_3_9838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_3_9839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_3_9840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_2_9841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_2_9842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_2_9843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_2_9844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_3_9845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_3_9846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_9847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_9848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_9849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_9850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_9851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_3_9852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_3_9853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_3_9854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2_9855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2_9856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2_9857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2_9858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_3_9859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_3_9860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_9861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_9862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_9863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_9864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_9865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_3_9866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_3_9867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_3_9868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2_9869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2_9870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2_9871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2_9872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_3_9873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_3_9874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_9875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_9876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_9877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_9878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_9879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_3_9880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_3_9881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_3_9882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2_9883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2_9884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2_9885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2_9886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_3_9887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_3_9888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_9889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_9890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_9891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_9892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_9893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_3_9894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_3_9895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_3_9896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2_9897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2_9898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2_9899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2_9900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_3_9901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_3_9902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_9903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_9904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_9905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_9906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_9907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_3_9908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_3_9909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_3_9910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2_9911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2_9912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2_9913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2_9914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_3_9915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_3_9916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_9917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_9918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_9919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_9920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_9921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_3_9922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_3_9923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_3_9924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2_9925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2_9926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2_9927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2_9928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_3_9929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_3_9930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_9931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_9932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_9933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_9934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_9935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_3_9936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_3_9937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_3_9938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2_9939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2_9940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2_9941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2_9942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_3_9943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_3_9944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_9945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_9946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_9947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_9948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_9949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_3_9950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_3_9951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_3_9952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2_9953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2_9954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2_9955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2_9956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_3_9957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_3_9958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_9959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_9960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_9961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_9962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_9963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_3_9964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_3_9965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_3_9966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2_9967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2_9968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2_9969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2_9970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_3_9971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_3_9972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_9973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_9974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_9975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_9976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_9977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_3_9978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_3_9979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_3_9980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2_9981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2_9982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2_9983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2_9984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_3_9985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_3_9986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_9987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_9988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_9989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_9990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_9991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_3_9992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_3_9993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_3_9994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2_9995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2_9996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2_9997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2_9998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_3_9999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_3_10000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_10001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_10002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_10003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_10004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_10005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_3_10006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_3_10007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_3_10008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2_10009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2_10010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2_10011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2_10012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_3_10013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_3_10014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_10015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_10016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_10017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_10018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_10019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_3_10020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_3_10021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_3_10022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2_10023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2_10024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2_10025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2_10026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_3_10027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_3_10028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_10029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_10030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_10031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_10032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_10033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_3_10034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_3_10035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_3_10036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2_10037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2_10038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2_10039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2_10040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_3_10041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_3_10042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_10043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_10044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_10045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_10046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_10047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_3_10048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_3_10049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_3_10050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2_10051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2_10052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2_10053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2_10054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_3_10055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_3_10056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_10057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_10058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_10059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_10060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_10061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_3_10062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_3_10063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_3_10064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2_10065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2_10066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2_10067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2_10068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_3_10069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_3_10070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_10071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_10072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_10073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_10074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_10075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_3_10076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_3_10077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_3_10078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2_10079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2_10080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2_10081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2_10082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_3_10083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_3_10084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_10085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_10086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_10087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_10088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_10089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_3_10090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_3_10091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_3_10092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2_10093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2_10094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2_10095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2_10096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_3_10097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_3_10098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_10099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_10100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_10101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_10102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_10103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_3_10104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_3_10105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_3_10106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2_10107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2_10108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2_10109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2_10110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_3_10111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_3_10112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_10113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_10114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_10115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_10116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_10117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_3_10118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_3_10119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_3_10120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2_10121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2_10122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2_10123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2_10124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3_10125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3_10126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_10127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_10128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_10129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_10130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_10131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3_10132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3_10133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3_10134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2_10135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2_10136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2_10137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2_10138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3_10139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3_10140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_10141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_10142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_10143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_10144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_10145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3_10146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3_10147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3_10148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2_10149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2_10150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2_10151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2_10152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3_10153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3_10154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_10155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_10156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_10157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_10158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_10159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3_10160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3_10161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3_10162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2_10163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2_10164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2_10165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2_10166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3_10167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3_10168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_10169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_10170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_10171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_10172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_10173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3_10174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3_10175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3_10176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2_10177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2_10178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2_10179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2_10180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3_10181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3_10182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_10183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_10184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_10185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_10186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_10187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3_10188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3_10189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3_10190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2_10191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2_10192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2_10193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2_10194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3_10195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3_10196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_10197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_10198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_10199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_10200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_10201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3_10202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3_10203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3_10204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2_10205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2_10206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2_10207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2_10208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3_10209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3_10210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_10211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_10212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_10213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_10214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_10215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3_10216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3_10217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3_10218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2_10219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2_10220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2_10221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2_10222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3_10223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3_10224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_10225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_10226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_10227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_10228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_10229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3_10230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3_10231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3_10232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2_10233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2_10234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2_10235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2_10236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3_10237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3_10238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_10239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_10240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_10241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_10242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_10243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3_10244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3_10245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3_10246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2_10247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2_10248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2_10249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2_10250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3_10251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3_10252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_10253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_10254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_10255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_10256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_10257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3_10258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3_10259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3_10260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2_10261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2_10262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2_10263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2_10264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3_10265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3_10266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_10267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_10268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_10269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_10270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_10271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3_10272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3_10273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3_10274 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(addr00[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(addr00[1]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(addr00[2]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(addr00[3]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(addr00[4]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(addr00[5]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(addr00[6]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(addr00[7]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(addr01[0]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(addr01[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(addr01[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(addr01[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(addr01[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(addr01[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(addr01[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(addr01[7]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(csb00),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(csb01),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(din00[0]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(din00[10]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(din00[11]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(din00[12]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(din00[13]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(din00[14]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(din00[15]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(din00[1]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(din00[2]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(din00[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(din00[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(din00[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(din00[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(din00[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(din00[8]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(din00[9]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(din01[0]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(din01[10]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(din01[11]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(din01[12]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(din01[13]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(din01[14]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(din01[15]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(din01[1]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(din01[2]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(din01[3]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(din01[4]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(din01[5]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(din01[6]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(din01[7]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(din01[8]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(din01[9]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(rst),
    .X(net51));
 sky130_fd_sc_hd__buf_1 output52 (.A(net52),
    .X(sine_out[0]));
 sky130_fd_sc_hd__buf_1 output53 (.A(net53),
    .X(sine_out[10]));
 sky130_fd_sc_hd__buf_1 output54 (.A(net54),
    .X(sine_out[11]));
 sky130_fd_sc_hd__buf_1 output55 (.A(net55),
    .X(sine_out[12]));
 sky130_fd_sc_hd__buf_1 output56 (.A(net56),
    .X(sine_out[13]));
 sky130_fd_sc_hd__buf_1 output57 (.A(net57),
    .X(sine_out[14]));
 sky130_fd_sc_hd__buf_1 output58 (.A(net58),
    .X(sine_out[15]));
 sky130_fd_sc_hd__buf_1 output59 (.A(net59),
    .X(sine_out[1]));
 sky130_fd_sc_hd__buf_1 output60 (.A(net60),
    .X(sine_out[2]));
 sky130_fd_sc_hd__buf_1 output61 (.A(net61),
    .X(sine_out[3]));
 sky130_fd_sc_hd__buf_1 output62 (.A(net62),
    .X(sine_out[4]));
 sky130_fd_sc_hd__buf_1 output63 (.A(net63),
    .X(sine_out[5]));
 sky130_fd_sc_hd__buf_1 output64 (.A(net64),
    .X(sine_out[6]));
 sky130_fd_sc_hd__buf_1 output65 (.A(net65),
    .X(sine_out[7]));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(sine_out[8]));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(sine_out[9]));
 sky130_fd_sc_hd__clkbuf_2 wire68 (.A(\sine_out_temp1[9] ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 wire69 (.A(\sine_out_temp1[8] ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 wire70 (.A(\sine_out_temp1[7] ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 wire71 (.A(\sine_out_temp1[6] ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 wire72 (.A(\sine_out_temp1[5] ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 wire73 (.A(\sine_out_temp1[4] ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 wire74 (.A(\sine_out_temp1[3] ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 wire75 (.A(\sine_out_temp1[2] ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 wire76 (.A(\sine_out_temp1[1] ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 wire77 (.A(\sine_out_temp1[15] ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 wire78 (.A(\sine_out_temp1[14] ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 wire79 (.A(\sine_out_temp1[13] ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 wire80 (.A(\sine_out_temp1[12] ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 wire81 (.A(\sine_out_temp1[11] ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 wire82 (.A(\sine_out_temp1[10] ),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 wire83 (.A(\sine_out_temp1[0] ),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 wire84 (.A(\sine_out_temp0[9] ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 wire85 (.A(\sine_out_temp0[8] ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 wire86 (.A(\sine_out_temp0[7] ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 wire87 (.A(\sine_out_temp0[6] ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 wire88 (.A(\sine_out_temp0[5] ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 wire89 (.A(\sine_out_temp0[4] ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 wire90 (.A(\sine_out_temp0[3] ),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 wire91 (.A(\sine_out_temp0[2] ),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 wire92 (.A(\sine_out_temp0[1] ),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 wire93 (.A(\sine_out_temp0[15] ),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 wire94 (.A(\sine_out_temp0[14] ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 wire95 (.A(\sine_out_temp0[13] ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 wire96 (.A(\sine_out_temp0[12] ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 wire97 (.A(\sine_out_temp0[11] ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 wire98 (.A(\sine_out_temp0[10] ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 wire99 (.A(\sine_out_temp0[0] ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 fanout100 (.A(\tcout[8] ),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 fanout101 (.A(\tcout[8] ),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 wire102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_2 load_slew103 (.A(\tcout[7] ),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 load_slew104 (.A(\tcout[7] ),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 wire105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__buf_2 load_slew106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_1 load_slew107 (.A(\tcout[6] ),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 load_slew108 (.A(\tcout[6] ),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 wire109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 load_slew110 (.A(\tcout[5] ),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 load_slew111 (.A(\tcout[5] ),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 wire112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_4 load_slew113 (.A(net115),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 load_slew114 (.A(\tcout[4] ),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 load_slew115 (.A(\tcout[4] ),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 wire116 (.A(net118),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 load_slew117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_4 load_slew118 (.A(\tcout[3] ),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 wire119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__buf_4 load_slew120 (.A(\tcout[2] ),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 load_slew121 (.A(\tcout[2] ),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 wire122 (.A(net124),
    .X(net122));
 sky130_fd_sc_hd__buf_4 load_slew123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_4 load_slew124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_1 load_slew125 (.A(\tcout[1] ),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 wire126 (.A(net128),
    .X(net126));
 sky130_fd_sc_hd__buf_4 load_slew127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_4 load_slew128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__buf_1 load_slew129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__buf_1 load_slew130 (.A(\tcout[0] ),
    .X(net130));
 sky130_fd_sc_hd__buf_4 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_4 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net51),
    .X(net133));
 sky130_fd_sc_hd__conb_1 mem_i0_134 (.LO(net134));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload1 (.A(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload2 (.A(clknet_2_2_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\tcout[6] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\tcout[4] ),
    .X(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__D (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__063__X (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__D (.DIODE(_001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__X (.DIODE(_001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__D (.DIODE(_002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__074__X (.DIODE(_002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__D (.DIODE(_003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__X (.DIODE(_003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__D (.DIODE(_004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__076__X (.DIODE(_004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__D (.DIODE(_005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__077__X (.DIODE(_005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__D (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__078__X (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__D (.DIODE(_007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__064__X (.DIODE(_007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__D (.DIODE(_008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__065__X (.DIODE(_008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__D (.DIODE(_009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__066__X (.DIODE(_009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__D (.DIODE(_010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__X (.DIODE(_010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__D (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__X (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__D (.DIODE(_012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__X (.DIODE(_012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__D (.DIODE(_013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__X (.DIODE(_013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__D (.DIODE(_014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__X (.DIODE(_014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__D (.DIODE(_015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__072__X (.DIODE(_015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__092__D (.DIODE(_056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__091__X (.DIODE(_056_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(addr00[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(addr00[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(addr00[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(addr00[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(addr00[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(addr00[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(addr00[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(addr00[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(addr01[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(addr01[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(addr01[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(addr01[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(addr01[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(addr01[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(addr01[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(addr01[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(csb00));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(csb01));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(din00[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(din00[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(din00[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(din00[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(din00[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(din00[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(din00[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(din00[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(din00[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(din00[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(din00[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(din00[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(din00[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(din00[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(din00[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(din00[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(din01[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(din01[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(din01[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(din01[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(din01[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(din01[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(din01[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(din01[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(din01[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(din01[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(din01[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(din01[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(din01[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(din01[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(din01[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(din01[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire99_A (.DIODE(\sine_out_temp0[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[0]  (.DIODE(\sine_out_temp0[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire98_A (.DIODE(\sine_out_temp0[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[10]  (.DIODE(\sine_out_temp0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire97_A (.DIODE(\sine_out_temp0[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[11]  (.DIODE(\sine_out_temp0[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire96_A (.DIODE(\sine_out_temp0[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[12]  (.DIODE(\sine_out_temp0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire95_A (.DIODE(\sine_out_temp0[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[13]  (.DIODE(\sine_out_temp0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire94_A (.DIODE(\sine_out_temp0[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[14]  (.DIODE(\sine_out_temp0[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire93_A (.DIODE(\sine_out_temp0[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[15]  (.DIODE(\sine_out_temp0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire92_A (.DIODE(\sine_out_temp0[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[1]  (.DIODE(\sine_out_temp0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire91_A (.DIODE(\sine_out_temp0[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[2]  (.DIODE(\sine_out_temp0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire90_A (.DIODE(\sine_out_temp0[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[3]  (.DIODE(\sine_out_temp0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire89_A (.DIODE(\sine_out_temp0[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[4]  (.DIODE(\sine_out_temp0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire88_A (.DIODE(\sine_out_temp0[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[5]  (.DIODE(\sine_out_temp0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire87_A (.DIODE(\sine_out_temp0[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[6]  (.DIODE(\sine_out_temp0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire86_A (.DIODE(\sine_out_temp0[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[7]  (.DIODE(\sine_out_temp0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire85_A (.DIODE(\sine_out_temp0[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[8]  (.DIODE(\sine_out_temp0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire84_A (.DIODE(\sine_out_temp0[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[9]  (.DIODE(\sine_out_temp0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire83_A (.DIODE(\sine_out_temp1[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[0]  (.DIODE(\sine_out_temp1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire82_A (.DIODE(\sine_out_temp1[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[10]  (.DIODE(\sine_out_temp1[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire81_A (.DIODE(\sine_out_temp1[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[11]  (.DIODE(\sine_out_temp1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire80_A (.DIODE(\sine_out_temp1[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[12]  (.DIODE(\sine_out_temp1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire79_A (.DIODE(\sine_out_temp1[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[13]  (.DIODE(\sine_out_temp1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire78_A (.DIODE(\sine_out_temp1[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[14]  (.DIODE(\sine_out_temp1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire77_A (.DIODE(\sine_out_temp1[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[15]  (.DIODE(\sine_out_temp1[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire76_A (.DIODE(\sine_out_temp1[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[1]  (.DIODE(\sine_out_temp1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire75_A (.DIODE(\sine_out_temp1[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[2]  (.DIODE(\sine_out_temp1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire74_A (.DIODE(\sine_out_temp1[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[3]  (.DIODE(\sine_out_temp1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire73_A (.DIODE(\sine_out_temp1[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[4]  (.DIODE(\sine_out_temp1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire72_A (.DIODE(\sine_out_temp1[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[5]  (.DIODE(\sine_out_temp1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire71_A (.DIODE(\sine_out_temp1[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[6]  (.DIODE(\sine_out_temp1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire70_A (.DIODE(\sine_out_temp1[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[7]  (.DIODE(\sine_out_temp1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire69_A (.DIODE(\sine_out_temp1[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[8]  (.DIODE(\sine_out_temp1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire68_A (.DIODE(\sine_out_temp1[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_dout1[9]  (.DIODE(\sine_out_temp1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(\tcout[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(\tcout[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__Q (.DIODE(\tcout[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[0]  (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[1]  (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[2]  (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[3]  (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[4]  (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[5]  (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[6]  (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr0[7]  (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr0[2]  (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr0[3]  (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr0[4]  (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr0[5]  (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr0[6]  (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr0[7]  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[0]  (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[1]  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[2]  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[3]  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[4]  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[5]  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[6]  (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[7]  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_din0[8]  (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__Q (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__Q (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__Q (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__Q (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__Q (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output57_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__Q (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_output58_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__Q (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_output59_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__Q (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__Q (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_output61_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__Q (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__Q (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__Q (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__Q (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__Q (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__Q (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__Q (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire68_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__072__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire69_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire70_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire71_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire72_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire73_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire74_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__066__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire75_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__065__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire76_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__064__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire77_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__078__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire78_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__077__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire79_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__076__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire80_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire81_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__074__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire82_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire83_X (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__063__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire84_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__072__A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire85_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire86_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire87_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire88_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire89_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire90_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__066__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire91_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__065__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire92_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__064__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire93_X (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__078__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire94_X (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__077__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire95_X (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__076__A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire96_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire97_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__074__A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire98_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire99_X (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__063__A0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__095__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__078__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__077__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__076__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__074__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew103_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire102_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__091__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew104_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[7]  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew106_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__091__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew107_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew106_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__A3 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew108_X (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[6]  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew110_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew111_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[5]  (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew113_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__092__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew114_X (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[4]  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew117_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[3]  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew118_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire116_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew117_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew120_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire119_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__083__C (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew121_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[2]  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew123_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[1]  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew124_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire122_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew123_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew127_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[0]  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew128_X (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire126_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew127_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__107__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__119__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__118__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__117__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__116__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__115__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__114__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__113__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__112__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__111__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__105__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__104__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__103__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__106__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__102__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload0_A (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__CLK (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__CLK (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__CLK (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__CLK (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i0_clk0 (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_clk_X (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload1_A (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__CLK (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__CLK (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__CLK (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__CLK (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__CLK (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__CLK (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i0_clk1 (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_clk_X (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload2_A (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__CLK (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__CLK (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__132__CLK (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__133__CLK (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__134__CLK (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__CLK (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i1_clk0 (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_clk_X (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__CLK (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__CLK (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__CLK (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__CLK (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__128__CLK (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__129__CLK (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__CLK (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__131__CLK (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__CLK (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i1_clk1 (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_clk_X (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net128));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1425 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1433 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1442 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1509 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1521 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1543 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1555 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1579 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1591 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2169 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1476 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1480 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1494 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1506 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1517 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2199 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2573 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1340 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1363 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1330 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1328 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1344 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2580 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1328 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2434 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_2446 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2434 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2446 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2458 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_2470 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1316 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1178 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1272 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1279 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1336 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2434 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_2446 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1356 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1368 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1316 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1312 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1344 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1232 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1356 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1344 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1364 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1344 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1364 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1328 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1344 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1340 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1366 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1344 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1367 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1342 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1260 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1303 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1316 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2429 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_2441 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_2474 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_2478 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2492 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2516 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_2528 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_2534 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2438 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2476 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2488 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_2506 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2508 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2532 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2544 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_2562 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_2576 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1509 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1567 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1578 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1590 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1601 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1613 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1622 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1625 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1633 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1650 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1664 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1687 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1695 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1705 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1714 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1734 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1750 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1769 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1779 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1795 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1807 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1823 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1835 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1851 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1863 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1879 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1891 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1899 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1917 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1953 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1958 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1973 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1981 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_2001 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2009 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_2012 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_2029 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2037 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_2040 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_2057 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_2067 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2073 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_2085 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2091 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2125 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2129 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_2138 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2321 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_2325 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_2333 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_2573 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_2575 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_2573 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_2577 ();
endmodule
